//=========================================================
//File name    : rename_in_agent_monitor.sv
//Author       : nanyunhao
//Module name  : rename_in_agent_monitor
//Discribution : rename_in_agent_monitor : monitor
//Date         : 2026-01-22
//=========================================================
`ifndef RENAME_IN_AGENT_MONITOR__SV
`define RENAME_IN_AGENT_MONITOR__SV

class rename_in_agent_monitor  extends tcnt_monitor_base#(virtual rename_in_agent_interface,rename_in_agent_cfg,rename_in_agent_xaction);

    `uvm_component_utils(rename_in_agent_monitor)

    extern function new(string name, uvm_component parent);
    extern virtual function void build_phase(uvm_phase phase);
    extern task run_phase(uvm_phase phase);
    extern task mon_data();
endclass:rename_in_agent_monitor

function rename_in_agent_monitor::new(string name, uvm_component parent);
    super.new(name,parent);
endfunction:new

function void rename_in_agent_monitor::build_phase(uvm_phase phase);
    super.build_phase(phase);
endfunction:build_phase

task rename_in_agent_monitor::run_phase(uvm_phase phase);
    super.run_phase(phase);
    this.mon_data();
endtask:run_phase

task rename_in_agent_monitor::mon_data();

    logic         clock                ;
    logic         reset                ;
    logic [5:0]   io_hartId            ;
    logic         io_enq_req_0_valid   ;
    logic [31:0]  io_enq_req_0_bits_instr;
    logic [49:0]  io_enq_req_0_bits_pc ;
    logic         io_enq_req_0_bits_exceptionVec_0;
    logic         io_enq_req_0_bits_exceptionVec_1;
    logic         io_enq_req_0_bits_exceptionVec_2;
    logic         io_enq_req_0_bits_exceptionVec_3;
    logic         io_enq_req_0_bits_exceptionVec_12;
    logic         io_enq_req_0_bits_exceptionVec_20;
    logic         io_enq_req_0_bits_exceptionVec_22;
    logic         io_enq_req_0_bits_isFetchMalAddr;
    logic         io_enq_req_0_bits_hasException;
    logic [3:0]   io_enq_req_0_bits_trigger;
    logic         io_enq_req_0_bits_preDecodeInfo_isRVC;
    logic         io_enq_req_0_bits_crossPageIPFFix;
    logic         io_enq_req_0_bits_ftqPtr_flag;
    logic [5:0]   io_enq_req_0_bits_ftqPtr_value;
    logic [3:0]   io_enq_req_0_bits_ftqOffset;
    logic [5:0]   io_enq_req_0_bits_ldest;
    logic [34:0]  io_enq_req_0_bits_fuType;
    logic [8:0]   io_enq_req_0_bits_fuOpType;
    logic         io_enq_req_0_bits_rfWen;
    logic         io_enq_req_0_bits_fpWen;
    logic         io_enq_req_0_bits_vecWen;
    logic         io_enq_req_0_bits_v0Wen;
    logic         io_enq_req_0_bits_vlWen;
    logic         io_enq_req_0_bits_isXSTrap;
    logic         io_enq_req_0_bits_waitForward;
    logic         io_enq_req_0_bits_blockBackward;
    logic         io_enq_req_0_bits_flushPipe;
    logic         io_enq_req_0_bits_vpu_vill;
    logic         io_enq_req_0_bits_vpu_vma;
    logic         io_enq_req_0_bits_vpu_vta;
    logic [1:0]   io_enq_req_0_bits_vpu_vsew;
    logic [2:0]   io_enq_req_0_bits_vpu_vlmul;
    logic         io_enq_req_0_bits_vpu_specVill;
    logic         io_enq_req_0_bits_vpu_specVma;
    logic         io_enq_req_0_bits_vpu_specVta;
    logic [1:0]   io_enq_req_0_bits_vpu_specVsew;
    logic [2:0]   io_enq_req_0_bits_vpu_specVlmul;
    logic         io_enq_req_0_bits_vlsInstr;
    logic         io_enq_req_0_bits_wfflags;
    logic         io_enq_req_0_bits_isMove;
    logic         io_enq_req_0_bits_isVset;
    logic         io_enq_req_0_bits_firstUop;
    logic         io_enq_req_0_bits_lastUop;
    logic [6:0]   io_enq_req_0_bits_numWB;
    logic [2:0]   io_enq_req_0_bits_commitType;
    logic [7:0]   io_enq_req_0_bits_pdest;
    logic         io_enq_req_0_bits_robIdx_flag;
    logic [7:0]   io_enq_req_0_bits_robIdx_value;
    logic [2:0]   io_enq_req_0_bits_instrSize;
    logic         io_enq_req_0_bits_dirtyFs;
    logic         io_enq_req_0_bits_dirtyVs;
    logic [3:0]   io_enq_req_0_bits_traceBlockInPipe_itype;
    logic [3:0]   io_enq_req_0_bits_traceBlockInPipe_iretire;
    logic         io_enq_req_0_bits_traceBlockInPipe_ilastsize;
    logic         io_enq_req_0_bits_eliminatedMove;
    logic         io_enq_req_0_bits_snapshot;
    logic [6:0]   io_enq_req_0_bits_lqIdx_value;
    logic [5:0]   io_enq_req_0_bits_sqIdx_value;
    logic         io_enq_req_0_bits_singleStep;
    logic         io_enq_req_0_bits_debug_sim_trig;
    logic         io_enq_req_1_valid   ;
    logic [31:0]  io_enq_req_1_bits_instr;
    logic [49:0]  io_enq_req_1_bits_pc ;
    logic         io_enq_req_1_bits_exceptionVec_0;
    logic         io_enq_req_1_bits_exceptionVec_1;
    logic         io_enq_req_1_bits_exceptionVec_2;
    logic         io_enq_req_1_bits_exceptionVec_3;
    logic         io_enq_req_1_bits_exceptionVec_12;
    logic         io_enq_req_1_bits_exceptionVec_20;
    logic         io_enq_req_1_bits_exceptionVec_22;
    logic         io_enq_req_1_bits_isFetchMalAddr;
    logic         io_enq_req_1_bits_hasException;
    logic [3:0]   io_enq_req_1_bits_trigger;
    logic         io_enq_req_1_bits_preDecodeInfo_isRVC;
    logic         io_enq_req_1_bits_crossPageIPFFix;
    logic         io_enq_req_1_bits_ftqPtr_flag;
    logic [5:0]   io_enq_req_1_bits_ftqPtr_value;
    logic [3:0]   io_enq_req_1_bits_ftqOffset;
    logic [5:0]   io_enq_req_1_bits_ldest;
    logic [34:0]  io_enq_req_1_bits_fuType;
    logic [8:0]   io_enq_req_1_bits_fuOpType;
    logic         io_enq_req_1_bits_rfWen;
    logic         io_enq_req_1_bits_fpWen;
    logic         io_enq_req_1_bits_vecWen;
    logic         io_enq_req_1_bits_v0Wen;
    logic         io_enq_req_1_bits_vlWen;
    logic         io_enq_req_1_bits_isXSTrap;
    logic         io_enq_req_1_bits_waitForward;
    logic         io_enq_req_1_bits_blockBackward;
    logic         io_enq_req_1_bits_flushPipe;
    logic         io_enq_req_1_bits_vpu_vill;
    logic         io_enq_req_1_bits_vpu_vma;
    logic         io_enq_req_1_bits_vpu_vta;
    logic [1:0]   io_enq_req_1_bits_vpu_vsew;
    logic [2:0]   io_enq_req_1_bits_vpu_vlmul;
    logic         io_enq_req_1_bits_vpu_specVill;
    logic         io_enq_req_1_bits_vpu_specVma;
    logic         io_enq_req_1_bits_vpu_specVta;
    logic [1:0]   io_enq_req_1_bits_vpu_specVsew;
    logic [2:0]   io_enq_req_1_bits_vpu_specVlmul;
    logic         io_enq_req_1_bits_vlsInstr;
    logic         io_enq_req_1_bits_wfflags;
    logic         io_enq_req_1_bits_isMove;
    logic         io_enq_req_1_bits_isVset;
    logic         io_enq_req_1_bits_firstUop;
    logic         io_enq_req_1_bits_lastUop;
    logic [6:0]   io_enq_req_1_bits_numWB;
    logic [2:0]   io_enq_req_1_bits_commitType;
    logic [7:0]   io_enq_req_1_bits_pdest;
    logic         io_enq_req_1_bits_robIdx_flag;
    logic [7:0]   io_enq_req_1_bits_robIdx_value;
    logic [2:0]   io_enq_req_1_bits_instrSize;
    logic         io_enq_req_1_bits_dirtyFs;
    logic         io_enq_req_1_bits_dirtyVs;
    logic [3:0]   io_enq_req_1_bits_traceBlockInPipe_itype;
    logic [3:0]   io_enq_req_1_bits_traceBlockInPipe_iretire;
    logic         io_enq_req_1_bits_traceBlockInPipe_ilastsize;
    logic         io_enq_req_1_bits_eliminatedMove;
    logic         io_enq_req_1_bits_snapshot;
    logic [6:0]   io_enq_req_1_bits_lqIdx_value;
    logic [5:0]   io_enq_req_1_bits_sqIdx_value;
    logic         io_enq_req_1_bits_singleStep;
    logic         io_enq_req_1_bits_debug_sim_trig;
    logic         io_enq_req_2_valid   ;
    logic [31:0]  io_enq_req_2_bits_instr;
    logic [49:0]  io_enq_req_2_bits_pc ;
    logic         io_enq_req_2_bits_exceptionVec_0;
    logic         io_enq_req_2_bits_exceptionVec_1;
    logic         io_enq_req_2_bits_exceptionVec_2;
    logic         io_enq_req_2_bits_exceptionVec_3;
    logic         io_enq_req_2_bits_exceptionVec_12;
    logic         io_enq_req_2_bits_exceptionVec_20;
    logic         io_enq_req_2_bits_exceptionVec_22;
    logic         io_enq_req_2_bits_isFetchMalAddr;
    logic         io_enq_req_2_bits_hasException;
    logic [3:0]   io_enq_req_2_bits_trigger;
    logic         io_enq_req_2_bits_preDecodeInfo_isRVC;
    logic         io_enq_req_2_bits_crossPageIPFFix;
    logic         io_enq_req_2_bits_ftqPtr_flag;
    logic [5:0]   io_enq_req_2_bits_ftqPtr_value;
    logic [3:0]   io_enq_req_2_bits_ftqOffset;
    logic [5:0]   io_enq_req_2_bits_ldest;
    logic [34:0]  io_enq_req_2_bits_fuType;
    logic [8:0]   io_enq_req_2_bits_fuOpType;
    logic         io_enq_req_2_bits_rfWen;
    logic         io_enq_req_2_bits_fpWen;
    logic         io_enq_req_2_bits_vecWen;
    logic         io_enq_req_2_bits_v0Wen;
    logic         io_enq_req_2_bits_vlWen;
    logic         io_enq_req_2_bits_isXSTrap;
    logic         io_enq_req_2_bits_waitForward;
    logic         io_enq_req_2_bits_blockBackward;
    logic         io_enq_req_2_bits_flushPipe;
    logic         io_enq_req_2_bits_vpu_vill;
    logic         io_enq_req_2_bits_vpu_vma;
    logic         io_enq_req_2_bits_vpu_vta;
    logic [1:0]   io_enq_req_2_bits_vpu_vsew;
    logic [2:0]   io_enq_req_2_bits_vpu_vlmul;
    logic         io_enq_req_2_bits_vpu_specVill;
    logic         io_enq_req_2_bits_vpu_specVma;
    logic         io_enq_req_2_bits_vpu_specVta;
    logic [1:0]   io_enq_req_2_bits_vpu_specVsew;
    logic [2:0]   io_enq_req_2_bits_vpu_specVlmul;
    logic         io_enq_req_2_bits_vlsInstr;
    logic         io_enq_req_2_bits_wfflags;
    logic         io_enq_req_2_bits_isMove;
    logic         io_enq_req_2_bits_isVset;
    logic         io_enq_req_2_bits_firstUop;
    logic         io_enq_req_2_bits_lastUop;
    logic [6:0]   io_enq_req_2_bits_numWB;
    logic [2:0]   io_enq_req_2_bits_commitType;
    logic [7:0]   io_enq_req_2_bits_pdest;
    logic         io_enq_req_2_bits_robIdx_flag;
    logic [7:0]   io_enq_req_2_bits_robIdx_value;
    logic [2:0]   io_enq_req_2_bits_instrSize;
    logic         io_enq_req_2_bits_dirtyFs;
    logic         io_enq_req_2_bits_dirtyVs;
    logic [3:0]   io_enq_req_2_bits_traceBlockInPipe_itype;
    logic [3:0]   io_enq_req_2_bits_traceBlockInPipe_iretire;
    logic         io_enq_req_2_bits_traceBlockInPipe_ilastsize;
    logic         io_enq_req_2_bits_eliminatedMove;
    logic         io_enq_req_2_bits_snapshot;
    logic [6:0]   io_enq_req_2_bits_lqIdx_value;
    logic [5:0]   io_enq_req_2_bits_sqIdx_value;
    logic         io_enq_req_2_bits_singleStep;
    logic         io_enq_req_2_bits_debug_sim_trig;
    logic         io_enq_req_3_valid   ;
    logic [31:0]  io_enq_req_3_bits_instr;
    logic [49:0]  io_enq_req_3_bits_pc ;
    logic         io_enq_req_3_bits_exceptionVec_0;
    logic         io_enq_req_3_bits_exceptionVec_1;
    logic         io_enq_req_3_bits_exceptionVec_2;
    logic         io_enq_req_3_bits_exceptionVec_3;
    logic         io_enq_req_3_bits_exceptionVec_12;
    logic         io_enq_req_3_bits_exceptionVec_20;
    logic         io_enq_req_3_bits_exceptionVec_22;
    logic         io_enq_req_3_bits_isFetchMalAddr;
    logic         io_enq_req_3_bits_hasException;
    logic [3:0]   io_enq_req_3_bits_trigger;
    logic         io_enq_req_3_bits_preDecodeInfo_isRVC;
    logic         io_enq_req_3_bits_crossPageIPFFix;
    logic         io_enq_req_3_bits_ftqPtr_flag;
    logic [5:0]   io_enq_req_3_bits_ftqPtr_value;
    logic [3:0]   io_enq_req_3_bits_ftqOffset;
    logic [5:0]   io_enq_req_3_bits_ldest;
    logic [34:0]  io_enq_req_3_bits_fuType;
    logic [8:0]   io_enq_req_3_bits_fuOpType;
    logic         io_enq_req_3_bits_rfWen;
    logic         io_enq_req_3_bits_fpWen;
    logic         io_enq_req_3_bits_vecWen;
    logic         io_enq_req_3_bits_v0Wen;
    logic         io_enq_req_3_bits_vlWen;
    logic         io_enq_req_3_bits_isXSTrap;
    logic         io_enq_req_3_bits_waitForward;
    logic         io_enq_req_3_bits_blockBackward;
    logic         io_enq_req_3_bits_flushPipe;
    logic         io_enq_req_3_bits_vpu_vill;
    logic         io_enq_req_3_bits_vpu_vma;
    logic         io_enq_req_3_bits_vpu_vta;
    logic [1:0]   io_enq_req_3_bits_vpu_vsew;
    logic [2:0]   io_enq_req_3_bits_vpu_vlmul;
    logic         io_enq_req_3_bits_vpu_specVill;
    logic         io_enq_req_3_bits_vpu_specVma;
    logic         io_enq_req_3_bits_vpu_specVta;
    logic [1:0]   io_enq_req_3_bits_vpu_specVsew;
    logic [2:0]   io_enq_req_3_bits_vpu_specVlmul;
    logic         io_enq_req_3_bits_vlsInstr;
    logic         io_enq_req_3_bits_wfflags;
    logic         io_enq_req_3_bits_isMove;
    logic         io_enq_req_3_bits_isVset;
    logic         io_enq_req_3_bits_firstUop;
    logic         io_enq_req_3_bits_lastUop;
    logic [6:0]   io_enq_req_3_bits_numWB;
    logic [2:0]   io_enq_req_3_bits_commitType;
    logic [7:0]   io_enq_req_3_bits_pdest;
    logic         io_enq_req_3_bits_robIdx_flag;
    logic [7:0]   io_enq_req_3_bits_robIdx_value;
    logic [2:0]   io_enq_req_3_bits_instrSize;
    logic         io_enq_req_3_bits_dirtyFs;
    logic         io_enq_req_3_bits_dirtyVs;
    logic [3:0]   io_enq_req_3_bits_traceBlockInPipe_itype;
    logic [3:0]   io_enq_req_3_bits_traceBlockInPipe_iretire;
    logic         io_enq_req_3_bits_traceBlockInPipe_ilastsize;
    logic         io_enq_req_3_bits_eliminatedMove;
    logic         io_enq_req_3_bits_snapshot;
    logic [6:0]   io_enq_req_3_bits_lqIdx_value;
    logic [5:0]   io_enq_req_3_bits_sqIdx_value;
    logic         io_enq_req_3_bits_singleStep;
    logic         io_enq_req_3_bits_debug_sim_trig;
    logic         io_enq_req_4_valid   ;
    logic [31:0]  io_enq_req_4_bits_instr;
    logic [49:0]  io_enq_req_4_bits_pc ;
    logic         io_enq_req_4_bits_exceptionVec_0;
    logic         io_enq_req_4_bits_exceptionVec_1;
    logic         io_enq_req_4_bits_exceptionVec_2;
    logic         io_enq_req_4_bits_exceptionVec_3;
    logic         io_enq_req_4_bits_exceptionVec_12;
    logic         io_enq_req_4_bits_exceptionVec_20;
    logic         io_enq_req_4_bits_exceptionVec_22;
    logic         io_enq_req_4_bits_isFetchMalAddr;
    logic         io_enq_req_4_bits_hasException;
    logic [3:0]   io_enq_req_4_bits_trigger;
    logic         io_enq_req_4_bits_preDecodeInfo_isRVC;
    logic         io_enq_req_4_bits_crossPageIPFFix;
    logic         io_enq_req_4_bits_ftqPtr_flag;
    logic [5:0]   io_enq_req_4_bits_ftqPtr_value;
    logic [3:0]   io_enq_req_4_bits_ftqOffset;
    logic [5:0]   io_enq_req_4_bits_ldest;
    logic [34:0]  io_enq_req_4_bits_fuType;
    logic [8:0]   io_enq_req_4_bits_fuOpType;
    logic         io_enq_req_4_bits_rfWen;
    logic         io_enq_req_4_bits_fpWen;
    logic         io_enq_req_4_bits_vecWen;
    logic         io_enq_req_4_bits_v0Wen;
    logic         io_enq_req_4_bits_vlWen;
    logic         io_enq_req_4_bits_isXSTrap;
    logic         io_enq_req_4_bits_waitForward;
    logic         io_enq_req_4_bits_blockBackward;
    logic         io_enq_req_4_bits_flushPipe;
    logic         io_enq_req_4_bits_vpu_vill;
    logic         io_enq_req_4_bits_vpu_vma;
    logic         io_enq_req_4_bits_vpu_vta;
    logic [1:0]   io_enq_req_4_bits_vpu_vsew;
    logic [2:0]   io_enq_req_4_bits_vpu_vlmul;
    logic         io_enq_req_4_bits_vpu_specVill;
    logic         io_enq_req_4_bits_vpu_specVma;
    logic         io_enq_req_4_bits_vpu_specVta;
    logic [1:0]   io_enq_req_4_bits_vpu_specVsew;
    logic [2:0]   io_enq_req_4_bits_vpu_specVlmul;
    logic         io_enq_req_4_bits_vlsInstr;
    logic         io_enq_req_4_bits_wfflags;
    logic         io_enq_req_4_bits_isMove;
    logic         io_enq_req_4_bits_isVset;
    logic         io_enq_req_4_bits_firstUop;
    logic         io_enq_req_4_bits_lastUop;
    logic [6:0]   io_enq_req_4_bits_numWB;
    logic [2:0]   io_enq_req_4_bits_commitType;
    logic [7:0]   io_enq_req_4_bits_pdest;
    logic         io_enq_req_4_bits_robIdx_flag;
    logic [7:0]   io_enq_req_4_bits_robIdx_value;
    logic [2:0]   io_enq_req_4_bits_instrSize;
    logic         io_enq_req_4_bits_dirtyFs;
    logic         io_enq_req_4_bits_dirtyVs;
    logic [3:0]   io_enq_req_4_bits_traceBlockInPipe_itype;
    logic [3:0]   io_enq_req_4_bits_traceBlockInPipe_iretire;
    logic         io_enq_req_4_bits_traceBlockInPipe_ilastsize;
    logic         io_enq_req_4_bits_eliminatedMove;
    logic         io_enq_req_4_bits_snapshot;
    logic [6:0]   io_enq_req_4_bits_lqIdx_value;
    logic [5:0]   io_enq_req_4_bits_sqIdx_value;
    logic         io_enq_req_4_bits_singleStep;
    logic         io_enq_req_4_bits_debug_sim_trig;
    logic         io_enq_req_5_valid   ;
    logic [31:0]  io_enq_req_5_bits_instr;
    logic [49:0]  io_enq_req_5_bits_pc ;
    logic         io_enq_req_5_bits_exceptionVec_0;
    logic         io_enq_req_5_bits_exceptionVec_1;
    logic         io_enq_req_5_bits_exceptionVec_2;
    logic         io_enq_req_5_bits_exceptionVec_3;
    logic         io_enq_req_5_bits_exceptionVec_12;
    logic         io_enq_req_5_bits_exceptionVec_20;
    logic         io_enq_req_5_bits_exceptionVec_22;
    logic         io_enq_req_5_bits_isFetchMalAddr;
    logic         io_enq_req_5_bits_hasException;
    logic [3:0]   io_enq_req_5_bits_trigger;
    logic         io_enq_req_5_bits_preDecodeInfo_isRVC;
    logic         io_enq_req_5_bits_crossPageIPFFix;
    logic         io_enq_req_5_bits_ftqPtr_flag;
    logic [5:0]   io_enq_req_5_bits_ftqPtr_value;
    logic [3:0]   io_enq_req_5_bits_ftqOffset;
    logic [5:0]   io_enq_req_5_bits_ldest;
    logic [34:0]  io_enq_req_5_bits_fuType;
    logic [8:0]   io_enq_req_5_bits_fuOpType;
    logic         io_enq_req_5_bits_rfWen;
    logic         io_enq_req_5_bits_fpWen;
    logic         io_enq_req_5_bits_vecWen;
    logic         io_enq_req_5_bits_v0Wen;
    logic         io_enq_req_5_bits_vlWen;
    logic         io_enq_req_5_bits_isXSTrap;
    logic         io_enq_req_5_bits_waitForward;
    logic         io_enq_req_5_bits_blockBackward;
    logic         io_enq_req_5_bits_flushPipe;
    logic         io_enq_req_5_bits_vpu_vill;
    logic         io_enq_req_5_bits_vpu_vma;
    logic         io_enq_req_5_bits_vpu_vta;
    logic [1:0]   io_enq_req_5_bits_vpu_vsew;
    logic [2:0]   io_enq_req_5_bits_vpu_vlmul;
    logic         io_enq_req_5_bits_vpu_specVill;
    logic         io_enq_req_5_bits_vpu_specVma;
    logic         io_enq_req_5_bits_vpu_specVta;
    logic [1:0]   io_enq_req_5_bits_vpu_specVsew;
    logic [2:0]   io_enq_req_5_bits_vpu_specVlmul;
    logic         io_enq_req_5_bits_vlsInstr;
    logic         io_enq_req_5_bits_wfflags;
    logic         io_enq_req_5_bits_isMove;
    logic         io_enq_req_5_bits_isVset;
    logic         io_enq_req_5_bits_firstUop;
    logic         io_enq_req_5_bits_lastUop;
    logic [6:0]   io_enq_req_5_bits_numWB;
    logic [2:0]   io_enq_req_5_bits_commitType;
    logic [7:0]   io_enq_req_5_bits_pdest;
    logic         io_enq_req_5_bits_robIdx_flag;
    logic [7:0]   io_enq_req_5_bits_robIdx_value;
    logic [2:0]   io_enq_req_5_bits_instrSize;
    logic         io_enq_req_5_bits_dirtyFs;
    logic         io_enq_req_5_bits_dirtyVs;
    logic [3:0]   io_enq_req_5_bits_traceBlockInPipe_itype;
    logic [3:0]   io_enq_req_5_bits_traceBlockInPipe_iretire;
    logic         io_enq_req_5_bits_traceBlockInPipe_ilastsize;
    logic         io_enq_req_5_bits_eliminatedMove;
    logic         io_enq_req_5_bits_snapshot;
    logic [6:0]   io_enq_req_5_bits_lqIdx_value;
    logic [5:0]   io_enq_req_5_bits_sqIdx_value;
    logic         io_enq_req_5_bits_singleStep;
    logic         io_enq_req_5_bits_debug_sim_trig;

    rename_in_agent_xaction  mon_tr;
    while(1) begin
        @this.vif.mon_mp.mon_cb;
        clock = this.vif.mon_mp.mon_cb.clock;
        reset = this.vif.mon_mp.mon_cb.reset;
        io_hartId = this.vif.mon_mp.mon_cb.io_hartId;
        io_enq_req_0_valid = this.vif.mon_mp.mon_cb.io_enq_req_0_valid;
        io_enq_req_0_bits_instr = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_instr;
        io_enq_req_0_bits_pc = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_pc;
        io_enq_req_0_bits_exceptionVec_0 = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_exceptionVec_0;
        io_enq_req_0_bits_exceptionVec_1 = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_exceptionVec_1;
        io_enq_req_0_bits_exceptionVec_2 = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_exceptionVec_2;
        io_enq_req_0_bits_exceptionVec_3 = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_exceptionVec_3;
        io_enq_req_0_bits_exceptionVec_12 = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_exceptionVec_12;
        io_enq_req_0_bits_exceptionVec_20 = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_exceptionVec_20;
        io_enq_req_0_bits_exceptionVec_22 = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_exceptionVec_22;
        io_enq_req_0_bits_isFetchMalAddr = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_isFetchMalAddr;
        io_enq_req_0_bits_hasException = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_hasException;
        io_enq_req_0_bits_trigger = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_trigger;
        io_enq_req_0_bits_preDecodeInfo_isRVC = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_preDecodeInfo_isRVC;
        io_enq_req_0_bits_crossPageIPFFix = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_crossPageIPFFix;
        io_enq_req_0_bits_ftqPtr_flag = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_ftqPtr_flag;
        io_enq_req_0_bits_ftqPtr_value = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_ftqPtr_value;
        io_enq_req_0_bits_ftqOffset = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_ftqOffset;
        io_enq_req_0_bits_ldest = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_ldest;
        io_enq_req_0_bits_fuType = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_fuType;
        io_enq_req_0_bits_fuOpType = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_fuOpType;
        io_enq_req_0_bits_rfWen = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_rfWen;
        io_enq_req_0_bits_fpWen = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_fpWen;
        io_enq_req_0_bits_vecWen = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_vecWen;
        io_enq_req_0_bits_v0Wen = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_v0Wen;
        io_enq_req_0_bits_vlWen = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_vlWen;
        io_enq_req_0_bits_isXSTrap = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_isXSTrap;
        io_enq_req_0_bits_waitForward = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_waitForward;
        io_enq_req_0_bits_blockBackward = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_blockBackward;
        io_enq_req_0_bits_flushPipe = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_flushPipe;
        io_enq_req_0_bits_vpu_vill = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_vpu_vill;
        io_enq_req_0_bits_vpu_vma = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_vpu_vma;
        io_enq_req_0_bits_vpu_vta = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_vpu_vta;
        io_enq_req_0_bits_vpu_vsew = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_vpu_vsew;
        io_enq_req_0_bits_vpu_vlmul = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_vpu_vlmul;
        io_enq_req_0_bits_vpu_specVill = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_vpu_specVill;
        io_enq_req_0_bits_vpu_specVma = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_vpu_specVma;
        io_enq_req_0_bits_vpu_specVta = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_vpu_specVta;
        io_enq_req_0_bits_vpu_specVsew = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_vpu_specVsew;
        io_enq_req_0_bits_vpu_specVlmul = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_vpu_specVlmul;
        io_enq_req_0_bits_vlsInstr = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_vlsInstr;
        io_enq_req_0_bits_wfflags = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_wfflags;
        io_enq_req_0_bits_isMove = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_isMove;
        io_enq_req_0_bits_isVset = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_isVset;
        io_enq_req_0_bits_firstUop = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_firstUop;
        io_enq_req_0_bits_lastUop = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_lastUop;
        io_enq_req_0_bits_numWB = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_numWB;
        io_enq_req_0_bits_commitType = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_commitType;
        io_enq_req_0_bits_pdest = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_pdest;
        io_enq_req_0_bits_robIdx_flag = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_robIdx_flag;
        io_enq_req_0_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_robIdx_value;
        io_enq_req_0_bits_instrSize = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_instrSize;
        io_enq_req_0_bits_dirtyFs = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_dirtyFs;
        io_enq_req_0_bits_dirtyVs = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_dirtyVs;
        io_enq_req_0_bits_traceBlockInPipe_itype = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_traceBlockInPipe_itype;
        io_enq_req_0_bits_traceBlockInPipe_iretire = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_traceBlockInPipe_iretire;
        io_enq_req_0_bits_traceBlockInPipe_ilastsize = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_traceBlockInPipe_ilastsize;
        io_enq_req_0_bits_eliminatedMove = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_eliminatedMove;
        io_enq_req_0_bits_snapshot = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_snapshot;
        io_enq_req_0_bits_lqIdx_value = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_lqIdx_value;
        io_enq_req_0_bits_sqIdx_value = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_sqIdx_value;
        io_enq_req_0_bits_singleStep = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_singleStep;
        io_enq_req_0_bits_debug_sim_trig = this.vif.mon_mp.mon_cb.io_enq_req_0_bits_debug_sim_trig;
        io_enq_req_1_valid = this.vif.mon_mp.mon_cb.io_enq_req_1_valid;
        io_enq_req_1_bits_instr = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_instr;
        io_enq_req_1_bits_pc = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_pc;
        io_enq_req_1_bits_exceptionVec_0 = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_exceptionVec_0;
        io_enq_req_1_bits_exceptionVec_1 = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_exceptionVec_1;
        io_enq_req_1_bits_exceptionVec_2 = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_exceptionVec_2;
        io_enq_req_1_bits_exceptionVec_3 = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_exceptionVec_3;
        io_enq_req_1_bits_exceptionVec_12 = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_exceptionVec_12;
        io_enq_req_1_bits_exceptionVec_20 = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_exceptionVec_20;
        io_enq_req_1_bits_exceptionVec_22 = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_exceptionVec_22;
        io_enq_req_1_bits_isFetchMalAddr = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_isFetchMalAddr;
        io_enq_req_1_bits_hasException = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_hasException;
        io_enq_req_1_bits_trigger = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_trigger;
        io_enq_req_1_bits_preDecodeInfo_isRVC = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_preDecodeInfo_isRVC;
        io_enq_req_1_bits_crossPageIPFFix = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_crossPageIPFFix;
        io_enq_req_1_bits_ftqPtr_flag = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_ftqPtr_flag;
        io_enq_req_1_bits_ftqPtr_value = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_ftqPtr_value;
        io_enq_req_1_bits_ftqOffset = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_ftqOffset;
        io_enq_req_1_bits_ldest = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_ldest;
        io_enq_req_1_bits_fuType = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_fuType;
        io_enq_req_1_bits_fuOpType = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_fuOpType;
        io_enq_req_1_bits_rfWen = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_rfWen;
        io_enq_req_1_bits_fpWen = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_fpWen;
        io_enq_req_1_bits_vecWen = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_vecWen;
        io_enq_req_1_bits_v0Wen = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_v0Wen;
        io_enq_req_1_bits_vlWen = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_vlWen;
        io_enq_req_1_bits_isXSTrap = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_isXSTrap;
        io_enq_req_1_bits_waitForward = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_waitForward;
        io_enq_req_1_bits_blockBackward = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_blockBackward;
        io_enq_req_1_bits_flushPipe = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_flushPipe;
        io_enq_req_1_bits_vpu_vill = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_vpu_vill;
        io_enq_req_1_bits_vpu_vma = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_vpu_vma;
        io_enq_req_1_bits_vpu_vta = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_vpu_vta;
        io_enq_req_1_bits_vpu_vsew = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_vpu_vsew;
        io_enq_req_1_bits_vpu_vlmul = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_vpu_vlmul;
        io_enq_req_1_bits_vpu_specVill = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_vpu_specVill;
        io_enq_req_1_bits_vpu_specVma = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_vpu_specVma;
        io_enq_req_1_bits_vpu_specVta = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_vpu_specVta;
        io_enq_req_1_bits_vpu_specVsew = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_vpu_specVsew;
        io_enq_req_1_bits_vpu_specVlmul = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_vpu_specVlmul;
        io_enq_req_1_bits_vlsInstr = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_vlsInstr;
        io_enq_req_1_bits_wfflags = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_wfflags;
        io_enq_req_1_bits_isMove = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_isMove;
        io_enq_req_1_bits_isVset = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_isVset;
        io_enq_req_1_bits_firstUop = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_firstUop;
        io_enq_req_1_bits_lastUop = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_lastUop;
        io_enq_req_1_bits_numWB = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_numWB;
        io_enq_req_1_bits_commitType = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_commitType;
        io_enq_req_1_bits_pdest = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_pdest;
        io_enq_req_1_bits_robIdx_flag = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_robIdx_flag;
        io_enq_req_1_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_robIdx_value;
        io_enq_req_1_bits_instrSize = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_instrSize;
        io_enq_req_1_bits_dirtyFs = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_dirtyFs;
        io_enq_req_1_bits_dirtyVs = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_dirtyVs;
        io_enq_req_1_bits_traceBlockInPipe_itype = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_traceBlockInPipe_itype;
        io_enq_req_1_bits_traceBlockInPipe_iretire = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_traceBlockInPipe_iretire;
        io_enq_req_1_bits_traceBlockInPipe_ilastsize = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_traceBlockInPipe_ilastsize;
        io_enq_req_1_bits_eliminatedMove = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_eliminatedMove;
        io_enq_req_1_bits_snapshot = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_snapshot;
        io_enq_req_1_bits_lqIdx_value = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_lqIdx_value;
        io_enq_req_1_bits_sqIdx_value = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_sqIdx_value;
        io_enq_req_1_bits_singleStep = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_singleStep;
        io_enq_req_1_bits_debug_sim_trig = this.vif.mon_mp.mon_cb.io_enq_req_1_bits_debug_sim_trig;
        io_enq_req_2_valid = this.vif.mon_mp.mon_cb.io_enq_req_2_valid;
        io_enq_req_2_bits_instr = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_instr;
        io_enq_req_2_bits_pc = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_pc;
        io_enq_req_2_bits_exceptionVec_0 = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_exceptionVec_0;
        io_enq_req_2_bits_exceptionVec_1 = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_exceptionVec_1;
        io_enq_req_2_bits_exceptionVec_2 = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_exceptionVec_2;
        io_enq_req_2_bits_exceptionVec_3 = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_exceptionVec_3;
        io_enq_req_2_bits_exceptionVec_12 = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_exceptionVec_12;
        io_enq_req_2_bits_exceptionVec_20 = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_exceptionVec_20;
        io_enq_req_2_bits_exceptionVec_22 = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_exceptionVec_22;
        io_enq_req_2_bits_isFetchMalAddr = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_isFetchMalAddr;
        io_enq_req_2_bits_hasException = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_hasException;
        io_enq_req_2_bits_trigger = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_trigger;
        io_enq_req_2_bits_preDecodeInfo_isRVC = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_preDecodeInfo_isRVC;
        io_enq_req_2_bits_crossPageIPFFix = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_crossPageIPFFix;
        io_enq_req_2_bits_ftqPtr_flag = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_ftqPtr_flag;
        io_enq_req_2_bits_ftqPtr_value = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_ftqPtr_value;
        io_enq_req_2_bits_ftqOffset = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_ftqOffset;
        io_enq_req_2_bits_ldest = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_ldest;
        io_enq_req_2_bits_fuType = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_fuType;
        io_enq_req_2_bits_fuOpType = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_fuOpType;
        io_enq_req_2_bits_rfWen = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_rfWen;
        io_enq_req_2_bits_fpWen = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_fpWen;
        io_enq_req_2_bits_vecWen = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_vecWen;
        io_enq_req_2_bits_v0Wen = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_v0Wen;
        io_enq_req_2_bits_vlWen = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_vlWen;
        io_enq_req_2_bits_isXSTrap = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_isXSTrap;
        io_enq_req_2_bits_waitForward = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_waitForward;
        io_enq_req_2_bits_blockBackward = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_blockBackward;
        io_enq_req_2_bits_flushPipe = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_flushPipe;
        io_enq_req_2_bits_vpu_vill = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_vpu_vill;
        io_enq_req_2_bits_vpu_vma = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_vpu_vma;
        io_enq_req_2_bits_vpu_vta = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_vpu_vta;
        io_enq_req_2_bits_vpu_vsew = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_vpu_vsew;
        io_enq_req_2_bits_vpu_vlmul = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_vpu_vlmul;
        io_enq_req_2_bits_vpu_specVill = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_vpu_specVill;
        io_enq_req_2_bits_vpu_specVma = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_vpu_specVma;
        io_enq_req_2_bits_vpu_specVta = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_vpu_specVta;
        io_enq_req_2_bits_vpu_specVsew = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_vpu_specVsew;
        io_enq_req_2_bits_vpu_specVlmul = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_vpu_specVlmul;
        io_enq_req_2_bits_vlsInstr = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_vlsInstr;
        io_enq_req_2_bits_wfflags = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_wfflags;
        io_enq_req_2_bits_isMove = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_isMove;
        io_enq_req_2_bits_isVset = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_isVset;
        io_enq_req_2_bits_firstUop = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_firstUop;
        io_enq_req_2_bits_lastUop = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_lastUop;
        io_enq_req_2_bits_numWB = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_numWB;
        io_enq_req_2_bits_commitType = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_commitType;
        io_enq_req_2_bits_pdest = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_pdest;
        io_enq_req_2_bits_robIdx_flag = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_robIdx_flag;
        io_enq_req_2_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_robIdx_value;
        io_enq_req_2_bits_instrSize = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_instrSize;
        io_enq_req_2_bits_dirtyFs = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_dirtyFs;
        io_enq_req_2_bits_dirtyVs = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_dirtyVs;
        io_enq_req_2_bits_traceBlockInPipe_itype = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_traceBlockInPipe_itype;
        io_enq_req_2_bits_traceBlockInPipe_iretire = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_traceBlockInPipe_iretire;
        io_enq_req_2_bits_traceBlockInPipe_ilastsize = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_traceBlockInPipe_ilastsize;
        io_enq_req_2_bits_eliminatedMove = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_eliminatedMove;
        io_enq_req_2_bits_snapshot = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_snapshot;
        io_enq_req_2_bits_lqIdx_value = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_lqIdx_value;
        io_enq_req_2_bits_sqIdx_value = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_sqIdx_value;
        io_enq_req_2_bits_singleStep = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_singleStep;
        io_enq_req_2_bits_debug_sim_trig = this.vif.mon_mp.mon_cb.io_enq_req_2_bits_debug_sim_trig;
        io_enq_req_3_valid = this.vif.mon_mp.mon_cb.io_enq_req_3_valid;
        io_enq_req_3_bits_instr = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_instr;
        io_enq_req_3_bits_pc = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_pc;
        io_enq_req_3_bits_exceptionVec_0 = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_exceptionVec_0;
        io_enq_req_3_bits_exceptionVec_1 = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_exceptionVec_1;
        io_enq_req_3_bits_exceptionVec_2 = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_exceptionVec_2;
        io_enq_req_3_bits_exceptionVec_3 = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_exceptionVec_3;
        io_enq_req_3_bits_exceptionVec_12 = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_exceptionVec_12;
        io_enq_req_3_bits_exceptionVec_20 = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_exceptionVec_20;
        io_enq_req_3_bits_exceptionVec_22 = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_exceptionVec_22;
        io_enq_req_3_bits_isFetchMalAddr = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_isFetchMalAddr;
        io_enq_req_3_bits_hasException = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_hasException;
        io_enq_req_3_bits_trigger = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_trigger;
        io_enq_req_3_bits_preDecodeInfo_isRVC = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_preDecodeInfo_isRVC;
        io_enq_req_3_bits_crossPageIPFFix = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_crossPageIPFFix;
        io_enq_req_3_bits_ftqPtr_flag = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_ftqPtr_flag;
        io_enq_req_3_bits_ftqPtr_value = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_ftqPtr_value;
        io_enq_req_3_bits_ftqOffset = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_ftqOffset;
        io_enq_req_3_bits_ldest = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_ldest;
        io_enq_req_3_bits_fuType = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_fuType;
        io_enq_req_3_bits_fuOpType = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_fuOpType;
        io_enq_req_3_bits_rfWen = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_rfWen;
        io_enq_req_3_bits_fpWen = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_fpWen;
        io_enq_req_3_bits_vecWen = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_vecWen;
        io_enq_req_3_bits_v0Wen = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_v0Wen;
        io_enq_req_3_bits_vlWen = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_vlWen;
        io_enq_req_3_bits_isXSTrap = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_isXSTrap;
        io_enq_req_3_bits_waitForward = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_waitForward;
        io_enq_req_3_bits_blockBackward = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_blockBackward;
        io_enq_req_3_bits_flushPipe = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_flushPipe;
        io_enq_req_3_bits_vpu_vill = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_vpu_vill;
        io_enq_req_3_bits_vpu_vma = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_vpu_vma;
        io_enq_req_3_bits_vpu_vta = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_vpu_vta;
        io_enq_req_3_bits_vpu_vsew = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_vpu_vsew;
        io_enq_req_3_bits_vpu_vlmul = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_vpu_vlmul;
        io_enq_req_3_bits_vpu_specVill = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_vpu_specVill;
        io_enq_req_3_bits_vpu_specVma = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_vpu_specVma;
        io_enq_req_3_bits_vpu_specVta = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_vpu_specVta;
        io_enq_req_3_bits_vpu_specVsew = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_vpu_specVsew;
        io_enq_req_3_bits_vpu_specVlmul = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_vpu_specVlmul;
        io_enq_req_3_bits_vlsInstr = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_vlsInstr;
        io_enq_req_3_bits_wfflags = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_wfflags;
        io_enq_req_3_bits_isMove = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_isMove;
        io_enq_req_3_bits_isVset = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_isVset;
        io_enq_req_3_bits_firstUop = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_firstUop;
        io_enq_req_3_bits_lastUop = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_lastUop;
        io_enq_req_3_bits_numWB = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_numWB;
        io_enq_req_3_bits_commitType = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_commitType;
        io_enq_req_3_bits_pdest = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_pdest;
        io_enq_req_3_bits_robIdx_flag = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_robIdx_flag;
        io_enq_req_3_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_robIdx_value;
        io_enq_req_3_bits_instrSize = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_instrSize;
        io_enq_req_3_bits_dirtyFs = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_dirtyFs;
        io_enq_req_3_bits_dirtyVs = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_dirtyVs;
        io_enq_req_3_bits_traceBlockInPipe_itype = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_traceBlockInPipe_itype;
        io_enq_req_3_bits_traceBlockInPipe_iretire = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_traceBlockInPipe_iretire;
        io_enq_req_3_bits_traceBlockInPipe_ilastsize = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_traceBlockInPipe_ilastsize;
        io_enq_req_3_bits_eliminatedMove = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_eliminatedMove;
        io_enq_req_3_bits_snapshot = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_snapshot;
        io_enq_req_3_bits_lqIdx_value = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_lqIdx_value;
        io_enq_req_3_bits_sqIdx_value = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_sqIdx_value;
        io_enq_req_3_bits_singleStep = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_singleStep;
        io_enq_req_3_bits_debug_sim_trig = this.vif.mon_mp.mon_cb.io_enq_req_3_bits_debug_sim_trig;
        io_enq_req_4_valid = this.vif.mon_mp.mon_cb.io_enq_req_4_valid;
        io_enq_req_4_bits_instr = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_instr;
        io_enq_req_4_bits_pc = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_pc;
        io_enq_req_4_bits_exceptionVec_0 = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_exceptionVec_0;
        io_enq_req_4_bits_exceptionVec_1 = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_exceptionVec_1;
        io_enq_req_4_bits_exceptionVec_2 = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_exceptionVec_2;
        io_enq_req_4_bits_exceptionVec_3 = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_exceptionVec_3;
        io_enq_req_4_bits_exceptionVec_12 = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_exceptionVec_12;
        io_enq_req_4_bits_exceptionVec_20 = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_exceptionVec_20;
        io_enq_req_4_bits_exceptionVec_22 = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_exceptionVec_22;
        io_enq_req_4_bits_isFetchMalAddr = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_isFetchMalAddr;
        io_enq_req_4_bits_hasException = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_hasException;
        io_enq_req_4_bits_trigger = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_trigger;
        io_enq_req_4_bits_preDecodeInfo_isRVC = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_preDecodeInfo_isRVC;
        io_enq_req_4_bits_crossPageIPFFix = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_crossPageIPFFix;
        io_enq_req_4_bits_ftqPtr_flag = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_ftqPtr_flag;
        io_enq_req_4_bits_ftqPtr_value = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_ftqPtr_value;
        io_enq_req_4_bits_ftqOffset = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_ftqOffset;
        io_enq_req_4_bits_ldest = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_ldest;
        io_enq_req_4_bits_fuType = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_fuType;
        io_enq_req_4_bits_fuOpType = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_fuOpType;
        io_enq_req_4_bits_rfWen = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_rfWen;
        io_enq_req_4_bits_fpWen = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_fpWen;
        io_enq_req_4_bits_vecWen = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_vecWen;
        io_enq_req_4_bits_v0Wen = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_v0Wen;
        io_enq_req_4_bits_vlWen = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_vlWen;
        io_enq_req_4_bits_isXSTrap = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_isXSTrap;
        io_enq_req_4_bits_waitForward = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_waitForward;
        io_enq_req_4_bits_blockBackward = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_blockBackward;
        io_enq_req_4_bits_flushPipe = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_flushPipe;
        io_enq_req_4_bits_vpu_vill = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_vpu_vill;
        io_enq_req_4_bits_vpu_vma = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_vpu_vma;
        io_enq_req_4_bits_vpu_vta = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_vpu_vta;
        io_enq_req_4_bits_vpu_vsew = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_vpu_vsew;
        io_enq_req_4_bits_vpu_vlmul = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_vpu_vlmul;
        io_enq_req_4_bits_vpu_specVill = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_vpu_specVill;
        io_enq_req_4_bits_vpu_specVma = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_vpu_specVma;
        io_enq_req_4_bits_vpu_specVta = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_vpu_specVta;
        io_enq_req_4_bits_vpu_specVsew = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_vpu_specVsew;
        io_enq_req_4_bits_vpu_specVlmul = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_vpu_specVlmul;
        io_enq_req_4_bits_vlsInstr = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_vlsInstr;
        io_enq_req_4_bits_wfflags = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_wfflags;
        io_enq_req_4_bits_isMove = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_isMove;
        io_enq_req_4_bits_isVset = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_isVset;
        io_enq_req_4_bits_firstUop = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_firstUop;
        io_enq_req_4_bits_lastUop = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_lastUop;
        io_enq_req_4_bits_numWB = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_numWB;
        io_enq_req_4_bits_commitType = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_commitType;
        io_enq_req_4_bits_pdest = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_pdest;
        io_enq_req_4_bits_robIdx_flag = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_robIdx_flag;
        io_enq_req_4_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_robIdx_value;
        io_enq_req_4_bits_instrSize = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_instrSize;
        io_enq_req_4_bits_dirtyFs = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_dirtyFs;
        io_enq_req_4_bits_dirtyVs = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_dirtyVs;
        io_enq_req_4_bits_traceBlockInPipe_itype = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_traceBlockInPipe_itype;
        io_enq_req_4_bits_traceBlockInPipe_iretire = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_traceBlockInPipe_iretire;
        io_enq_req_4_bits_traceBlockInPipe_ilastsize = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_traceBlockInPipe_ilastsize;
        io_enq_req_4_bits_eliminatedMove = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_eliminatedMove;
        io_enq_req_4_bits_snapshot = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_snapshot;
        io_enq_req_4_bits_lqIdx_value = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_lqIdx_value;
        io_enq_req_4_bits_sqIdx_value = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_sqIdx_value;
        io_enq_req_4_bits_singleStep = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_singleStep;
        io_enq_req_4_bits_debug_sim_trig = this.vif.mon_mp.mon_cb.io_enq_req_4_bits_debug_sim_trig;
        io_enq_req_5_valid = this.vif.mon_mp.mon_cb.io_enq_req_5_valid;
        io_enq_req_5_bits_instr = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_instr;
        io_enq_req_5_bits_pc = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_pc;
        io_enq_req_5_bits_exceptionVec_0 = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_exceptionVec_0;
        io_enq_req_5_bits_exceptionVec_1 = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_exceptionVec_1;
        io_enq_req_5_bits_exceptionVec_2 = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_exceptionVec_2;
        io_enq_req_5_bits_exceptionVec_3 = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_exceptionVec_3;
        io_enq_req_5_bits_exceptionVec_12 = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_exceptionVec_12;
        io_enq_req_5_bits_exceptionVec_20 = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_exceptionVec_20;
        io_enq_req_5_bits_exceptionVec_22 = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_exceptionVec_22;
        io_enq_req_5_bits_isFetchMalAddr = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_isFetchMalAddr;
        io_enq_req_5_bits_hasException = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_hasException;
        io_enq_req_5_bits_trigger = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_trigger;
        io_enq_req_5_bits_preDecodeInfo_isRVC = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_preDecodeInfo_isRVC;
        io_enq_req_5_bits_crossPageIPFFix = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_crossPageIPFFix;
        io_enq_req_5_bits_ftqPtr_flag = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_ftqPtr_flag;
        io_enq_req_5_bits_ftqPtr_value = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_ftqPtr_value;
        io_enq_req_5_bits_ftqOffset = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_ftqOffset;
        io_enq_req_5_bits_ldest = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_ldest;
        io_enq_req_5_bits_fuType = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_fuType;
        io_enq_req_5_bits_fuOpType = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_fuOpType;
        io_enq_req_5_bits_rfWen = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_rfWen;
        io_enq_req_5_bits_fpWen = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_fpWen;
        io_enq_req_5_bits_vecWen = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_vecWen;
        io_enq_req_5_bits_v0Wen = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_v0Wen;
        io_enq_req_5_bits_vlWen = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_vlWen;
        io_enq_req_5_bits_isXSTrap = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_isXSTrap;
        io_enq_req_5_bits_waitForward = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_waitForward;
        io_enq_req_5_bits_blockBackward = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_blockBackward;
        io_enq_req_5_bits_flushPipe = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_flushPipe;
        io_enq_req_5_bits_vpu_vill = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_vpu_vill;
        io_enq_req_5_bits_vpu_vma = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_vpu_vma;
        io_enq_req_5_bits_vpu_vta = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_vpu_vta;
        io_enq_req_5_bits_vpu_vsew = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_vpu_vsew;
        io_enq_req_5_bits_vpu_vlmul = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_vpu_vlmul;
        io_enq_req_5_bits_vpu_specVill = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_vpu_specVill;
        io_enq_req_5_bits_vpu_specVma = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_vpu_specVma;
        io_enq_req_5_bits_vpu_specVta = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_vpu_specVta;
        io_enq_req_5_bits_vpu_specVsew = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_vpu_specVsew;
        io_enq_req_5_bits_vpu_specVlmul = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_vpu_specVlmul;
        io_enq_req_5_bits_vlsInstr = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_vlsInstr;
        io_enq_req_5_bits_wfflags = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_wfflags;
        io_enq_req_5_bits_isMove = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_isMove;
        io_enq_req_5_bits_isVset = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_isVset;
        io_enq_req_5_bits_firstUop = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_firstUop;
        io_enq_req_5_bits_lastUop = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_lastUop;
        io_enq_req_5_bits_numWB = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_numWB;
        io_enq_req_5_bits_commitType = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_commitType;
        io_enq_req_5_bits_pdest = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_pdest;
        io_enq_req_5_bits_robIdx_flag = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_robIdx_flag;
        io_enq_req_5_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_robIdx_value;
        io_enq_req_5_bits_instrSize = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_instrSize;
        io_enq_req_5_bits_dirtyFs = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_dirtyFs;
        io_enq_req_5_bits_dirtyVs = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_dirtyVs;
        io_enq_req_5_bits_traceBlockInPipe_itype = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_traceBlockInPipe_itype;
        io_enq_req_5_bits_traceBlockInPipe_iretire = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_traceBlockInPipe_iretire;
        io_enq_req_5_bits_traceBlockInPipe_ilastsize = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_traceBlockInPipe_ilastsize;
        io_enq_req_5_bits_eliminatedMove = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_eliminatedMove;
        io_enq_req_5_bits_snapshot = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_snapshot;
        io_enq_req_5_bits_lqIdx_value = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_lqIdx_value;
        io_enq_req_5_bits_sqIdx_value = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_sqIdx_value;
        io_enq_req_5_bits_singleStep = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_singleStep;
        io_enq_req_5_bits_debug_sim_trig = this.vif.mon_mp.mon_cb.io_enq_req_5_bits_debug_sim_trig;

        // if(this.cfg.xz_sw==tcnt_dec_base::ON & this.vif.rst_n==1'b1) begin
        //     `TCNT_CHECK_SIG_XZ(clock,clock,1);
        //     `TCNT_CHECK_SIG_XZ(reset,reset,1);
        //     `TCNT_CHECK_SIG_XZ(io_hartId,io_hartId,6);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_valid,io_enq_req_0_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_instr,io_enq_req_0_bits_instr,32);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_pc,io_enq_req_0_bits_pc,50);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_exceptionVec_0,io_enq_req_0_bits_exceptionVec_0,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_exceptionVec_1,io_enq_req_0_bits_exceptionVec_1,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_exceptionVec_2,io_enq_req_0_bits_exceptionVec_2,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_exceptionVec_3,io_enq_req_0_bits_exceptionVec_3,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_exceptionVec_12,io_enq_req_0_bits_exceptionVec_12,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_exceptionVec_20,io_enq_req_0_bits_exceptionVec_20,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_exceptionVec_22,io_enq_req_0_bits_exceptionVec_22,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_isFetchMalAddr,io_enq_req_0_bits_isFetchMalAddr,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_hasException,io_enq_req_0_bits_hasException,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_trigger,io_enq_req_0_bits_trigger,4);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_preDecodeInfo_isRVC,io_enq_req_0_bits_preDecodeInfo_isRVC,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_crossPageIPFFix,io_enq_req_0_bits_crossPageIPFFix,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_ftqPtr_flag,io_enq_req_0_bits_ftqPtr_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_ftqPtr_value,io_enq_req_0_bits_ftqPtr_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_ftqOffset,io_enq_req_0_bits_ftqOffset,4);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_ldest,io_enq_req_0_bits_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_fuType,io_enq_req_0_bits_fuType,35);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_fuOpType,io_enq_req_0_bits_fuOpType,9);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_rfWen,io_enq_req_0_bits_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_fpWen,io_enq_req_0_bits_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_vecWen,io_enq_req_0_bits_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_v0Wen,io_enq_req_0_bits_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_vlWen,io_enq_req_0_bits_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_isXSTrap,io_enq_req_0_bits_isXSTrap,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_waitForward,io_enq_req_0_bits_waitForward,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_blockBackward,io_enq_req_0_bits_blockBackward,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_flushPipe,io_enq_req_0_bits_flushPipe,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_vpu_vill,io_enq_req_0_bits_vpu_vill,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_vpu_vma,io_enq_req_0_bits_vpu_vma,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_vpu_vta,io_enq_req_0_bits_vpu_vta,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_vpu_vsew,io_enq_req_0_bits_vpu_vsew,2);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_vpu_vlmul,io_enq_req_0_bits_vpu_vlmul,3);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_vpu_specVill,io_enq_req_0_bits_vpu_specVill,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_vpu_specVma,io_enq_req_0_bits_vpu_specVma,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_vpu_specVta,io_enq_req_0_bits_vpu_specVta,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_vpu_specVsew,io_enq_req_0_bits_vpu_specVsew,2);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_vpu_specVlmul,io_enq_req_0_bits_vpu_specVlmul,3);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_vlsInstr,io_enq_req_0_bits_vlsInstr,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_wfflags,io_enq_req_0_bits_wfflags,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_isMove,io_enq_req_0_bits_isMove,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_isVset,io_enq_req_0_bits_isVset,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_firstUop,io_enq_req_0_bits_firstUop,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_lastUop,io_enq_req_0_bits_lastUop,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_numWB,io_enq_req_0_bits_numWB,7);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_commitType,io_enq_req_0_bits_commitType,3);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_pdest,io_enq_req_0_bits_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_robIdx_flag,io_enq_req_0_bits_robIdx_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_robIdx_value,io_enq_req_0_bits_robIdx_value,8);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_instrSize,io_enq_req_0_bits_instrSize,3);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_dirtyFs,io_enq_req_0_bits_dirtyFs,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_dirtyVs,io_enq_req_0_bits_dirtyVs,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_traceBlockInPipe_itype,io_enq_req_0_bits_traceBlockInPipe_itype,4);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_traceBlockInPipe_iretire,io_enq_req_0_bits_traceBlockInPipe_iretire,4);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_traceBlockInPipe_ilastsize,io_enq_req_0_bits_traceBlockInPipe_ilastsize,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_eliminatedMove,io_enq_req_0_bits_eliminatedMove,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_snapshot,io_enq_req_0_bits_snapshot,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_lqIdx_value,io_enq_req_0_bits_lqIdx_value,7);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_sqIdx_value,io_enq_req_0_bits_sqIdx_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_singleStep,io_enq_req_0_bits_singleStep,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_0_bits_debug_sim_trig,io_enq_req_0_bits_debug_sim_trig,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_valid,io_enq_req_1_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_instr,io_enq_req_1_bits_instr,32);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_pc,io_enq_req_1_bits_pc,50);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_exceptionVec_0,io_enq_req_1_bits_exceptionVec_0,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_exceptionVec_1,io_enq_req_1_bits_exceptionVec_1,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_exceptionVec_2,io_enq_req_1_bits_exceptionVec_2,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_exceptionVec_3,io_enq_req_1_bits_exceptionVec_3,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_exceptionVec_12,io_enq_req_1_bits_exceptionVec_12,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_exceptionVec_20,io_enq_req_1_bits_exceptionVec_20,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_exceptionVec_22,io_enq_req_1_bits_exceptionVec_22,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_isFetchMalAddr,io_enq_req_1_bits_isFetchMalAddr,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_hasException,io_enq_req_1_bits_hasException,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_trigger,io_enq_req_1_bits_trigger,4);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_preDecodeInfo_isRVC,io_enq_req_1_bits_preDecodeInfo_isRVC,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_crossPageIPFFix,io_enq_req_1_bits_crossPageIPFFix,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_ftqPtr_flag,io_enq_req_1_bits_ftqPtr_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_ftqPtr_value,io_enq_req_1_bits_ftqPtr_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_ftqOffset,io_enq_req_1_bits_ftqOffset,4);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_ldest,io_enq_req_1_bits_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_fuType,io_enq_req_1_bits_fuType,35);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_fuOpType,io_enq_req_1_bits_fuOpType,9);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_rfWen,io_enq_req_1_bits_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_fpWen,io_enq_req_1_bits_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_vecWen,io_enq_req_1_bits_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_v0Wen,io_enq_req_1_bits_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_vlWen,io_enq_req_1_bits_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_isXSTrap,io_enq_req_1_bits_isXSTrap,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_waitForward,io_enq_req_1_bits_waitForward,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_blockBackward,io_enq_req_1_bits_blockBackward,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_flushPipe,io_enq_req_1_bits_flushPipe,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_vpu_vill,io_enq_req_1_bits_vpu_vill,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_vpu_vma,io_enq_req_1_bits_vpu_vma,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_vpu_vta,io_enq_req_1_bits_vpu_vta,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_vpu_vsew,io_enq_req_1_bits_vpu_vsew,2);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_vpu_vlmul,io_enq_req_1_bits_vpu_vlmul,3);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_vpu_specVill,io_enq_req_1_bits_vpu_specVill,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_vpu_specVma,io_enq_req_1_bits_vpu_specVma,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_vpu_specVta,io_enq_req_1_bits_vpu_specVta,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_vpu_specVsew,io_enq_req_1_bits_vpu_specVsew,2);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_vpu_specVlmul,io_enq_req_1_bits_vpu_specVlmul,3);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_vlsInstr,io_enq_req_1_bits_vlsInstr,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_wfflags,io_enq_req_1_bits_wfflags,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_isMove,io_enq_req_1_bits_isMove,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_isVset,io_enq_req_1_bits_isVset,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_firstUop,io_enq_req_1_bits_firstUop,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_lastUop,io_enq_req_1_bits_lastUop,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_numWB,io_enq_req_1_bits_numWB,7);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_commitType,io_enq_req_1_bits_commitType,3);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_pdest,io_enq_req_1_bits_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_robIdx_flag,io_enq_req_1_bits_robIdx_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_robIdx_value,io_enq_req_1_bits_robIdx_value,8);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_instrSize,io_enq_req_1_bits_instrSize,3);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_dirtyFs,io_enq_req_1_bits_dirtyFs,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_dirtyVs,io_enq_req_1_bits_dirtyVs,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_traceBlockInPipe_itype,io_enq_req_1_bits_traceBlockInPipe_itype,4);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_traceBlockInPipe_iretire,io_enq_req_1_bits_traceBlockInPipe_iretire,4);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_traceBlockInPipe_ilastsize,io_enq_req_1_bits_traceBlockInPipe_ilastsize,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_eliminatedMove,io_enq_req_1_bits_eliminatedMove,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_snapshot,io_enq_req_1_bits_snapshot,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_lqIdx_value,io_enq_req_1_bits_lqIdx_value,7);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_sqIdx_value,io_enq_req_1_bits_sqIdx_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_singleStep,io_enq_req_1_bits_singleStep,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_1_bits_debug_sim_trig,io_enq_req_1_bits_debug_sim_trig,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_valid,io_enq_req_2_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_instr,io_enq_req_2_bits_instr,32);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_pc,io_enq_req_2_bits_pc,50);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_exceptionVec_0,io_enq_req_2_bits_exceptionVec_0,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_exceptionVec_1,io_enq_req_2_bits_exceptionVec_1,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_exceptionVec_2,io_enq_req_2_bits_exceptionVec_2,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_exceptionVec_3,io_enq_req_2_bits_exceptionVec_3,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_exceptionVec_12,io_enq_req_2_bits_exceptionVec_12,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_exceptionVec_20,io_enq_req_2_bits_exceptionVec_20,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_exceptionVec_22,io_enq_req_2_bits_exceptionVec_22,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_isFetchMalAddr,io_enq_req_2_bits_isFetchMalAddr,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_hasException,io_enq_req_2_bits_hasException,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_trigger,io_enq_req_2_bits_trigger,4);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_preDecodeInfo_isRVC,io_enq_req_2_bits_preDecodeInfo_isRVC,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_crossPageIPFFix,io_enq_req_2_bits_crossPageIPFFix,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_ftqPtr_flag,io_enq_req_2_bits_ftqPtr_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_ftqPtr_value,io_enq_req_2_bits_ftqPtr_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_ftqOffset,io_enq_req_2_bits_ftqOffset,4);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_ldest,io_enq_req_2_bits_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_fuType,io_enq_req_2_bits_fuType,35);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_fuOpType,io_enq_req_2_bits_fuOpType,9);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_rfWen,io_enq_req_2_bits_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_fpWen,io_enq_req_2_bits_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_vecWen,io_enq_req_2_bits_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_v0Wen,io_enq_req_2_bits_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_vlWen,io_enq_req_2_bits_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_isXSTrap,io_enq_req_2_bits_isXSTrap,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_waitForward,io_enq_req_2_bits_waitForward,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_blockBackward,io_enq_req_2_bits_blockBackward,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_flushPipe,io_enq_req_2_bits_flushPipe,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_vpu_vill,io_enq_req_2_bits_vpu_vill,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_vpu_vma,io_enq_req_2_bits_vpu_vma,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_vpu_vta,io_enq_req_2_bits_vpu_vta,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_vpu_vsew,io_enq_req_2_bits_vpu_vsew,2);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_vpu_vlmul,io_enq_req_2_bits_vpu_vlmul,3);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_vpu_specVill,io_enq_req_2_bits_vpu_specVill,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_vpu_specVma,io_enq_req_2_bits_vpu_specVma,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_vpu_specVta,io_enq_req_2_bits_vpu_specVta,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_vpu_specVsew,io_enq_req_2_bits_vpu_specVsew,2);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_vpu_specVlmul,io_enq_req_2_bits_vpu_specVlmul,3);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_vlsInstr,io_enq_req_2_bits_vlsInstr,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_wfflags,io_enq_req_2_bits_wfflags,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_isMove,io_enq_req_2_bits_isMove,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_isVset,io_enq_req_2_bits_isVset,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_firstUop,io_enq_req_2_bits_firstUop,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_lastUop,io_enq_req_2_bits_lastUop,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_numWB,io_enq_req_2_bits_numWB,7);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_commitType,io_enq_req_2_bits_commitType,3);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_pdest,io_enq_req_2_bits_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_robIdx_flag,io_enq_req_2_bits_robIdx_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_robIdx_value,io_enq_req_2_bits_robIdx_value,8);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_instrSize,io_enq_req_2_bits_instrSize,3);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_dirtyFs,io_enq_req_2_bits_dirtyFs,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_dirtyVs,io_enq_req_2_bits_dirtyVs,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_traceBlockInPipe_itype,io_enq_req_2_bits_traceBlockInPipe_itype,4);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_traceBlockInPipe_iretire,io_enq_req_2_bits_traceBlockInPipe_iretire,4);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_traceBlockInPipe_ilastsize,io_enq_req_2_bits_traceBlockInPipe_ilastsize,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_eliminatedMove,io_enq_req_2_bits_eliminatedMove,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_snapshot,io_enq_req_2_bits_snapshot,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_lqIdx_value,io_enq_req_2_bits_lqIdx_value,7);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_sqIdx_value,io_enq_req_2_bits_sqIdx_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_singleStep,io_enq_req_2_bits_singleStep,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_2_bits_debug_sim_trig,io_enq_req_2_bits_debug_sim_trig,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_valid,io_enq_req_3_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_instr,io_enq_req_3_bits_instr,32);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_pc,io_enq_req_3_bits_pc,50);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_exceptionVec_0,io_enq_req_3_bits_exceptionVec_0,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_exceptionVec_1,io_enq_req_3_bits_exceptionVec_1,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_exceptionVec_2,io_enq_req_3_bits_exceptionVec_2,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_exceptionVec_3,io_enq_req_3_bits_exceptionVec_3,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_exceptionVec_12,io_enq_req_3_bits_exceptionVec_12,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_exceptionVec_20,io_enq_req_3_bits_exceptionVec_20,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_exceptionVec_22,io_enq_req_3_bits_exceptionVec_22,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_isFetchMalAddr,io_enq_req_3_bits_isFetchMalAddr,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_hasException,io_enq_req_3_bits_hasException,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_trigger,io_enq_req_3_bits_trigger,4);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_preDecodeInfo_isRVC,io_enq_req_3_bits_preDecodeInfo_isRVC,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_crossPageIPFFix,io_enq_req_3_bits_crossPageIPFFix,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_ftqPtr_flag,io_enq_req_3_bits_ftqPtr_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_ftqPtr_value,io_enq_req_3_bits_ftqPtr_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_ftqOffset,io_enq_req_3_bits_ftqOffset,4);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_ldest,io_enq_req_3_bits_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_fuType,io_enq_req_3_bits_fuType,35);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_fuOpType,io_enq_req_3_bits_fuOpType,9);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_rfWen,io_enq_req_3_bits_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_fpWen,io_enq_req_3_bits_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_vecWen,io_enq_req_3_bits_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_v0Wen,io_enq_req_3_bits_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_vlWen,io_enq_req_3_bits_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_isXSTrap,io_enq_req_3_bits_isXSTrap,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_waitForward,io_enq_req_3_bits_waitForward,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_blockBackward,io_enq_req_3_bits_blockBackward,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_flushPipe,io_enq_req_3_bits_flushPipe,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_vpu_vill,io_enq_req_3_bits_vpu_vill,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_vpu_vma,io_enq_req_3_bits_vpu_vma,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_vpu_vta,io_enq_req_3_bits_vpu_vta,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_vpu_vsew,io_enq_req_3_bits_vpu_vsew,2);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_vpu_vlmul,io_enq_req_3_bits_vpu_vlmul,3);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_vpu_specVill,io_enq_req_3_bits_vpu_specVill,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_vpu_specVma,io_enq_req_3_bits_vpu_specVma,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_vpu_specVta,io_enq_req_3_bits_vpu_specVta,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_vpu_specVsew,io_enq_req_3_bits_vpu_specVsew,2);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_vpu_specVlmul,io_enq_req_3_bits_vpu_specVlmul,3);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_vlsInstr,io_enq_req_3_bits_vlsInstr,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_wfflags,io_enq_req_3_bits_wfflags,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_isMove,io_enq_req_3_bits_isMove,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_isVset,io_enq_req_3_bits_isVset,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_firstUop,io_enq_req_3_bits_firstUop,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_lastUop,io_enq_req_3_bits_lastUop,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_numWB,io_enq_req_3_bits_numWB,7);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_commitType,io_enq_req_3_bits_commitType,3);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_pdest,io_enq_req_3_bits_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_robIdx_flag,io_enq_req_3_bits_robIdx_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_robIdx_value,io_enq_req_3_bits_robIdx_value,8);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_instrSize,io_enq_req_3_bits_instrSize,3);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_dirtyFs,io_enq_req_3_bits_dirtyFs,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_dirtyVs,io_enq_req_3_bits_dirtyVs,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_traceBlockInPipe_itype,io_enq_req_3_bits_traceBlockInPipe_itype,4);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_traceBlockInPipe_iretire,io_enq_req_3_bits_traceBlockInPipe_iretire,4);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_traceBlockInPipe_ilastsize,io_enq_req_3_bits_traceBlockInPipe_ilastsize,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_eliminatedMove,io_enq_req_3_bits_eliminatedMove,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_snapshot,io_enq_req_3_bits_snapshot,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_lqIdx_value,io_enq_req_3_bits_lqIdx_value,7);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_sqIdx_value,io_enq_req_3_bits_sqIdx_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_singleStep,io_enq_req_3_bits_singleStep,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_3_bits_debug_sim_trig,io_enq_req_3_bits_debug_sim_trig,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_valid,io_enq_req_4_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_instr,io_enq_req_4_bits_instr,32);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_pc,io_enq_req_4_bits_pc,50);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_exceptionVec_0,io_enq_req_4_bits_exceptionVec_0,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_exceptionVec_1,io_enq_req_4_bits_exceptionVec_1,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_exceptionVec_2,io_enq_req_4_bits_exceptionVec_2,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_exceptionVec_3,io_enq_req_4_bits_exceptionVec_3,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_exceptionVec_12,io_enq_req_4_bits_exceptionVec_12,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_exceptionVec_20,io_enq_req_4_bits_exceptionVec_20,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_exceptionVec_22,io_enq_req_4_bits_exceptionVec_22,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_isFetchMalAddr,io_enq_req_4_bits_isFetchMalAddr,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_hasException,io_enq_req_4_bits_hasException,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_trigger,io_enq_req_4_bits_trigger,4);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_preDecodeInfo_isRVC,io_enq_req_4_bits_preDecodeInfo_isRVC,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_crossPageIPFFix,io_enq_req_4_bits_crossPageIPFFix,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_ftqPtr_flag,io_enq_req_4_bits_ftqPtr_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_ftqPtr_value,io_enq_req_4_bits_ftqPtr_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_ftqOffset,io_enq_req_4_bits_ftqOffset,4);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_ldest,io_enq_req_4_bits_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_fuType,io_enq_req_4_bits_fuType,35);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_fuOpType,io_enq_req_4_bits_fuOpType,9);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_rfWen,io_enq_req_4_bits_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_fpWen,io_enq_req_4_bits_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_vecWen,io_enq_req_4_bits_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_v0Wen,io_enq_req_4_bits_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_vlWen,io_enq_req_4_bits_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_isXSTrap,io_enq_req_4_bits_isXSTrap,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_waitForward,io_enq_req_4_bits_waitForward,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_blockBackward,io_enq_req_4_bits_blockBackward,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_flushPipe,io_enq_req_4_bits_flushPipe,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_vpu_vill,io_enq_req_4_bits_vpu_vill,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_vpu_vma,io_enq_req_4_bits_vpu_vma,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_vpu_vta,io_enq_req_4_bits_vpu_vta,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_vpu_vsew,io_enq_req_4_bits_vpu_vsew,2);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_vpu_vlmul,io_enq_req_4_bits_vpu_vlmul,3);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_vpu_specVill,io_enq_req_4_bits_vpu_specVill,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_vpu_specVma,io_enq_req_4_bits_vpu_specVma,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_vpu_specVta,io_enq_req_4_bits_vpu_specVta,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_vpu_specVsew,io_enq_req_4_bits_vpu_specVsew,2);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_vpu_specVlmul,io_enq_req_4_bits_vpu_specVlmul,3);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_vlsInstr,io_enq_req_4_bits_vlsInstr,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_wfflags,io_enq_req_4_bits_wfflags,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_isMove,io_enq_req_4_bits_isMove,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_isVset,io_enq_req_4_bits_isVset,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_firstUop,io_enq_req_4_bits_firstUop,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_lastUop,io_enq_req_4_bits_lastUop,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_numWB,io_enq_req_4_bits_numWB,7);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_commitType,io_enq_req_4_bits_commitType,3);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_pdest,io_enq_req_4_bits_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_robIdx_flag,io_enq_req_4_bits_robIdx_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_robIdx_value,io_enq_req_4_bits_robIdx_value,8);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_instrSize,io_enq_req_4_bits_instrSize,3);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_dirtyFs,io_enq_req_4_bits_dirtyFs,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_dirtyVs,io_enq_req_4_bits_dirtyVs,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_traceBlockInPipe_itype,io_enq_req_4_bits_traceBlockInPipe_itype,4);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_traceBlockInPipe_iretire,io_enq_req_4_bits_traceBlockInPipe_iretire,4);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_traceBlockInPipe_ilastsize,io_enq_req_4_bits_traceBlockInPipe_ilastsize,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_eliminatedMove,io_enq_req_4_bits_eliminatedMove,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_snapshot,io_enq_req_4_bits_snapshot,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_lqIdx_value,io_enq_req_4_bits_lqIdx_value,7);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_sqIdx_value,io_enq_req_4_bits_sqIdx_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_singleStep,io_enq_req_4_bits_singleStep,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_4_bits_debug_sim_trig,io_enq_req_4_bits_debug_sim_trig,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_valid,io_enq_req_5_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_instr,io_enq_req_5_bits_instr,32);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_pc,io_enq_req_5_bits_pc,50);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_exceptionVec_0,io_enq_req_5_bits_exceptionVec_0,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_exceptionVec_1,io_enq_req_5_bits_exceptionVec_1,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_exceptionVec_2,io_enq_req_5_bits_exceptionVec_2,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_exceptionVec_3,io_enq_req_5_bits_exceptionVec_3,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_exceptionVec_12,io_enq_req_5_bits_exceptionVec_12,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_exceptionVec_20,io_enq_req_5_bits_exceptionVec_20,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_exceptionVec_22,io_enq_req_5_bits_exceptionVec_22,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_isFetchMalAddr,io_enq_req_5_bits_isFetchMalAddr,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_hasException,io_enq_req_5_bits_hasException,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_trigger,io_enq_req_5_bits_trigger,4);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_preDecodeInfo_isRVC,io_enq_req_5_bits_preDecodeInfo_isRVC,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_crossPageIPFFix,io_enq_req_5_bits_crossPageIPFFix,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_ftqPtr_flag,io_enq_req_5_bits_ftqPtr_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_ftqPtr_value,io_enq_req_5_bits_ftqPtr_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_ftqOffset,io_enq_req_5_bits_ftqOffset,4);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_ldest,io_enq_req_5_bits_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_fuType,io_enq_req_5_bits_fuType,35);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_fuOpType,io_enq_req_5_bits_fuOpType,9);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_rfWen,io_enq_req_5_bits_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_fpWen,io_enq_req_5_bits_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_vecWen,io_enq_req_5_bits_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_v0Wen,io_enq_req_5_bits_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_vlWen,io_enq_req_5_bits_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_isXSTrap,io_enq_req_5_bits_isXSTrap,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_waitForward,io_enq_req_5_bits_waitForward,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_blockBackward,io_enq_req_5_bits_blockBackward,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_flushPipe,io_enq_req_5_bits_flushPipe,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_vpu_vill,io_enq_req_5_bits_vpu_vill,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_vpu_vma,io_enq_req_5_bits_vpu_vma,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_vpu_vta,io_enq_req_5_bits_vpu_vta,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_vpu_vsew,io_enq_req_5_bits_vpu_vsew,2);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_vpu_vlmul,io_enq_req_5_bits_vpu_vlmul,3);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_vpu_specVill,io_enq_req_5_bits_vpu_specVill,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_vpu_specVma,io_enq_req_5_bits_vpu_specVma,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_vpu_specVta,io_enq_req_5_bits_vpu_specVta,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_vpu_specVsew,io_enq_req_5_bits_vpu_specVsew,2);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_vpu_specVlmul,io_enq_req_5_bits_vpu_specVlmul,3);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_vlsInstr,io_enq_req_5_bits_vlsInstr,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_wfflags,io_enq_req_5_bits_wfflags,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_isMove,io_enq_req_5_bits_isMove,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_isVset,io_enq_req_5_bits_isVset,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_firstUop,io_enq_req_5_bits_firstUop,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_lastUop,io_enq_req_5_bits_lastUop,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_numWB,io_enq_req_5_bits_numWB,7);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_commitType,io_enq_req_5_bits_commitType,3);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_pdest,io_enq_req_5_bits_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_robIdx_flag,io_enq_req_5_bits_robIdx_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_robIdx_value,io_enq_req_5_bits_robIdx_value,8);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_instrSize,io_enq_req_5_bits_instrSize,3);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_dirtyFs,io_enq_req_5_bits_dirtyFs,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_dirtyVs,io_enq_req_5_bits_dirtyVs,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_traceBlockInPipe_itype,io_enq_req_5_bits_traceBlockInPipe_itype,4);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_traceBlockInPipe_iretire,io_enq_req_5_bits_traceBlockInPipe_iretire,4);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_traceBlockInPipe_ilastsize,io_enq_req_5_bits_traceBlockInPipe_ilastsize,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_eliminatedMove,io_enq_req_5_bits_eliminatedMove,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_snapshot,io_enq_req_5_bits_snapshot,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_lqIdx_value,io_enq_req_5_bits_lqIdx_value,7);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_sqIdx_value,io_enq_req_5_bits_sqIdx_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_singleStep,io_enq_req_5_bits_singleStep,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_req_5_bits_debug_sim_trig,io_enq_req_5_bits_debug_sim_trig,1);

        //end
        //if(xxxTODOxxx==1'b1) begin
        //    mon_tr = rename_in_agent_xaction::type_id::create("mon_tr");
        //    mon_tr.clock = clock;
        //    mon_tr.reset = reset;
        //    mon_tr.io_hartId = io_hartId;
        //    mon_tr.io_enq_req_0_valid = io_enq_req_0_valid;
        //    mon_tr.io_enq_req_0_bits_instr = io_enq_req_0_bits_instr;
        //    mon_tr.io_enq_req_0_bits_pc = io_enq_req_0_bits_pc;
        //    mon_tr.io_enq_req_0_bits_exceptionVec_0 = io_enq_req_0_bits_exceptionVec_0;
        //    mon_tr.io_enq_req_0_bits_exceptionVec_1 = io_enq_req_0_bits_exceptionVec_1;
        //    mon_tr.io_enq_req_0_bits_exceptionVec_2 = io_enq_req_0_bits_exceptionVec_2;
        //    mon_tr.io_enq_req_0_bits_exceptionVec_3 = io_enq_req_0_bits_exceptionVec_3;
        //    mon_tr.io_enq_req_0_bits_exceptionVec_12 = io_enq_req_0_bits_exceptionVec_12;
        //    mon_tr.io_enq_req_0_bits_exceptionVec_20 = io_enq_req_0_bits_exceptionVec_20;
        //    mon_tr.io_enq_req_0_bits_exceptionVec_22 = io_enq_req_0_bits_exceptionVec_22;
        //    mon_tr.io_enq_req_0_bits_isFetchMalAddr = io_enq_req_0_bits_isFetchMalAddr;
        //    mon_tr.io_enq_req_0_bits_hasException = io_enq_req_0_bits_hasException;
        //    mon_tr.io_enq_req_0_bits_trigger = io_enq_req_0_bits_trigger;
        //    mon_tr.io_enq_req_0_bits_preDecodeInfo_isRVC = io_enq_req_0_bits_preDecodeInfo_isRVC;
        //    mon_tr.io_enq_req_0_bits_crossPageIPFFix = io_enq_req_0_bits_crossPageIPFFix;
        //    mon_tr.io_enq_req_0_bits_ftqPtr_flag = io_enq_req_0_bits_ftqPtr_flag;
        //    mon_tr.io_enq_req_0_bits_ftqPtr_value = io_enq_req_0_bits_ftqPtr_value;
        //    mon_tr.io_enq_req_0_bits_ftqOffset = io_enq_req_0_bits_ftqOffset;
        //    mon_tr.io_enq_req_0_bits_ldest = io_enq_req_0_bits_ldest;
        //    mon_tr.io_enq_req_0_bits_fuType = io_enq_req_0_bits_fuType;
        //    mon_tr.io_enq_req_0_bits_fuOpType = io_enq_req_0_bits_fuOpType;
        //    mon_tr.io_enq_req_0_bits_rfWen = io_enq_req_0_bits_rfWen;
        //    mon_tr.io_enq_req_0_bits_fpWen = io_enq_req_0_bits_fpWen;
        //    mon_tr.io_enq_req_0_bits_vecWen = io_enq_req_0_bits_vecWen;
        //    mon_tr.io_enq_req_0_bits_v0Wen = io_enq_req_0_bits_v0Wen;
        //    mon_tr.io_enq_req_0_bits_vlWen = io_enq_req_0_bits_vlWen;
        //    mon_tr.io_enq_req_0_bits_isXSTrap = io_enq_req_0_bits_isXSTrap;
        //    mon_tr.io_enq_req_0_bits_waitForward = io_enq_req_0_bits_waitForward;
        //    mon_tr.io_enq_req_0_bits_blockBackward = io_enq_req_0_bits_blockBackward;
        //    mon_tr.io_enq_req_0_bits_flushPipe = io_enq_req_0_bits_flushPipe;
        //    mon_tr.io_enq_req_0_bits_vpu_vill = io_enq_req_0_bits_vpu_vill;
        //    mon_tr.io_enq_req_0_bits_vpu_vma = io_enq_req_0_bits_vpu_vma;
        //    mon_tr.io_enq_req_0_bits_vpu_vta = io_enq_req_0_bits_vpu_vta;
        //    mon_tr.io_enq_req_0_bits_vpu_vsew = io_enq_req_0_bits_vpu_vsew;
        //    mon_tr.io_enq_req_0_bits_vpu_vlmul = io_enq_req_0_bits_vpu_vlmul;
        //    mon_tr.io_enq_req_0_bits_vpu_specVill = io_enq_req_0_bits_vpu_specVill;
        //    mon_tr.io_enq_req_0_bits_vpu_specVma = io_enq_req_0_bits_vpu_specVma;
        //    mon_tr.io_enq_req_0_bits_vpu_specVta = io_enq_req_0_bits_vpu_specVta;
        //    mon_tr.io_enq_req_0_bits_vpu_specVsew = io_enq_req_0_bits_vpu_specVsew;
        //    mon_tr.io_enq_req_0_bits_vpu_specVlmul = io_enq_req_0_bits_vpu_specVlmul;
        //    mon_tr.io_enq_req_0_bits_vlsInstr = io_enq_req_0_bits_vlsInstr;
        //    mon_tr.io_enq_req_0_bits_wfflags = io_enq_req_0_bits_wfflags;
        //    mon_tr.io_enq_req_0_bits_isMove = io_enq_req_0_bits_isMove;
        //    mon_tr.io_enq_req_0_bits_isVset = io_enq_req_0_bits_isVset;
        //    mon_tr.io_enq_req_0_bits_firstUop = io_enq_req_0_bits_firstUop;
        //    mon_tr.io_enq_req_0_bits_lastUop = io_enq_req_0_bits_lastUop;
        //    mon_tr.io_enq_req_0_bits_numWB = io_enq_req_0_bits_numWB;
        //    mon_tr.io_enq_req_0_bits_commitType = io_enq_req_0_bits_commitType;
        //    mon_tr.io_enq_req_0_bits_pdest = io_enq_req_0_bits_pdest;
        //    mon_tr.io_enq_req_0_bits_robIdx_flag = io_enq_req_0_bits_robIdx_flag;
        //    mon_tr.io_enq_req_0_bits_robIdx_value = io_enq_req_0_bits_robIdx_value;
        //    mon_tr.io_enq_req_0_bits_instrSize = io_enq_req_0_bits_instrSize;
        //    mon_tr.io_enq_req_0_bits_dirtyFs = io_enq_req_0_bits_dirtyFs;
        //    mon_tr.io_enq_req_0_bits_dirtyVs = io_enq_req_0_bits_dirtyVs;
        //    mon_tr.io_enq_req_0_bits_traceBlockInPipe_itype = io_enq_req_0_bits_traceBlockInPipe_itype;
        //    mon_tr.io_enq_req_0_bits_traceBlockInPipe_iretire = io_enq_req_0_bits_traceBlockInPipe_iretire;
        //    mon_tr.io_enq_req_0_bits_traceBlockInPipe_ilastsize = io_enq_req_0_bits_traceBlockInPipe_ilastsize;
        //    mon_tr.io_enq_req_0_bits_eliminatedMove = io_enq_req_0_bits_eliminatedMove;
        //    mon_tr.io_enq_req_0_bits_snapshot = io_enq_req_0_bits_snapshot;
        //    mon_tr.io_enq_req_0_bits_lqIdx_value = io_enq_req_0_bits_lqIdx_value;
        //    mon_tr.io_enq_req_0_bits_sqIdx_value = io_enq_req_0_bits_sqIdx_value;
        //    mon_tr.io_enq_req_0_bits_singleStep = io_enq_req_0_bits_singleStep;
        //    mon_tr.io_enq_req_0_bits_debug_sim_trig = io_enq_req_0_bits_debug_sim_trig;
        //    mon_tr.io_enq_req_1_valid = io_enq_req_1_valid;
        //    mon_tr.io_enq_req_1_bits_instr = io_enq_req_1_bits_instr;
        //    mon_tr.io_enq_req_1_bits_pc = io_enq_req_1_bits_pc;
        //    mon_tr.io_enq_req_1_bits_exceptionVec_0 = io_enq_req_1_bits_exceptionVec_0;
        //    mon_tr.io_enq_req_1_bits_exceptionVec_1 = io_enq_req_1_bits_exceptionVec_1;
        //    mon_tr.io_enq_req_1_bits_exceptionVec_2 = io_enq_req_1_bits_exceptionVec_2;
        //    mon_tr.io_enq_req_1_bits_exceptionVec_3 = io_enq_req_1_bits_exceptionVec_3;
        //    mon_tr.io_enq_req_1_bits_exceptionVec_12 = io_enq_req_1_bits_exceptionVec_12;
        //    mon_tr.io_enq_req_1_bits_exceptionVec_20 = io_enq_req_1_bits_exceptionVec_20;
        //    mon_tr.io_enq_req_1_bits_exceptionVec_22 = io_enq_req_1_bits_exceptionVec_22;
        //    mon_tr.io_enq_req_1_bits_isFetchMalAddr = io_enq_req_1_bits_isFetchMalAddr;
        //    mon_tr.io_enq_req_1_bits_hasException = io_enq_req_1_bits_hasException;
        //    mon_tr.io_enq_req_1_bits_trigger = io_enq_req_1_bits_trigger;
        //    mon_tr.io_enq_req_1_bits_preDecodeInfo_isRVC = io_enq_req_1_bits_preDecodeInfo_isRVC;
        //    mon_tr.io_enq_req_1_bits_crossPageIPFFix = io_enq_req_1_bits_crossPageIPFFix;
        //    mon_tr.io_enq_req_1_bits_ftqPtr_flag = io_enq_req_1_bits_ftqPtr_flag;
        //    mon_tr.io_enq_req_1_bits_ftqPtr_value = io_enq_req_1_bits_ftqPtr_value;
        //    mon_tr.io_enq_req_1_bits_ftqOffset = io_enq_req_1_bits_ftqOffset;
        //    mon_tr.io_enq_req_1_bits_ldest = io_enq_req_1_bits_ldest;
        //    mon_tr.io_enq_req_1_bits_fuType = io_enq_req_1_bits_fuType;
        //    mon_tr.io_enq_req_1_bits_fuOpType = io_enq_req_1_bits_fuOpType;
        //    mon_tr.io_enq_req_1_bits_rfWen = io_enq_req_1_bits_rfWen;
        //    mon_tr.io_enq_req_1_bits_fpWen = io_enq_req_1_bits_fpWen;
        //    mon_tr.io_enq_req_1_bits_vecWen = io_enq_req_1_bits_vecWen;
        //    mon_tr.io_enq_req_1_bits_v0Wen = io_enq_req_1_bits_v0Wen;
        //    mon_tr.io_enq_req_1_bits_vlWen = io_enq_req_1_bits_vlWen;
        //    mon_tr.io_enq_req_1_bits_isXSTrap = io_enq_req_1_bits_isXSTrap;
        //    mon_tr.io_enq_req_1_bits_waitForward = io_enq_req_1_bits_waitForward;
        //    mon_tr.io_enq_req_1_bits_blockBackward = io_enq_req_1_bits_blockBackward;
        //    mon_tr.io_enq_req_1_bits_flushPipe = io_enq_req_1_bits_flushPipe;
        //    mon_tr.io_enq_req_1_bits_vpu_vill = io_enq_req_1_bits_vpu_vill;
        //    mon_tr.io_enq_req_1_bits_vpu_vma = io_enq_req_1_bits_vpu_vma;
        //    mon_tr.io_enq_req_1_bits_vpu_vta = io_enq_req_1_bits_vpu_vta;
        //    mon_tr.io_enq_req_1_bits_vpu_vsew = io_enq_req_1_bits_vpu_vsew;
        //    mon_tr.io_enq_req_1_bits_vpu_vlmul = io_enq_req_1_bits_vpu_vlmul;
        //    mon_tr.io_enq_req_1_bits_vpu_specVill = io_enq_req_1_bits_vpu_specVill;
        //    mon_tr.io_enq_req_1_bits_vpu_specVma = io_enq_req_1_bits_vpu_specVma;
        //    mon_tr.io_enq_req_1_bits_vpu_specVta = io_enq_req_1_bits_vpu_specVta;
        //    mon_tr.io_enq_req_1_bits_vpu_specVsew = io_enq_req_1_bits_vpu_specVsew;
        //    mon_tr.io_enq_req_1_bits_vpu_specVlmul = io_enq_req_1_bits_vpu_specVlmul;
        //    mon_tr.io_enq_req_1_bits_vlsInstr = io_enq_req_1_bits_vlsInstr;
        //    mon_tr.io_enq_req_1_bits_wfflags = io_enq_req_1_bits_wfflags;
        //    mon_tr.io_enq_req_1_bits_isMove = io_enq_req_1_bits_isMove;
        //    mon_tr.io_enq_req_1_bits_isVset = io_enq_req_1_bits_isVset;
        //    mon_tr.io_enq_req_1_bits_firstUop = io_enq_req_1_bits_firstUop;
        //    mon_tr.io_enq_req_1_bits_lastUop = io_enq_req_1_bits_lastUop;
        //    mon_tr.io_enq_req_1_bits_numWB = io_enq_req_1_bits_numWB;
        //    mon_tr.io_enq_req_1_bits_commitType = io_enq_req_1_bits_commitType;
        //    mon_tr.io_enq_req_1_bits_pdest = io_enq_req_1_bits_pdest;
        //    mon_tr.io_enq_req_1_bits_robIdx_flag = io_enq_req_1_bits_robIdx_flag;
        //    mon_tr.io_enq_req_1_bits_robIdx_value = io_enq_req_1_bits_robIdx_value;
        //    mon_tr.io_enq_req_1_bits_instrSize = io_enq_req_1_bits_instrSize;
        //    mon_tr.io_enq_req_1_bits_dirtyFs = io_enq_req_1_bits_dirtyFs;
        //    mon_tr.io_enq_req_1_bits_dirtyVs = io_enq_req_1_bits_dirtyVs;
        //    mon_tr.io_enq_req_1_bits_traceBlockInPipe_itype = io_enq_req_1_bits_traceBlockInPipe_itype;
        //    mon_tr.io_enq_req_1_bits_traceBlockInPipe_iretire = io_enq_req_1_bits_traceBlockInPipe_iretire;
        //    mon_tr.io_enq_req_1_bits_traceBlockInPipe_ilastsize = io_enq_req_1_bits_traceBlockInPipe_ilastsize;
        //    mon_tr.io_enq_req_1_bits_eliminatedMove = io_enq_req_1_bits_eliminatedMove;
        //    mon_tr.io_enq_req_1_bits_snapshot = io_enq_req_1_bits_snapshot;
        //    mon_tr.io_enq_req_1_bits_lqIdx_value = io_enq_req_1_bits_lqIdx_value;
        //    mon_tr.io_enq_req_1_bits_sqIdx_value = io_enq_req_1_bits_sqIdx_value;
        //    mon_tr.io_enq_req_1_bits_singleStep = io_enq_req_1_bits_singleStep;
        //    mon_tr.io_enq_req_1_bits_debug_sim_trig = io_enq_req_1_bits_debug_sim_trig;
        //    mon_tr.io_enq_req_2_valid = io_enq_req_2_valid;
        //    mon_tr.io_enq_req_2_bits_instr = io_enq_req_2_bits_instr;
        //    mon_tr.io_enq_req_2_bits_pc = io_enq_req_2_bits_pc;
        //    mon_tr.io_enq_req_2_bits_exceptionVec_0 = io_enq_req_2_bits_exceptionVec_0;
        //    mon_tr.io_enq_req_2_bits_exceptionVec_1 = io_enq_req_2_bits_exceptionVec_1;
        //    mon_tr.io_enq_req_2_bits_exceptionVec_2 = io_enq_req_2_bits_exceptionVec_2;
        //    mon_tr.io_enq_req_2_bits_exceptionVec_3 = io_enq_req_2_bits_exceptionVec_3;
        //    mon_tr.io_enq_req_2_bits_exceptionVec_12 = io_enq_req_2_bits_exceptionVec_12;
        //    mon_tr.io_enq_req_2_bits_exceptionVec_20 = io_enq_req_2_bits_exceptionVec_20;
        //    mon_tr.io_enq_req_2_bits_exceptionVec_22 = io_enq_req_2_bits_exceptionVec_22;
        //    mon_tr.io_enq_req_2_bits_isFetchMalAddr = io_enq_req_2_bits_isFetchMalAddr;
        //    mon_tr.io_enq_req_2_bits_hasException = io_enq_req_2_bits_hasException;
        //    mon_tr.io_enq_req_2_bits_trigger = io_enq_req_2_bits_trigger;
        //    mon_tr.io_enq_req_2_bits_preDecodeInfo_isRVC = io_enq_req_2_bits_preDecodeInfo_isRVC;
        //    mon_tr.io_enq_req_2_bits_crossPageIPFFix = io_enq_req_2_bits_crossPageIPFFix;
        //    mon_tr.io_enq_req_2_bits_ftqPtr_flag = io_enq_req_2_bits_ftqPtr_flag;
        //    mon_tr.io_enq_req_2_bits_ftqPtr_value = io_enq_req_2_bits_ftqPtr_value;
        //    mon_tr.io_enq_req_2_bits_ftqOffset = io_enq_req_2_bits_ftqOffset;
        //    mon_tr.io_enq_req_2_bits_ldest = io_enq_req_2_bits_ldest;
        //    mon_tr.io_enq_req_2_bits_fuType = io_enq_req_2_bits_fuType;
        //    mon_tr.io_enq_req_2_bits_fuOpType = io_enq_req_2_bits_fuOpType;
        //    mon_tr.io_enq_req_2_bits_rfWen = io_enq_req_2_bits_rfWen;
        //    mon_tr.io_enq_req_2_bits_fpWen = io_enq_req_2_bits_fpWen;
        //    mon_tr.io_enq_req_2_bits_vecWen = io_enq_req_2_bits_vecWen;
        //    mon_tr.io_enq_req_2_bits_v0Wen = io_enq_req_2_bits_v0Wen;
        //    mon_tr.io_enq_req_2_bits_vlWen = io_enq_req_2_bits_vlWen;
        //    mon_tr.io_enq_req_2_bits_isXSTrap = io_enq_req_2_bits_isXSTrap;
        //    mon_tr.io_enq_req_2_bits_waitForward = io_enq_req_2_bits_waitForward;
        //    mon_tr.io_enq_req_2_bits_blockBackward = io_enq_req_2_bits_blockBackward;
        //    mon_tr.io_enq_req_2_bits_flushPipe = io_enq_req_2_bits_flushPipe;
        //    mon_tr.io_enq_req_2_bits_vpu_vill = io_enq_req_2_bits_vpu_vill;
        //    mon_tr.io_enq_req_2_bits_vpu_vma = io_enq_req_2_bits_vpu_vma;
        //    mon_tr.io_enq_req_2_bits_vpu_vta = io_enq_req_2_bits_vpu_vta;
        //    mon_tr.io_enq_req_2_bits_vpu_vsew = io_enq_req_2_bits_vpu_vsew;
        //    mon_tr.io_enq_req_2_bits_vpu_vlmul = io_enq_req_2_bits_vpu_vlmul;
        //    mon_tr.io_enq_req_2_bits_vpu_specVill = io_enq_req_2_bits_vpu_specVill;
        //    mon_tr.io_enq_req_2_bits_vpu_specVma = io_enq_req_2_bits_vpu_specVma;
        //    mon_tr.io_enq_req_2_bits_vpu_specVta = io_enq_req_2_bits_vpu_specVta;
        //    mon_tr.io_enq_req_2_bits_vpu_specVsew = io_enq_req_2_bits_vpu_specVsew;
        //    mon_tr.io_enq_req_2_bits_vpu_specVlmul = io_enq_req_2_bits_vpu_specVlmul;
        //    mon_tr.io_enq_req_2_bits_vlsInstr = io_enq_req_2_bits_vlsInstr;
        //    mon_tr.io_enq_req_2_bits_wfflags = io_enq_req_2_bits_wfflags;
        //    mon_tr.io_enq_req_2_bits_isMove = io_enq_req_2_bits_isMove;
        //    mon_tr.io_enq_req_2_bits_isVset = io_enq_req_2_bits_isVset;
        //    mon_tr.io_enq_req_2_bits_firstUop = io_enq_req_2_bits_firstUop;
        //    mon_tr.io_enq_req_2_bits_lastUop = io_enq_req_2_bits_lastUop;
        //    mon_tr.io_enq_req_2_bits_numWB = io_enq_req_2_bits_numWB;
        //    mon_tr.io_enq_req_2_bits_commitType = io_enq_req_2_bits_commitType;
        //    mon_tr.io_enq_req_2_bits_pdest = io_enq_req_2_bits_pdest;
        //    mon_tr.io_enq_req_2_bits_robIdx_flag = io_enq_req_2_bits_robIdx_flag;
        //    mon_tr.io_enq_req_2_bits_robIdx_value = io_enq_req_2_bits_robIdx_value;
        //    mon_tr.io_enq_req_2_bits_instrSize = io_enq_req_2_bits_instrSize;
        //    mon_tr.io_enq_req_2_bits_dirtyFs = io_enq_req_2_bits_dirtyFs;
        //    mon_tr.io_enq_req_2_bits_dirtyVs = io_enq_req_2_bits_dirtyVs;
        //    mon_tr.io_enq_req_2_bits_traceBlockInPipe_itype = io_enq_req_2_bits_traceBlockInPipe_itype;
        //    mon_tr.io_enq_req_2_bits_traceBlockInPipe_iretire = io_enq_req_2_bits_traceBlockInPipe_iretire;
        //    mon_tr.io_enq_req_2_bits_traceBlockInPipe_ilastsize = io_enq_req_2_bits_traceBlockInPipe_ilastsize;
        //    mon_tr.io_enq_req_2_bits_eliminatedMove = io_enq_req_2_bits_eliminatedMove;
        //    mon_tr.io_enq_req_2_bits_snapshot = io_enq_req_2_bits_snapshot;
        //    mon_tr.io_enq_req_2_bits_lqIdx_value = io_enq_req_2_bits_lqIdx_value;
        //    mon_tr.io_enq_req_2_bits_sqIdx_value = io_enq_req_2_bits_sqIdx_value;
        //    mon_tr.io_enq_req_2_bits_singleStep = io_enq_req_2_bits_singleStep;
        //    mon_tr.io_enq_req_2_bits_debug_sim_trig = io_enq_req_2_bits_debug_sim_trig;
        //    mon_tr.io_enq_req_3_valid = io_enq_req_3_valid;
        //    mon_tr.io_enq_req_3_bits_instr = io_enq_req_3_bits_instr;
        //    mon_tr.io_enq_req_3_bits_pc = io_enq_req_3_bits_pc;
        //    mon_tr.io_enq_req_3_bits_exceptionVec_0 = io_enq_req_3_bits_exceptionVec_0;
        //    mon_tr.io_enq_req_3_bits_exceptionVec_1 = io_enq_req_3_bits_exceptionVec_1;
        //    mon_tr.io_enq_req_3_bits_exceptionVec_2 = io_enq_req_3_bits_exceptionVec_2;
        //    mon_tr.io_enq_req_3_bits_exceptionVec_3 = io_enq_req_3_bits_exceptionVec_3;
        //    mon_tr.io_enq_req_3_bits_exceptionVec_12 = io_enq_req_3_bits_exceptionVec_12;
        //    mon_tr.io_enq_req_3_bits_exceptionVec_20 = io_enq_req_3_bits_exceptionVec_20;
        //    mon_tr.io_enq_req_3_bits_exceptionVec_22 = io_enq_req_3_bits_exceptionVec_22;
        //    mon_tr.io_enq_req_3_bits_isFetchMalAddr = io_enq_req_3_bits_isFetchMalAddr;
        //    mon_tr.io_enq_req_3_bits_hasException = io_enq_req_3_bits_hasException;
        //    mon_tr.io_enq_req_3_bits_trigger = io_enq_req_3_bits_trigger;
        //    mon_tr.io_enq_req_3_bits_preDecodeInfo_isRVC = io_enq_req_3_bits_preDecodeInfo_isRVC;
        //    mon_tr.io_enq_req_3_bits_crossPageIPFFix = io_enq_req_3_bits_crossPageIPFFix;
        //    mon_tr.io_enq_req_3_bits_ftqPtr_flag = io_enq_req_3_bits_ftqPtr_flag;
        //    mon_tr.io_enq_req_3_bits_ftqPtr_value = io_enq_req_3_bits_ftqPtr_value;
        //    mon_tr.io_enq_req_3_bits_ftqOffset = io_enq_req_3_bits_ftqOffset;
        //    mon_tr.io_enq_req_3_bits_ldest = io_enq_req_3_bits_ldest;
        //    mon_tr.io_enq_req_3_bits_fuType = io_enq_req_3_bits_fuType;
        //    mon_tr.io_enq_req_3_bits_fuOpType = io_enq_req_3_bits_fuOpType;
        //    mon_tr.io_enq_req_3_bits_rfWen = io_enq_req_3_bits_rfWen;
        //    mon_tr.io_enq_req_3_bits_fpWen = io_enq_req_3_bits_fpWen;
        //    mon_tr.io_enq_req_3_bits_vecWen = io_enq_req_3_bits_vecWen;
        //    mon_tr.io_enq_req_3_bits_v0Wen = io_enq_req_3_bits_v0Wen;
        //    mon_tr.io_enq_req_3_bits_vlWen = io_enq_req_3_bits_vlWen;
        //    mon_tr.io_enq_req_3_bits_isXSTrap = io_enq_req_3_bits_isXSTrap;
        //    mon_tr.io_enq_req_3_bits_waitForward = io_enq_req_3_bits_waitForward;
        //    mon_tr.io_enq_req_3_bits_blockBackward = io_enq_req_3_bits_blockBackward;
        //    mon_tr.io_enq_req_3_bits_flushPipe = io_enq_req_3_bits_flushPipe;
        //    mon_tr.io_enq_req_3_bits_vpu_vill = io_enq_req_3_bits_vpu_vill;
        //    mon_tr.io_enq_req_3_bits_vpu_vma = io_enq_req_3_bits_vpu_vma;
        //    mon_tr.io_enq_req_3_bits_vpu_vta = io_enq_req_3_bits_vpu_vta;
        //    mon_tr.io_enq_req_3_bits_vpu_vsew = io_enq_req_3_bits_vpu_vsew;
        //    mon_tr.io_enq_req_3_bits_vpu_vlmul = io_enq_req_3_bits_vpu_vlmul;
        //    mon_tr.io_enq_req_3_bits_vpu_specVill = io_enq_req_3_bits_vpu_specVill;
        //    mon_tr.io_enq_req_3_bits_vpu_specVma = io_enq_req_3_bits_vpu_specVma;
        //    mon_tr.io_enq_req_3_bits_vpu_specVta = io_enq_req_3_bits_vpu_specVta;
        //    mon_tr.io_enq_req_3_bits_vpu_specVsew = io_enq_req_3_bits_vpu_specVsew;
        //    mon_tr.io_enq_req_3_bits_vpu_specVlmul = io_enq_req_3_bits_vpu_specVlmul;
        //    mon_tr.io_enq_req_3_bits_vlsInstr = io_enq_req_3_bits_vlsInstr;
        //    mon_tr.io_enq_req_3_bits_wfflags = io_enq_req_3_bits_wfflags;
        //    mon_tr.io_enq_req_3_bits_isMove = io_enq_req_3_bits_isMove;
        //    mon_tr.io_enq_req_3_bits_isVset = io_enq_req_3_bits_isVset;
        //    mon_tr.io_enq_req_3_bits_firstUop = io_enq_req_3_bits_firstUop;
        //    mon_tr.io_enq_req_3_bits_lastUop = io_enq_req_3_bits_lastUop;
        //    mon_tr.io_enq_req_3_bits_numWB = io_enq_req_3_bits_numWB;
        //    mon_tr.io_enq_req_3_bits_commitType = io_enq_req_3_bits_commitType;
        //    mon_tr.io_enq_req_3_bits_pdest = io_enq_req_3_bits_pdest;
        //    mon_tr.io_enq_req_3_bits_robIdx_flag = io_enq_req_3_bits_robIdx_flag;
        //    mon_tr.io_enq_req_3_bits_robIdx_value = io_enq_req_3_bits_robIdx_value;
        //    mon_tr.io_enq_req_3_bits_instrSize = io_enq_req_3_bits_instrSize;
        //    mon_tr.io_enq_req_3_bits_dirtyFs = io_enq_req_3_bits_dirtyFs;
        //    mon_tr.io_enq_req_3_bits_dirtyVs = io_enq_req_3_bits_dirtyVs;
        //    mon_tr.io_enq_req_3_bits_traceBlockInPipe_itype = io_enq_req_3_bits_traceBlockInPipe_itype;
        //    mon_tr.io_enq_req_3_bits_traceBlockInPipe_iretire = io_enq_req_3_bits_traceBlockInPipe_iretire;
        //    mon_tr.io_enq_req_3_bits_traceBlockInPipe_ilastsize = io_enq_req_3_bits_traceBlockInPipe_ilastsize;
        //    mon_tr.io_enq_req_3_bits_eliminatedMove = io_enq_req_3_bits_eliminatedMove;
        //    mon_tr.io_enq_req_3_bits_snapshot = io_enq_req_3_bits_snapshot;
        //    mon_tr.io_enq_req_3_bits_lqIdx_value = io_enq_req_3_bits_lqIdx_value;
        //    mon_tr.io_enq_req_3_bits_sqIdx_value = io_enq_req_3_bits_sqIdx_value;
        //    mon_tr.io_enq_req_3_bits_singleStep = io_enq_req_3_bits_singleStep;
        //    mon_tr.io_enq_req_3_bits_debug_sim_trig = io_enq_req_3_bits_debug_sim_trig;
        //    mon_tr.io_enq_req_4_valid = io_enq_req_4_valid;
        //    mon_tr.io_enq_req_4_bits_instr = io_enq_req_4_bits_instr;
        //    mon_tr.io_enq_req_4_bits_pc = io_enq_req_4_bits_pc;
        //    mon_tr.io_enq_req_4_bits_exceptionVec_0 = io_enq_req_4_bits_exceptionVec_0;
        //    mon_tr.io_enq_req_4_bits_exceptionVec_1 = io_enq_req_4_bits_exceptionVec_1;
        //    mon_tr.io_enq_req_4_bits_exceptionVec_2 = io_enq_req_4_bits_exceptionVec_2;
        //    mon_tr.io_enq_req_4_bits_exceptionVec_3 = io_enq_req_4_bits_exceptionVec_3;
        //    mon_tr.io_enq_req_4_bits_exceptionVec_12 = io_enq_req_4_bits_exceptionVec_12;
        //    mon_tr.io_enq_req_4_bits_exceptionVec_20 = io_enq_req_4_bits_exceptionVec_20;
        //    mon_tr.io_enq_req_4_bits_exceptionVec_22 = io_enq_req_4_bits_exceptionVec_22;
        //    mon_tr.io_enq_req_4_bits_isFetchMalAddr = io_enq_req_4_bits_isFetchMalAddr;
        //    mon_tr.io_enq_req_4_bits_hasException = io_enq_req_4_bits_hasException;
        //    mon_tr.io_enq_req_4_bits_trigger = io_enq_req_4_bits_trigger;
        //    mon_tr.io_enq_req_4_bits_preDecodeInfo_isRVC = io_enq_req_4_bits_preDecodeInfo_isRVC;
        //    mon_tr.io_enq_req_4_bits_crossPageIPFFix = io_enq_req_4_bits_crossPageIPFFix;
        //    mon_tr.io_enq_req_4_bits_ftqPtr_flag = io_enq_req_4_bits_ftqPtr_flag;
        //    mon_tr.io_enq_req_4_bits_ftqPtr_value = io_enq_req_4_bits_ftqPtr_value;
        //    mon_tr.io_enq_req_4_bits_ftqOffset = io_enq_req_4_bits_ftqOffset;
        //    mon_tr.io_enq_req_4_bits_ldest = io_enq_req_4_bits_ldest;
        //    mon_tr.io_enq_req_4_bits_fuType = io_enq_req_4_bits_fuType;
        //    mon_tr.io_enq_req_4_bits_fuOpType = io_enq_req_4_bits_fuOpType;
        //    mon_tr.io_enq_req_4_bits_rfWen = io_enq_req_4_bits_rfWen;
        //    mon_tr.io_enq_req_4_bits_fpWen = io_enq_req_4_bits_fpWen;
        //    mon_tr.io_enq_req_4_bits_vecWen = io_enq_req_4_bits_vecWen;
        //    mon_tr.io_enq_req_4_bits_v0Wen = io_enq_req_4_bits_v0Wen;
        //    mon_tr.io_enq_req_4_bits_vlWen = io_enq_req_4_bits_vlWen;
        //    mon_tr.io_enq_req_4_bits_isXSTrap = io_enq_req_4_bits_isXSTrap;
        //    mon_tr.io_enq_req_4_bits_waitForward = io_enq_req_4_bits_waitForward;
        //    mon_tr.io_enq_req_4_bits_blockBackward = io_enq_req_4_bits_blockBackward;
        //    mon_tr.io_enq_req_4_bits_flushPipe = io_enq_req_4_bits_flushPipe;
        //    mon_tr.io_enq_req_4_bits_vpu_vill = io_enq_req_4_bits_vpu_vill;
        //    mon_tr.io_enq_req_4_bits_vpu_vma = io_enq_req_4_bits_vpu_vma;
        //    mon_tr.io_enq_req_4_bits_vpu_vta = io_enq_req_4_bits_vpu_vta;
        //    mon_tr.io_enq_req_4_bits_vpu_vsew = io_enq_req_4_bits_vpu_vsew;
        //    mon_tr.io_enq_req_4_bits_vpu_vlmul = io_enq_req_4_bits_vpu_vlmul;
        //    mon_tr.io_enq_req_4_bits_vpu_specVill = io_enq_req_4_bits_vpu_specVill;
        //    mon_tr.io_enq_req_4_bits_vpu_specVma = io_enq_req_4_bits_vpu_specVma;
        //    mon_tr.io_enq_req_4_bits_vpu_specVta = io_enq_req_4_bits_vpu_specVta;
        //    mon_tr.io_enq_req_4_bits_vpu_specVsew = io_enq_req_4_bits_vpu_specVsew;
        //    mon_tr.io_enq_req_4_bits_vpu_specVlmul = io_enq_req_4_bits_vpu_specVlmul;
        //    mon_tr.io_enq_req_4_bits_vlsInstr = io_enq_req_4_bits_vlsInstr;
        //    mon_tr.io_enq_req_4_bits_wfflags = io_enq_req_4_bits_wfflags;
        //    mon_tr.io_enq_req_4_bits_isMove = io_enq_req_4_bits_isMove;
        //    mon_tr.io_enq_req_4_bits_isVset = io_enq_req_4_bits_isVset;
        //    mon_tr.io_enq_req_4_bits_firstUop = io_enq_req_4_bits_firstUop;
        //    mon_tr.io_enq_req_4_bits_lastUop = io_enq_req_4_bits_lastUop;
        //    mon_tr.io_enq_req_4_bits_numWB = io_enq_req_4_bits_numWB;
        //    mon_tr.io_enq_req_4_bits_commitType = io_enq_req_4_bits_commitType;
        //    mon_tr.io_enq_req_4_bits_pdest = io_enq_req_4_bits_pdest;
        //    mon_tr.io_enq_req_4_bits_robIdx_flag = io_enq_req_4_bits_robIdx_flag;
        //    mon_tr.io_enq_req_4_bits_robIdx_value = io_enq_req_4_bits_robIdx_value;
        //    mon_tr.io_enq_req_4_bits_instrSize = io_enq_req_4_bits_instrSize;
        //    mon_tr.io_enq_req_4_bits_dirtyFs = io_enq_req_4_bits_dirtyFs;
        //    mon_tr.io_enq_req_4_bits_dirtyVs = io_enq_req_4_bits_dirtyVs;
        //    mon_tr.io_enq_req_4_bits_traceBlockInPipe_itype = io_enq_req_4_bits_traceBlockInPipe_itype;
        //    mon_tr.io_enq_req_4_bits_traceBlockInPipe_iretire = io_enq_req_4_bits_traceBlockInPipe_iretire;
        //    mon_tr.io_enq_req_4_bits_traceBlockInPipe_ilastsize = io_enq_req_4_bits_traceBlockInPipe_ilastsize;
        //    mon_tr.io_enq_req_4_bits_eliminatedMove = io_enq_req_4_bits_eliminatedMove;
        //    mon_tr.io_enq_req_4_bits_snapshot = io_enq_req_4_bits_snapshot;
        //    mon_tr.io_enq_req_4_bits_lqIdx_value = io_enq_req_4_bits_lqIdx_value;
        //    mon_tr.io_enq_req_4_bits_sqIdx_value = io_enq_req_4_bits_sqIdx_value;
        //    mon_tr.io_enq_req_4_bits_singleStep = io_enq_req_4_bits_singleStep;
        //    mon_tr.io_enq_req_4_bits_debug_sim_trig = io_enq_req_4_bits_debug_sim_trig;
        //    mon_tr.io_enq_req_5_valid = io_enq_req_5_valid;
        //    mon_tr.io_enq_req_5_bits_instr = io_enq_req_5_bits_instr;
        //    mon_tr.io_enq_req_5_bits_pc = io_enq_req_5_bits_pc;
        //    mon_tr.io_enq_req_5_bits_exceptionVec_0 = io_enq_req_5_bits_exceptionVec_0;
        //    mon_tr.io_enq_req_5_bits_exceptionVec_1 = io_enq_req_5_bits_exceptionVec_1;
        //    mon_tr.io_enq_req_5_bits_exceptionVec_2 = io_enq_req_5_bits_exceptionVec_2;
        //    mon_tr.io_enq_req_5_bits_exceptionVec_3 = io_enq_req_5_bits_exceptionVec_3;
        //    mon_tr.io_enq_req_5_bits_exceptionVec_12 = io_enq_req_5_bits_exceptionVec_12;
        //    mon_tr.io_enq_req_5_bits_exceptionVec_20 = io_enq_req_5_bits_exceptionVec_20;
        //    mon_tr.io_enq_req_5_bits_exceptionVec_22 = io_enq_req_5_bits_exceptionVec_22;
        //    mon_tr.io_enq_req_5_bits_isFetchMalAddr = io_enq_req_5_bits_isFetchMalAddr;
        //    mon_tr.io_enq_req_5_bits_hasException = io_enq_req_5_bits_hasException;
        //    mon_tr.io_enq_req_5_bits_trigger = io_enq_req_5_bits_trigger;
        //    mon_tr.io_enq_req_5_bits_preDecodeInfo_isRVC = io_enq_req_5_bits_preDecodeInfo_isRVC;
        //    mon_tr.io_enq_req_5_bits_crossPageIPFFix = io_enq_req_5_bits_crossPageIPFFix;
        //    mon_tr.io_enq_req_5_bits_ftqPtr_flag = io_enq_req_5_bits_ftqPtr_flag;
        //    mon_tr.io_enq_req_5_bits_ftqPtr_value = io_enq_req_5_bits_ftqPtr_value;
        //    mon_tr.io_enq_req_5_bits_ftqOffset = io_enq_req_5_bits_ftqOffset;
        //    mon_tr.io_enq_req_5_bits_ldest = io_enq_req_5_bits_ldest;
        //    mon_tr.io_enq_req_5_bits_fuType = io_enq_req_5_bits_fuType;
        //    mon_tr.io_enq_req_5_bits_fuOpType = io_enq_req_5_bits_fuOpType;
        //    mon_tr.io_enq_req_5_bits_rfWen = io_enq_req_5_bits_rfWen;
        //    mon_tr.io_enq_req_5_bits_fpWen = io_enq_req_5_bits_fpWen;
        //    mon_tr.io_enq_req_5_bits_vecWen = io_enq_req_5_bits_vecWen;
        //    mon_tr.io_enq_req_5_bits_v0Wen = io_enq_req_5_bits_v0Wen;
        //    mon_tr.io_enq_req_5_bits_vlWen = io_enq_req_5_bits_vlWen;
        //    mon_tr.io_enq_req_5_bits_isXSTrap = io_enq_req_5_bits_isXSTrap;
        //    mon_tr.io_enq_req_5_bits_waitForward = io_enq_req_5_bits_waitForward;
        //    mon_tr.io_enq_req_5_bits_blockBackward = io_enq_req_5_bits_blockBackward;
        //    mon_tr.io_enq_req_5_bits_flushPipe = io_enq_req_5_bits_flushPipe;
        //    mon_tr.io_enq_req_5_bits_vpu_vill = io_enq_req_5_bits_vpu_vill;
        //    mon_tr.io_enq_req_5_bits_vpu_vma = io_enq_req_5_bits_vpu_vma;
        //    mon_tr.io_enq_req_5_bits_vpu_vta = io_enq_req_5_bits_vpu_vta;
        //    mon_tr.io_enq_req_5_bits_vpu_vsew = io_enq_req_5_bits_vpu_vsew;
        //    mon_tr.io_enq_req_5_bits_vpu_vlmul = io_enq_req_5_bits_vpu_vlmul;
        //    mon_tr.io_enq_req_5_bits_vpu_specVill = io_enq_req_5_bits_vpu_specVill;
        //    mon_tr.io_enq_req_5_bits_vpu_specVma = io_enq_req_5_bits_vpu_specVma;
        //    mon_tr.io_enq_req_5_bits_vpu_specVta = io_enq_req_5_bits_vpu_specVta;
        //    mon_tr.io_enq_req_5_bits_vpu_specVsew = io_enq_req_5_bits_vpu_specVsew;
        //    mon_tr.io_enq_req_5_bits_vpu_specVlmul = io_enq_req_5_bits_vpu_specVlmul;
        //    mon_tr.io_enq_req_5_bits_vlsInstr = io_enq_req_5_bits_vlsInstr;
        //    mon_tr.io_enq_req_5_bits_wfflags = io_enq_req_5_bits_wfflags;
        //    mon_tr.io_enq_req_5_bits_isMove = io_enq_req_5_bits_isMove;
        //    mon_tr.io_enq_req_5_bits_isVset = io_enq_req_5_bits_isVset;
        //    mon_tr.io_enq_req_5_bits_firstUop = io_enq_req_5_bits_firstUop;
        //    mon_tr.io_enq_req_5_bits_lastUop = io_enq_req_5_bits_lastUop;
        //    mon_tr.io_enq_req_5_bits_numWB = io_enq_req_5_bits_numWB;
        //    mon_tr.io_enq_req_5_bits_commitType = io_enq_req_5_bits_commitType;
        //    mon_tr.io_enq_req_5_bits_pdest = io_enq_req_5_bits_pdest;
        //    mon_tr.io_enq_req_5_bits_robIdx_flag = io_enq_req_5_bits_robIdx_flag;
        //    mon_tr.io_enq_req_5_bits_robIdx_value = io_enq_req_5_bits_robIdx_value;
        //    mon_tr.io_enq_req_5_bits_instrSize = io_enq_req_5_bits_instrSize;
        //    mon_tr.io_enq_req_5_bits_dirtyFs = io_enq_req_5_bits_dirtyFs;
        //    mon_tr.io_enq_req_5_bits_dirtyVs = io_enq_req_5_bits_dirtyVs;
        //    mon_tr.io_enq_req_5_bits_traceBlockInPipe_itype = io_enq_req_5_bits_traceBlockInPipe_itype;
        //    mon_tr.io_enq_req_5_bits_traceBlockInPipe_iretire = io_enq_req_5_bits_traceBlockInPipe_iretire;
        //    mon_tr.io_enq_req_5_bits_traceBlockInPipe_ilastsize = io_enq_req_5_bits_traceBlockInPipe_ilastsize;
        //    mon_tr.io_enq_req_5_bits_eliminatedMove = io_enq_req_5_bits_eliminatedMove;
        //    mon_tr.io_enq_req_5_bits_snapshot = io_enq_req_5_bits_snapshot;
        //    mon_tr.io_enq_req_5_bits_lqIdx_value = io_enq_req_5_bits_lqIdx_value;
        //    mon_tr.io_enq_req_5_bits_sqIdx_value = io_enq_req_5_bits_sqIdx_value;
        //    mon_tr.io_enq_req_5_bits_singleStep = io_enq_req_5_bits_singleStep;
        //    mon_tr.io_enq_req_5_bits_debug_sim_trig = io_enq_req_5_bits_debug_sim_trig;

        //    mon_tr.channel_id = this.cfg.channel_id;
        //    mon_tr.unpack();
        //    this.mon_item_port.write(mon_tr);
        //end
    end
endtask:mon_data

`endif


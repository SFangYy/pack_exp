//=========================================================
//File name    : CSR_in_agent_dec.sv
//Author       : nanyunhao
//Module name  : CSR_in_agent_dec
//Discribution : CSR_in_agent_dec : parameter
//Date         : 2026-01-22
//=========================================================
`ifndef CSR_IN_AGENT_DEC__SV
`define CSR_IN_AGENT_DEC__SV

package CSR_in_agent_dec;

endpackage:CSR_in_agent_dec

import CSR_in_agent_dec::*;

`endif


//=========================================================
//File name    : Rob_dec.sv
//Author       : nanyunhao
//Module name  : Rob_dec
//Discribution : Rob_dec : common parameter
//Date         : 2026-01-22
//=========================================================
`ifndef ROB_DEC__SV
`define ROB_DEC__SV

package Rob_dec;

endpackage

import Rob_dec::*;

`endif


//=========================================================
//File name    : dut_inst.sv
//Author       : nanyunhao
//Module name  : dut_inst
//Discribution : dut_inst : DUT instance
//Date         : 2026-01-22
//=========================================================
`ifndef DUT_INST__SV
`define DUT_INST__SV

//rename_in
reg         clock                  ;
reg         reset                  ;
reg [5:0]   io_hartId              ;
reg         io_enq_req_0_valid     ;
reg [31:0]  io_enq_req_0_bits_instr;
reg [49:0]  io_enq_req_0_bits_pc   ;
reg         io_enq_req_0_bits_exceptionVec_0;
reg         io_enq_req_0_bits_exceptionVec_1;
reg         io_enq_req_0_bits_exceptionVec_2;
reg         io_enq_req_0_bits_exceptionVec_3;
reg         io_enq_req_0_bits_exceptionVec_12;
reg         io_enq_req_0_bits_exceptionVec_20;
reg         io_enq_req_0_bits_exceptionVec_22;
reg         io_enq_req_0_bits_isFetchMalAddr;
reg         io_enq_req_0_bits_hasException;
reg [3:0]   io_enq_req_0_bits_trigger;
reg         io_enq_req_0_bits_preDecodeInfo_isRVC;
reg         io_enq_req_0_bits_crossPageIPFFix;
reg         io_enq_req_0_bits_ftqPtr_flag;
reg [5:0]   io_enq_req_0_bits_ftqPtr_value;
reg [3:0]   io_enq_req_0_bits_ftqOffset;
reg [5:0]   io_enq_req_0_bits_ldest;
reg [34:0]  io_enq_req_0_bits_fuType;
reg [8:0]   io_enq_req_0_bits_fuOpType;
reg         io_enq_req_0_bits_rfWen;
reg         io_enq_req_0_bits_fpWen;
reg         io_enq_req_0_bits_vecWen;
reg         io_enq_req_0_bits_v0Wen;
reg         io_enq_req_0_bits_vlWen;
reg         io_enq_req_0_bits_isXSTrap;
reg         io_enq_req_0_bits_waitForward;
reg         io_enq_req_0_bits_blockBackward;
reg         io_enq_req_0_bits_flushPipe;
reg         io_enq_req_0_bits_vpu_vill;
reg         io_enq_req_0_bits_vpu_vma;
reg         io_enq_req_0_bits_vpu_vta;
reg [1:0]   io_enq_req_0_bits_vpu_vsew;
reg [2:0]   io_enq_req_0_bits_vpu_vlmul;
reg         io_enq_req_0_bits_vpu_specVill;
reg         io_enq_req_0_bits_vpu_specVma;
reg         io_enq_req_0_bits_vpu_specVta;
reg [1:0]   io_enq_req_0_bits_vpu_specVsew;
reg [2:0]   io_enq_req_0_bits_vpu_specVlmul;
reg         io_enq_req_0_bits_vlsInstr;
reg         io_enq_req_0_bits_wfflags;
reg         io_enq_req_0_bits_isMove;
reg         io_enq_req_0_bits_isVset;
reg         io_enq_req_0_bits_firstUop;
reg         io_enq_req_0_bits_lastUop;
reg [6:0]   io_enq_req_0_bits_numWB;
reg [2:0]   io_enq_req_0_bits_commitType;
reg [7:0]   io_enq_req_0_bits_pdest;
reg         io_enq_req_0_bits_robIdx_flag;
reg [7:0]   io_enq_req_0_bits_robIdx_value;
reg [2:0]   io_enq_req_0_bits_instrSize;
reg         io_enq_req_0_bits_dirtyFs;
reg         io_enq_req_0_bits_dirtyVs;
reg [3:0]   io_enq_req_0_bits_traceBlockInPipe_itype;
reg [3:0]   io_enq_req_0_bits_traceBlockInPipe_iretire;
reg         io_enq_req_0_bits_traceBlockInPipe_ilastsize;
reg         io_enq_req_0_bits_eliminatedMove;
reg         io_enq_req_0_bits_snapshot;
reg [6:0]   io_enq_req_0_bits_lqIdx_value;
reg [5:0]   io_enq_req_0_bits_sqIdx_value;
reg         io_enq_req_0_bits_singleStep;
reg         io_enq_req_0_bits_debug_sim_trig;
reg         io_enq_req_1_valid     ;
reg [31:0]  io_enq_req_1_bits_instr;
reg [49:0]  io_enq_req_1_bits_pc   ;
reg         io_enq_req_1_bits_exceptionVec_0;
reg         io_enq_req_1_bits_exceptionVec_1;
reg         io_enq_req_1_bits_exceptionVec_2;
reg         io_enq_req_1_bits_exceptionVec_3;
reg         io_enq_req_1_bits_exceptionVec_12;
reg         io_enq_req_1_bits_exceptionVec_20;
reg         io_enq_req_1_bits_exceptionVec_22;
reg         io_enq_req_1_bits_isFetchMalAddr;
reg         io_enq_req_1_bits_hasException;
reg [3:0]   io_enq_req_1_bits_trigger;
reg         io_enq_req_1_bits_preDecodeInfo_isRVC;
reg         io_enq_req_1_bits_crossPageIPFFix;
reg         io_enq_req_1_bits_ftqPtr_flag;
reg [5:0]   io_enq_req_1_bits_ftqPtr_value;
reg [3:0]   io_enq_req_1_bits_ftqOffset;
reg [5:0]   io_enq_req_1_bits_ldest;
reg [34:0]  io_enq_req_1_bits_fuType;
reg [8:0]   io_enq_req_1_bits_fuOpType;
reg         io_enq_req_1_bits_rfWen;
reg         io_enq_req_1_bits_fpWen;
reg         io_enq_req_1_bits_vecWen;
reg         io_enq_req_1_bits_v0Wen;
reg         io_enq_req_1_bits_vlWen;
reg         io_enq_req_1_bits_isXSTrap;
reg         io_enq_req_1_bits_waitForward;
reg         io_enq_req_1_bits_blockBackward;
reg         io_enq_req_1_bits_flushPipe;
reg         io_enq_req_1_bits_vpu_vill;
reg         io_enq_req_1_bits_vpu_vma;
reg         io_enq_req_1_bits_vpu_vta;
reg [1:0]   io_enq_req_1_bits_vpu_vsew;
reg [2:0]   io_enq_req_1_bits_vpu_vlmul;
reg         io_enq_req_1_bits_vpu_specVill;
reg         io_enq_req_1_bits_vpu_specVma;
reg         io_enq_req_1_bits_vpu_specVta;
reg [1:0]   io_enq_req_1_bits_vpu_specVsew;
reg [2:0]   io_enq_req_1_bits_vpu_specVlmul;
reg         io_enq_req_1_bits_vlsInstr;
reg         io_enq_req_1_bits_wfflags;
reg         io_enq_req_1_bits_isMove;
reg         io_enq_req_1_bits_isVset;
reg         io_enq_req_1_bits_firstUop;
reg         io_enq_req_1_bits_lastUop;
reg [6:0]   io_enq_req_1_bits_numWB;
reg [2:0]   io_enq_req_1_bits_commitType;
reg [7:0]   io_enq_req_1_bits_pdest;
reg         io_enq_req_1_bits_robIdx_flag;
reg [7:0]   io_enq_req_1_bits_robIdx_value;
reg [2:0]   io_enq_req_1_bits_instrSize;
reg         io_enq_req_1_bits_dirtyFs;
reg         io_enq_req_1_bits_dirtyVs;
reg [3:0]   io_enq_req_1_bits_traceBlockInPipe_itype;
reg [3:0]   io_enq_req_1_bits_traceBlockInPipe_iretire;
reg         io_enq_req_1_bits_traceBlockInPipe_ilastsize;
reg         io_enq_req_1_bits_eliminatedMove;
reg         io_enq_req_1_bits_snapshot;
reg [6:0]   io_enq_req_1_bits_lqIdx_value;
reg [5:0]   io_enq_req_1_bits_sqIdx_value;
reg         io_enq_req_1_bits_singleStep;
reg         io_enq_req_1_bits_debug_sim_trig;
reg         io_enq_req_2_valid     ;
reg [31:0]  io_enq_req_2_bits_instr;
reg [49:0]  io_enq_req_2_bits_pc   ;
reg         io_enq_req_2_bits_exceptionVec_0;
reg         io_enq_req_2_bits_exceptionVec_1;
reg         io_enq_req_2_bits_exceptionVec_2;
reg         io_enq_req_2_bits_exceptionVec_3;
reg         io_enq_req_2_bits_exceptionVec_12;
reg         io_enq_req_2_bits_exceptionVec_20;
reg         io_enq_req_2_bits_exceptionVec_22;
reg         io_enq_req_2_bits_isFetchMalAddr;
reg         io_enq_req_2_bits_hasException;
reg [3:0]   io_enq_req_2_bits_trigger;
reg         io_enq_req_2_bits_preDecodeInfo_isRVC;
reg         io_enq_req_2_bits_crossPageIPFFix;
reg         io_enq_req_2_bits_ftqPtr_flag;
reg [5:0]   io_enq_req_2_bits_ftqPtr_value;
reg [3:0]   io_enq_req_2_bits_ftqOffset;
reg [5:0]   io_enq_req_2_bits_ldest;
reg [34:0]  io_enq_req_2_bits_fuType;
reg [8:0]   io_enq_req_2_bits_fuOpType;
reg         io_enq_req_2_bits_rfWen;
reg         io_enq_req_2_bits_fpWen;
reg         io_enq_req_2_bits_vecWen;
reg         io_enq_req_2_bits_v0Wen;
reg         io_enq_req_2_bits_vlWen;
reg         io_enq_req_2_bits_isXSTrap;
reg         io_enq_req_2_bits_waitForward;
reg         io_enq_req_2_bits_blockBackward;
reg         io_enq_req_2_bits_flushPipe;
reg         io_enq_req_2_bits_vpu_vill;
reg         io_enq_req_2_bits_vpu_vma;
reg         io_enq_req_2_bits_vpu_vta;
reg [1:0]   io_enq_req_2_bits_vpu_vsew;
reg [2:0]   io_enq_req_2_bits_vpu_vlmul;
reg         io_enq_req_2_bits_vpu_specVill;
reg         io_enq_req_2_bits_vpu_specVma;
reg         io_enq_req_2_bits_vpu_specVta;
reg [1:0]   io_enq_req_2_bits_vpu_specVsew;
reg [2:0]   io_enq_req_2_bits_vpu_specVlmul;
reg         io_enq_req_2_bits_vlsInstr;
reg         io_enq_req_2_bits_wfflags;
reg         io_enq_req_2_bits_isMove;
reg         io_enq_req_2_bits_isVset;
reg         io_enq_req_2_bits_firstUop;
reg         io_enq_req_2_bits_lastUop;
reg [6:0]   io_enq_req_2_bits_numWB;
reg [2:0]   io_enq_req_2_bits_commitType;
reg [7:0]   io_enq_req_2_bits_pdest;
reg         io_enq_req_2_bits_robIdx_flag;
reg [7:0]   io_enq_req_2_bits_robIdx_value;
reg [2:0]   io_enq_req_2_bits_instrSize;
reg         io_enq_req_2_bits_dirtyFs;
reg         io_enq_req_2_bits_dirtyVs;
reg [3:0]   io_enq_req_2_bits_traceBlockInPipe_itype;
reg [3:0]   io_enq_req_2_bits_traceBlockInPipe_iretire;
reg         io_enq_req_2_bits_traceBlockInPipe_ilastsize;
reg         io_enq_req_2_bits_eliminatedMove;
reg         io_enq_req_2_bits_snapshot;
reg [6:0]   io_enq_req_2_bits_lqIdx_value;
reg [5:0]   io_enq_req_2_bits_sqIdx_value;
reg         io_enq_req_2_bits_singleStep;
reg         io_enq_req_2_bits_debug_sim_trig;
reg         io_enq_req_3_valid     ;
reg [31:0]  io_enq_req_3_bits_instr;
reg [49:0]  io_enq_req_3_bits_pc   ;
reg         io_enq_req_3_bits_exceptionVec_0;
reg         io_enq_req_3_bits_exceptionVec_1;
reg         io_enq_req_3_bits_exceptionVec_2;
reg         io_enq_req_3_bits_exceptionVec_3;
reg         io_enq_req_3_bits_exceptionVec_12;
reg         io_enq_req_3_bits_exceptionVec_20;
reg         io_enq_req_3_bits_exceptionVec_22;
reg         io_enq_req_3_bits_isFetchMalAddr;
reg         io_enq_req_3_bits_hasException;
reg [3:0]   io_enq_req_3_bits_trigger;
reg         io_enq_req_3_bits_preDecodeInfo_isRVC;
reg         io_enq_req_3_bits_crossPageIPFFix;
reg         io_enq_req_3_bits_ftqPtr_flag;
reg [5:0]   io_enq_req_3_bits_ftqPtr_value;
reg [3:0]   io_enq_req_3_bits_ftqOffset;
reg [5:0]   io_enq_req_3_bits_ldest;
reg [34:0]  io_enq_req_3_bits_fuType;
reg [8:0]   io_enq_req_3_bits_fuOpType;
reg         io_enq_req_3_bits_rfWen;
reg         io_enq_req_3_bits_fpWen;
reg         io_enq_req_3_bits_vecWen;
reg         io_enq_req_3_bits_v0Wen;
reg         io_enq_req_3_bits_vlWen;
reg         io_enq_req_3_bits_isXSTrap;
reg         io_enq_req_3_bits_waitForward;
reg         io_enq_req_3_bits_blockBackward;
reg         io_enq_req_3_bits_flushPipe;
reg         io_enq_req_3_bits_vpu_vill;
reg         io_enq_req_3_bits_vpu_vma;
reg         io_enq_req_3_bits_vpu_vta;
reg [1:0]   io_enq_req_3_bits_vpu_vsew;
reg [2:0]   io_enq_req_3_bits_vpu_vlmul;
reg         io_enq_req_3_bits_vpu_specVill;
reg         io_enq_req_3_bits_vpu_specVma;
reg         io_enq_req_3_bits_vpu_specVta;
reg [1:0]   io_enq_req_3_bits_vpu_specVsew;
reg [2:0]   io_enq_req_3_bits_vpu_specVlmul;
reg         io_enq_req_3_bits_vlsInstr;
reg         io_enq_req_3_bits_wfflags;
reg         io_enq_req_3_bits_isMove;
reg         io_enq_req_3_bits_isVset;
reg         io_enq_req_3_bits_firstUop;
reg         io_enq_req_3_bits_lastUop;
reg [6:0]   io_enq_req_3_bits_numWB;
reg [2:0]   io_enq_req_3_bits_commitType;
reg [7:0]   io_enq_req_3_bits_pdest;
reg         io_enq_req_3_bits_robIdx_flag;
reg [7:0]   io_enq_req_3_bits_robIdx_value;
reg [2:0]   io_enq_req_3_bits_instrSize;
reg         io_enq_req_3_bits_dirtyFs;
reg         io_enq_req_3_bits_dirtyVs;
reg [3:0]   io_enq_req_3_bits_traceBlockInPipe_itype;
reg [3:0]   io_enq_req_3_bits_traceBlockInPipe_iretire;
reg         io_enq_req_3_bits_traceBlockInPipe_ilastsize;
reg         io_enq_req_3_bits_eliminatedMove;
reg         io_enq_req_3_bits_snapshot;
reg [6:0]   io_enq_req_3_bits_lqIdx_value;
reg [5:0]   io_enq_req_3_bits_sqIdx_value;
reg         io_enq_req_3_bits_singleStep;
reg         io_enq_req_3_bits_debug_sim_trig;
reg         io_enq_req_4_valid     ;
reg [31:0]  io_enq_req_4_bits_instr;
reg [49:0]  io_enq_req_4_bits_pc   ;
reg         io_enq_req_4_bits_exceptionVec_0;
reg         io_enq_req_4_bits_exceptionVec_1;
reg         io_enq_req_4_bits_exceptionVec_2;
reg         io_enq_req_4_bits_exceptionVec_3;
reg         io_enq_req_4_bits_exceptionVec_12;
reg         io_enq_req_4_bits_exceptionVec_20;
reg         io_enq_req_4_bits_exceptionVec_22;
reg         io_enq_req_4_bits_isFetchMalAddr;
reg         io_enq_req_4_bits_hasException;
reg [3:0]   io_enq_req_4_bits_trigger;
reg         io_enq_req_4_bits_preDecodeInfo_isRVC;
reg         io_enq_req_4_bits_crossPageIPFFix;
reg         io_enq_req_4_bits_ftqPtr_flag;
reg [5:0]   io_enq_req_4_bits_ftqPtr_value;
reg [3:0]   io_enq_req_4_bits_ftqOffset;
reg [5:0]   io_enq_req_4_bits_ldest;
reg [34:0]  io_enq_req_4_bits_fuType;
reg [8:0]   io_enq_req_4_bits_fuOpType;
reg         io_enq_req_4_bits_rfWen;
reg         io_enq_req_4_bits_fpWen;
reg         io_enq_req_4_bits_vecWen;
reg         io_enq_req_4_bits_v0Wen;
reg         io_enq_req_4_bits_vlWen;
reg         io_enq_req_4_bits_isXSTrap;
reg         io_enq_req_4_bits_waitForward;
reg         io_enq_req_4_bits_blockBackward;
reg         io_enq_req_4_bits_flushPipe;
reg         io_enq_req_4_bits_vpu_vill;
reg         io_enq_req_4_bits_vpu_vma;
reg         io_enq_req_4_bits_vpu_vta;
reg [1:0]   io_enq_req_4_bits_vpu_vsew;
reg [2:0]   io_enq_req_4_bits_vpu_vlmul;
reg         io_enq_req_4_bits_vpu_specVill;
reg         io_enq_req_4_bits_vpu_specVma;
reg         io_enq_req_4_bits_vpu_specVta;
reg [1:0]   io_enq_req_4_bits_vpu_specVsew;
reg [2:0]   io_enq_req_4_bits_vpu_specVlmul;
reg         io_enq_req_4_bits_vlsInstr;
reg         io_enq_req_4_bits_wfflags;
reg         io_enq_req_4_bits_isMove;
reg         io_enq_req_4_bits_isVset;
reg         io_enq_req_4_bits_firstUop;
reg         io_enq_req_4_bits_lastUop;
reg [6:0]   io_enq_req_4_bits_numWB;
reg [2:0]   io_enq_req_4_bits_commitType;
reg [7:0]   io_enq_req_4_bits_pdest;
reg         io_enq_req_4_bits_robIdx_flag;
reg [7:0]   io_enq_req_4_bits_robIdx_value;
reg [2:0]   io_enq_req_4_bits_instrSize;
reg         io_enq_req_4_bits_dirtyFs;
reg         io_enq_req_4_bits_dirtyVs;
reg [3:0]   io_enq_req_4_bits_traceBlockInPipe_itype;
reg [3:0]   io_enq_req_4_bits_traceBlockInPipe_iretire;
reg         io_enq_req_4_bits_traceBlockInPipe_ilastsize;
reg         io_enq_req_4_bits_eliminatedMove;
reg         io_enq_req_4_bits_snapshot;
reg [6:0]   io_enq_req_4_bits_lqIdx_value;
reg [5:0]   io_enq_req_4_bits_sqIdx_value;
reg         io_enq_req_4_bits_singleStep;
reg         io_enq_req_4_bits_debug_sim_trig;
reg         io_enq_req_5_valid     ;
reg [31:0]  io_enq_req_5_bits_instr;
reg [49:0]  io_enq_req_5_bits_pc   ;
reg         io_enq_req_5_bits_exceptionVec_0;
reg         io_enq_req_5_bits_exceptionVec_1;
reg         io_enq_req_5_bits_exceptionVec_2;
reg         io_enq_req_5_bits_exceptionVec_3;
reg         io_enq_req_5_bits_exceptionVec_12;
reg         io_enq_req_5_bits_exceptionVec_20;
reg         io_enq_req_5_bits_exceptionVec_22;
reg         io_enq_req_5_bits_isFetchMalAddr;
reg         io_enq_req_5_bits_hasException;
reg [3:0]   io_enq_req_5_bits_trigger;
reg         io_enq_req_5_bits_preDecodeInfo_isRVC;
reg         io_enq_req_5_bits_crossPageIPFFix;
reg         io_enq_req_5_bits_ftqPtr_flag;
reg [5:0]   io_enq_req_5_bits_ftqPtr_value;
reg [3:0]   io_enq_req_5_bits_ftqOffset;
reg [5:0]   io_enq_req_5_bits_ldest;
reg [34:0]  io_enq_req_5_bits_fuType;
reg [8:0]   io_enq_req_5_bits_fuOpType;
reg         io_enq_req_5_bits_rfWen;
reg         io_enq_req_5_bits_fpWen;
reg         io_enq_req_5_bits_vecWen;
reg         io_enq_req_5_bits_v0Wen;
reg         io_enq_req_5_bits_vlWen;
reg         io_enq_req_5_bits_isXSTrap;
reg         io_enq_req_5_bits_waitForward;
reg         io_enq_req_5_bits_blockBackward;
reg         io_enq_req_5_bits_flushPipe;
reg         io_enq_req_5_bits_vpu_vill;
reg         io_enq_req_5_bits_vpu_vma;
reg         io_enq_req_5_bits_vpu_vta;
reg [1:0]   io_enq_req_5_bits_vpu_vsew;
reg [2:0]   io_enq_req_5_bits_vpu_vlmul;
reg         io_enq_req_5_bits_vpu_specVill;
reg         io_enq_req_5_bits_vpu_specVma;
reg         io_enq_req_5_bits_vpu_specVta;
reg [1:0]   io_enq_req_5_bits_vpu_specVsew;
reg [2:0]   io_enq_req_5_bits_vpu_specVlmul;
reg         io_enq_req_5_bits_vlsInstr;
reg         io_enq_req_5_bits_wfflags;
reg         io_enq_req_5_bits_isMove;
reg         io_enq_req_5_bits_isVset;
reg         io_enq_req_5_bits_firstUop;
reg         io_enq_req_5_bits_lastUop;
reg [6:0]   io_enq_req_5_bits_numWB;
reg [2:0]   io_enq_req_5_bits_commitType;
reg [7:0]   io_enq_req_5_bits_pdest;
reg         io_enq_req_5_bits_robIdx_flag;
reg [7:0]   io_enq_req_5_bits_robIdx_value;
reg [2:0]   io_enq_req_5_bits_instrSize;
reg         io_enq_req_5_bits_dirtyFs;
reg         io_enq_req_5_bits_dirtyVs;
reg [3:0]   io_enq_req_5_bits_traceBlockInPipe_itype;
reg [3:0]   io_enq_req_5_bits_traceBlockInPipe_iretire;
reg         io_enq_req_5_bits_traceBlockInPipe_ilastsize;
reg         io_enq_req_5_bits_eliminatedMove;
reg         io_enq_req_5_bits_snapshot;
reg [6:0]   io_enq_req_5_bits_lqIdx_value;
reg [5:0]   io_enq_req_5_bits_sqIdx_value;
reg         io_enq_req_5_bits_singleStep;
reg         io_enq_req_5_bits_debug_sim_trig;
//WriteBack_in
reg         io_writeback_24_valid  ;
reg [127:0] io_writeback_24_bits_data_0;
reg [6:0]   io_writeback_24_bits_pdest;
reg         io_writeback_24_bits_robIdx_flag;
reg [7:0]   io_writeback_24_bits_robIdx_value;
reg         io_writeback_24_bits_vecWen;
reg         io_writeback_24_bits_v0Wen;
reg         io_writeback_24_bits_vlWen;
reg         io_writeback_24_bits_exceptionVec_0;
reg         io_writeback_24_bits_exceptionVec_1;
reg         io_writeback_24_bits_exceptionVec_2;
reg         io_writeback_24_bits_exceptionVec_3;
reg         io_writeback_24_bits_exceptionVec_4;
reg         io_writeback_24_bits_exceptionVec_5;
reg         io_writeback_24_bits_exceptionVec_6;
reg         io_writeback_24_bits_exceptionVec_7;
reg         io_writeback_24_bits_exceptionVec_8;
reg         io_writeback_24_bits_exceptionVec_9;
reg         io_writeback_24_bits_exceptionVec_10;
reg         io_writeback_24_bits_exceptionVec_11;
reg         io_writeback_24_bits_exceptionVec_12;
reg         io_writeback_24_bits_exceptionVec_13;
reg         io_writeback_24_bits_exceptionVec_14;
reg         io_writeback_24_bits_exceptionVec_15;
reg         io_writeback_24_bits_exceptionVec_16;
reg         io_writeback_24_bits_exceptionVec_17;
reg         io_writeback_24_bits_exceptionVec_18;
reg         io_writeback_24_bits_exceptionVec_19;
reg         io_writeback_24_bits_exceptionVec_20;
reg         io_writeback_24_bits_exceptionVec_21;
reg         io_writeback_24_bits_exceptionVec_22;
reg         io_writeback_24_bits_exceptionVec_23;
reg         io_writeback_24_bits_flushPipe;
reg         io_writeback_24_bits_replay;
reg [3:0]   io_writeback_24_bits_trigger;
reg         io_writeback_24_bits_vls_vpu_vill;
reg         io_writeback_24_bits_vls_vpu_vma;
reg         io_writeback_24_bits_vls_vpu_vta;
reg [1:0]   io_writeback_24_bits_vls_vpu_vsew;
reg [2:0]   io_writeback_24_bits_vls_vpu_vlmul;
reg         io_writeback_24_bits_vls_vpu_specVill;
reg         io_writeback_24_bits_vls_vpu_specVma;
reg         io_writeback_24_bits_vls_vpu_specVta;
reg [1:0]   io_writeback_24_bits_vls_vpu_specVsew;
reg [2:0]   io_writeback_24_bits_vls_vpu_specVlmul;
reg         io_writeback_24_bits_vls_vpu_vm;
reg [7:0]   io_writeback_24_bits_vls_vpu_vstart;
reg [2:0]   io_writeback_24_bits_vls_vpu_frm;
reg         io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst;
reg         io_writeback_24_bits_vls_vpu_fpu_isFP32Instr;
reg         io_writeback_24_bits_vls_vpu_fpu_isFP64Instr;
reg         io_writeback_24_bits_vls_vpu_fpu_isReduction;
reg         io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2;
reg         io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4;
reg         io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8;
reg [1:0]   io_writeback_24_bits_vls_vpu_vxrm;
reg [6:0]   io_writeback_24_bits_vls_vpu_vuopIdx;
reg         io_writeback_24_bits_vls_vpu_lastUop;
reg [127:0] io_writeback_24_bits_vls_vpu_vmask;
reg [7:0]   io_writeback_24_bits_vls_vpu_vl;
reg [2:0]   io_writeback_24_bits_vls_vpu_nf;
reg [1:0]   io_writeback_24_bits_vls_vpu_veew;
reg         io_writeback_24_bits_vls_vpu_isReverse;
reg         io_writeback_24_bits_vls_vpu_isExt;
reg         io_writeback_24_bits_vls_vpu_isNarrow;
reg         io_writeback_24_bits_vls_vpu_isDstMask;
reg         io_writeback_24_bits_vls_vpu_isOpMask;
reg         io_writeback_24_bits_vls_vpu_isMove;
reg         io_writeback_24_bits_vls_vpu_isDependOldVd;
reg         io_writeback_24_bits_vls_vpu_isWritePartVd;
reg         io_writeback_24_bits_vls_vpu_isVleff;
reg [7:0]   io_writeback_24_bits_vls_oldVdPsrc;
reg [2:0]   io_writeback_24_bits_vls_vdIdx;
reg [2:0]   io_writeback_24_bits_vls_vdIdxInField;
reg         io_writeback_24_bits_vls_isIndexed;
reg         io_writeback_24_bits_vls_isMasked;
reg         io_writeback_24_bits_vls_isStrided;
reg         io_writeback_24_bits_vls_isWhole;
reg         io_writeback_24_bits_vls_isVecLoad;
reg         io_writeback_24_bits_vls_isVlm;
reg         io_writeback_24_bits_debug_isMMIO;
reg         io_writeback_24_bits_debug_isNCIO;
reg         io_writeback_24_bits_debug_isPerfCnt;
reg [47:0]  io_writeback_24_bits_debug_paddr;
reg [49:0]  io_writeback_24_bits_debug_vaddr;
reg         io_writeback_24_bits_debugInfo_eliminatedMove;
reg [63:0]  io_writeback_24_bits_debugInfo_renameTime;
reg [63:0]  io_writeback_24_bits_debugInfo_dispatchTime;
reg [63:0]  io_writeback_24_bits_debugInfo_enqRsTime;
reg [63:0]  io_writeback_24_bits_debugInfo_selectTime;
reg [63:0]  io_writeback_24_bits_debugInfo_issueTime;
reg [63:0]  io_writeback_24_bits_debugInfo_writebackTime;
reg [63:0]  io_writeback_24_bits_debugInfo_runahead_checkpoint_id;
reg [63:0]  io_writeback_24_bits_debugInfo_tlbFirstReqTime;
reg [63:0]  io_writeback_24_bits_debugInfo_tlbRespTime;
reg [63:0]  io_writeback_24_bits_debug_seqNum;
reg         io_writeback_23_valid  ;
reg [127:0] io_writeback_23_bits_data_0;
reg [6:0]   io_writeback_23_bits_pdest;
reg         io_writeback_23_bits_robIdx_flag;
reg [7:0]   io_writeback_23_bits_robIdx_value;
reg         io_writeback_23_bits_vecWen;
reg         io_writeback_23_bits_v0Wen;
reg         io_writeback_23_bits_vlWen;
reg         io_writeback_23_bits_exceptionVec_0;
reg         io_writeback_23_bits_exceptionVec_1;
reg         io_writeback_23_bits_exceptionVec_2;
reg         io_writeback_23_bits_exceptionVec_3;
reg         io_writeback_23_bits_exceptionVec_4;
reg         io_writeback_23_bits_exceptionVec_5;
reg         io_writeback_23_bits_exceptionVec_6;
reg         io_writeback_23_bits_exceptionVec_7;
reg         io_writeback_23_bits_exceptionVec_8;
reg         io_writeback_23_bits_exceptionVec_9;
reg         io_writeback_23_bits_exceptionVec_10;
reg         io_writeback_23_bits_exceptionVec_11;
reg         io_writeback_23_bits_exceptionVec_12;
reg         io_writeback_23_bits_exceptionVec_13;
reg         io_writeback_23_bits_exceptionVec_14;
reg         io_writeback_23_bits_exceptionVec_15;
reg         io_writeback_23_bits_exceptionVec_16;
reg         io_writeback_23_bits_exceptionVec_17;
reg         io_writeback_23_bits_exceptionVec_18;
reg         io_writeback_23_bits_exceptionVec_19;
reg         io_writeback_23_bits_exceptionVec_20;
reg         io_writeback_23_bits_exceptionVec_21;
reg         io_writeback_23_bits_exceptionVec_22;
reg         io_writeback_23_bits_exceptionVec_23;
reg         io_writeback_23_bits_flushPipe;
reg         io_writeback_23_bits_replay;
reg [3:0]   io_writeback_23_bits_trigger;
reg         io_writeback_23_bits_vls_vpu_vill;
reg         io_writeback_23_bits_vls_vpu_vma;
reg         io_writeback_23_bits_vls_vpu_vta;
reg [1:0]   io_writeback_23_bits_vls_vpu_vsew;
reg [2:0]   io_writeback_23_bits_vls_vpu_vlmul;
reg         io_writeback_23_bits_vls_vpu_specVill;
reg         io_writeback_23_bits_vls_vpu_specVma;
reg         io_writeback_23_bits_vls_vpu_specVta;
reg [1:0]   io_writeback_23_bits_vls_vpu_specVsew;
reg [2:0]   io_writeback_23_bits_vls_vpu_specVlmul;
reg         io_writeback_23_bits_vls_vpu_vm;
reg [7:0]   io_writeback_23_bits_vls_vpu_vstart;
reg [2:0]   io_writeback_23_bits_vls_vpu_frm;
reg         io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst;
reg         io_writeback_23_bits_vls_vpu_fpu_isFP32Instr;
reg         io_writeback_23_bits_vls_vpu_fpu_isFP64Instr;
reg         io_writeback_23_bits_vls_vpu_fpu_isReduction;
reg         io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2;
reg         io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4;
reg         io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8;
reg [1:0]   io_writeback_23_bits_vls_vpu_vxrm;
reg [6:0]   io_writeback_23_bits_vls_vpu_vuopIdx;
reg         io_writeback_23_bits_vls_vpu_lastUop;
reg [127:0] io_writeback_23_bits_vls_vpu_vmask;
reg [7:0]   io_writeback_23_bits_vls_vpu_vl;
reg [2:0]   io_writeback_23_bits_vls_vpu_nf;
reg [1:0]   io_writeback_23_bits_vls_vpu_veew;
reg         io_writeback_23_bits_vls_vpu_isReverse;
reg         io_writeback_23_bits_vls_vpu_isExt;
reg         io_writeback_23_bits_vls_vpu_isNarrow;
reg         io_writeback_23_bits_vls_vpu_isDstMask;
reg         io_writeback_23_bits_vls_vpu_isOpMask;
reg         io_writeback_23_bits_vls_vpu_isMove;
reg         io_writeback_23_bits_vls_vpu_isDependOldVd;
reg         io_writeback_23_bits_vls_vpu_isWritePartVd;
reg         io_writeback_23_bits_vls_vpu_isVleff;
reg [7:0]   io_writeback_23_bits_vls_oldVdPsrc;
reg [2:0]   io_writeback_23_bits_vls_vdIdx;
reg [2:0]   io_writeback_23_bits_vls_vdIdxInField;
reg         io_writeback_23_bits_vls_isIndexed;
reg         io_writeback_23_bits_vls_isMasked;
reg         io_writeback_23_bits_vls_isStrided;
reg         io_writeback_23_bits_vls_isWhole;
reg         io_writeback_23_bits_vls_isVecLoad;
reg         io_writeback_23_bits_vls_isVlm;
reg         io_writeback_23_bits_debug_isMMIO;
reg         io_writeback_23_bits_debug_isNCIO;
reg         io_writeback_23_bits_debug_isPerfCnt;
reg [47:0]  io_writeback_23_bits_debug_paddr;
reg [49:0]  io_writeback_23_bits_debug_vaddr;
reg         io_writeback_23_bits_debugInfo_eliminatedMove;
reg [63:0]  io_writeback_23_bits_debugInfo_renameTime;
reg [63:0]  io_writeback_23_bits_debugInfo_dispatchTime;
reg [63:0]  io_writeback_23_bits_debugInfo_enqRsTime;
reg [63:0]  io_writeback_23_bits_debugInfo_selectTime;
reg [63:0]  io_writeback_23_bits_debugInfo_issueTime;
reg [63:0]  io_writeback_23_bits_debugInfo_writebackTime;
reg [63:0]  io_writeback_23_bits_debugInfo_runahead_checkpoint_id;
reg [63:0]  io_writeback_23_bits_debugInfo_tlbFirstReqTime;
reg [63:0]  io_writeback_23_bits_debugInfo_tlbRespTime;
reg [63:0]  io_writeback_23_bits_debug_seqNum;
reg         io_writeback_22_valid  ;
reg [63:0]  io_writeback_22_bits_data_0;
reg [7:0]   io_writeback_22_bits_pdest;
reg         io_writeback_22_bits_robIdx_flag;
reg [7:0]   io_writeback_22_bits_robIdx_value;
reg         io_writeback_22_bits_intWen;
reg         io_writeback_22_bits_fpWen;
reg         io_writeback_22_bits_exceptionVec_0;
reg         io_writeback_22_bits_exceptionVec_1;
reg         io_writeback_22_bits_exceptionVec_2;
reg         io_writeback_22_bits_exceptionVec_3;
reg         io_writeback_22_bits_exceptionVec_4;
reg         io_writeback_22_bits_exceptionVec_5;
reg         io_writeback_22_bits_exceptionVec_6;
reg         io_writeback_22_bits_exceptionVec_7;
reg         io_writeback_22_bits_exceptionVec_8;
reg         io_writeback_22_bits_exceptionVec_9;
reg         io_writeback_22_bits_exceptionVec_10;
reg         io_writeback_22_bits_exceptionVec_11;
reg         io_writeback_22_bits_exceptionVec_12;
reg         io_writeback_22_bits_exceptionVec_13;
reg         io_writeback_22_bits_exceptionVec_14;
reg         io_writeback_22_bits_exceptionVec_15;
reg         io_writeback_22_bits_exceptionVec_16;
reg         io_writeback_22_bits_exceptionVec_17;
reg         io_writeback_22_bits_exceptionVec_18;
reg         io_writeback_22_bits_exceptionVec_19;
reg         io_writeback_22_bits_exceptionVec_20;
reg         io_writeback_22_bits_exceptionVec_21;
reg         io_writeback_22_bits_exceptionVec_22;
reg         io_writeback_22_bits_exceptionVec_23;
reg         io_writeback_22_bits_flushPipe;
reg         io_writeback_22_bits_replay;
reg         io_writeback_22_bits_lqIdx_flag;
reg [6:0]   io_writeback_22_bits_lqIdx_value;
reg [3:0]   io_writeback_22_bits_trigger;
reg         io_writeback_22_bits_predecodeInfo_valid;
reg         io_writeback_22_bits_predecodeInfo_isRVC;
reg [1:0]   io_writeback_22_bits_predecodeInfo_brType;
reg         io_writeback_22_bits_predecodeInfo_isCall;
reg         io_writeback_22_bits_predecodeInfo_isRet;
reg         io_writeback_22_bits_debug_isMMIO;
reg         io_writeback_22_bits_debug_isNCIO;
reg         io_writeback_22_bits_debug_isPerfCnt;
reg [47:0]  io_writeback_22_bits_debug_paddr;
reg [49:0]  io_writeback_22_bits_debug_vaddr;
reg         io_writeback_22_bits_debugInfo_eliminatedMove;
reg [63:0]  io_writeback_22_bits_debugInfo_renameTime;
reg [63:0]  io_writeback_22_bits_debugInfo_dispatchTime;
reg [63:0]  io_writeback_22_bits_debugInfo_enqRsTime;
reg [63:0]  io_writeback_22_bits_debugInfo_selectTime;
reg [63:0]  io_writeback_22_bits_debugInfo_issueTime;
reg [63:0]  io_writeback_22_bits_debugInfo_writebackTime;
reg [63:0]  io_writeback_22_bits_debugInfo_runahead_checkpoint_id;
reg [63:0]  io_writeback_22_bits_debugInfo_tlbFirstReqTime;
reg [63:0]  io_writeback_22_bits_debugInfo_tlbRespTime;
reg [63:0]  io_writeback_22_bits_debug_seqNum;
reg         io_writeback_21_valid  ;
reg [63:0]  io_writeback_21_bits_data_0;
reg [7:0]   io_writeback_21_bits_pdest;
reg         io_writeback_21_bits_robIdx_flag;
reg [7:0]   io_writeback_21_bits_robIdx_value;
reg         io_writeback_21_bits_intWen;
reg         io_writeback_21_bits_fpWen;
reg         io_writeback_21_bits_exceptionVec_0;
reg         io_writeback_21_bits_exceptionVec_1;
reg         io_writeback_21_bits_exceptionVec_2;
reg         io_writeback_21_bits_exceptionVec_3;
reg         io_writeback_21_bits_exceptionVec_4;
reg         io_writeback_21_bits_exceptionVec_5;
reg         io_writeback_21_bits_exceptionVec_6;
reg         io_writeback_21_bits_exceptionVec_7;
reg         io_writeback_21_bits_exceptionVec_8;
reg         io_writeback_21_bits_exceptionVec_9;
reg         io_writeback_21_bits_exceptionVec_10;
reg         io_writeback_21_bits_exceptionVec_11;
reg         io_writeback_21_bits_exceptionVec_12;
reg         io_writeback_21_bits_exceptionVec_13;
reg         io_writeback_21_bits_exceptionVec_14;
reg         io_writeback_21_bits_exceptionVec_15;
reg         io_writeback_21_bits_exceptionVec_16;
reg         io_writeback_21_bits_exceptionVec_17;
reg         io_writeback_21_bits_exceptionVec_18;
reg         io_writeback_21_bits_exceptionVec_19;
reg         io_writeback_21_bits_exceptionVec_20;
reg         io_writeback_21_bits_exceptionVec_21;
reg         io_writeback_21_bits_exceptionVec_22;
reg         io_writeback_21_bits_exceptionVec_23;
reg         io_writeback_21_bits_flushPipe;
reg         io_writeback_21_bits_replay;
reg         io_writeback_21_bits_lqIdx_flag;
reg [6:0]   io_writeback_21_bits_lqIdx_value;
reg [3:0]   io_writeback_21_bits_trigger;
reg         io_writeback_21_bits_predecodeInfo_valid;
reg         io_writeback_21_bits_predecodeInfo_isRVC;
reg [1:0]   io_writeback_21_bits_predecodeInfo_brType;
reg         io_writeback_21_bits_predecodeInfo_isCall;
reg         io_writeback_21_bits_predecodeInfo_isRet;
reg         io_writeback_21_bits_debug_isMMIO;
reg         io_writeback_21_bits_debug_isNCIO;
reg         io_writeback_21_bits_debug_isPerfCnt;
reg [47:0]  io_writeback_21_bits_debug_paddr;
reg [49:0]  io_writeback_21_bits_debug_vaddr;
reg         io_writeback_21_bits_debugInfo_eliminatedMove;
reg [63:0]  io_writeback_21_bits_debugInfo_renameTime;
reg [63:0]  io_writeback_21_bits_debugInfo_dispatchTime;
reg [63:0]  io_writeback_21_bits_debugInfo_enqRsTime;
reg [63:0]  io_writeback_21_bits_debugInfo_selectTime;
reg [63:0]  io_writeback_21_bits_debugInfo_issueTime;
reg [63:0]  io_writeback_21_bits_debugInfo_writebackTime;
reg [63:0]  io_writeback_21_bits_debugInfo_runahead_checkpoint_id;
reg [63:0]  io_writeback_21_bits_debugInfo_tlbFirstReqTime;
reg [63:0]  io_writeback_21_bits_debugInfo_tlbRespTime;
reg [63:0]  io_writeback_21_bits_debug_seqNum;
reg         io_writeback_20_valid  ;
reg [63:0]  io_writeback_20_bits_data_0;
reg [7:0]   io_writeback_20_bits_pdest;
reg         io_writeback_20_bits_robIdx_flag;
reg [7:0]   io_writeback_20_bits_robIdx_value;
reg         io_writeback_20_bits_intWen;
reg         io_writeback_20_bits_fpWen;
reg         io_writeback_20_bits_exceptionVec_0;
reg         io_writeback_20_bits_exceptionVec_1;
reg         io_writeback_20_bits_exceptionVec_2;
reg         io_writeback_20_bits_exceptionVec_3;
reg         io_writeback_20_bits_exceptionVec_4;
reg         io_writeback_20_bits_exceptionVec_5;
reg         io_writeback_20_bits_exceptionVec_6;
reg         io_writeback_20_bits_exceptionVec_7;
reg         io_writeback_20_bits_exceptionVec_8;
reg         io_writeback_20_bits_exceptionVec_9;
reg         io_writeback_20_bits_exceptionVec_10;
reg         io_writeback_20_bits_exceptionVec_11;
reg         io_writeback_20_bits_exceptionVec_12;
reg         io_writeback_20_bits_exceptionVec_13;
reg         io_writeback_20_bits_exceptionVec_14;
reg         io_writeback_20_bits_exceptionVec_15;
reg         io_writeback_20_bits_exceptionVec_16;
reg         io_writeback_20_bits_exceptionVec_17;
reg         io_writeback_20_bits_exceptionVec_18;
reg         io_writeback_20_bits_exceptionVec_19;
reg         io_writeback_20_bits_exceptionVec_20;
reg         io_writeback_20_bits_exceptionVec_21;
reg         io_writeback_20_bits_exceptionVec_22;
reg         io_writeback_20_bits_exceptionVec_23;
reg         io_writeback_20_bits_flushPipe;
reg         io_writeback_20_bits_replay;
reg         io_writeback_20_bits_lqIdx_flag;
reg [6:0]   io_writeback_20_bits_lqIdx_value;
reg [3:0]   io_writeback_20_bits_trigger;
reg         io_writeback_20_bits_predecodeInfo_valid;
reg         io_writeback_20_bits_predecodeInfo_isRVC;
reg [1:0]   io_writeback_20_bits_predecodeInfo_brType;
reg         io_writeback_20_bits_predecodeInfo_isCall;
reg         io_writeback_20_bits_predecodeInfo_isRet;
reg         io_writeback_20_bits_debug_isMMIO;
reg         io_writeback_20_bits_debug_isNCIO;
reg         io_writeback_20_bits_debug_isPerfCnt;
reg [47:0]  io_writeback_20_bits_debug_paddr;
reg [49:0]  io_writeback_20_bits_debug_vaddr;
reg         io_writeback_20_bits_debugInfo_eliminatedMove;
reg [63:0]  io_writeback_20_bits_debugInfo_renameTime;
reg [63:0]  io_writeback_20_bits_debugInfo_dispatchTime;
reg [63:0]  io_writeback_20_bits_debugInfo_enqRsTime;
reg [63:0]  io_writeback_20_bits_debugInfo_selectTime;
reg [63:0]  io_writeback_20_bits_debugInfo_issueTime;
reg [63:0]  io_writeback_20_bits_debugInfo_writebackTime;
reg [63:0]  io_writeback_20_bits_debugInfo_runahead_checkpoint_id;
reg [63:0]  io_writeback_20_bits_debugInfo_tlbFirstReqTime;
reg [63:0]  io_writeback_20_bits_debugInfo_tlbRespTime;
reg [63:0]  io_writeback_20_bits_debug_seqNum;
reg         io_writeback_19_valid  ;
reg [63:0]  io_writeback_19_bits_data_0;
reg [7:0]   io_writeback_19_bits_pdest;
reg         io_writeback_19_bits_robIdx_flag;
reg [7:0]   io_writeback_19_bits_robIdx_value;
reg         io_writeback_19_bits_intWen;
reg         io_writeback_19_bits_exceptionVec_0;
reg         io_writeback_19_bits_exceptionVec_1;
reg         io_writeback_19_bits_exceptionVec_2;
reg         io_writeback_19_bits_exceptionVec_3;
reg         io_writeback_19_bits_exceptionVec_4;
reg         io_writeback_19_bits_exceptionVec_5;
reg         io_writeback_19_bits_exceptionVec_6;
reg         io_writeback_19_bits_exceptionVec_7;
reg         io_writeback_19_bits_exceptionVec_8;
reg         io_writeback_19_bits_exceptionVec_9;
reg         io_writeback_19_bits_exceptionVec_10;
reg         io_writeback_19_bits_exceptionVec_11;
reg         io_writeback_19_bits_exceptionVec_12;
reg         io_writeback_19_bits_exceptionVec_13;
reg         io_writeback_19_bits_exceptionVec_14;
reg         io_writeback_19_bits_exceptionVec_15;
reg         io_writeback_19_bits_exceptionVec_16;
reg         io_writeback_19_bits_exceptionVec_17;
reg         io_writeback_19_bits_exceptionVec_18;
reg         io_writeback_19_bits_exceptionVec_19;
reg         io_writeback_19_bits_exceptionVec_20;
reg         io_writeback_19_bits_exceptionVec_21;
reg         io_writeback_19_bits_exceptionVec_22;
reg         io_writeback_19_bits_exceptionVec_23;
reg         io_writeback_19_bits_flushPipe;
reg         io_writeback_19_bits_sqIdx_flag;
reg [5:0]   io_writeback_19_bits_sqIdx_value;
reg [3:0]   io_writeback_19_bits_trigger;
reg         io_writeback_19_bits_debug_isMMIO;
reg         io_writeback_19_bits_debug_isNCIO;
reg         io_writeback_19_bits_debug_isPerfCnt;
reg [47:0]  io_writeback_19_bits_debug_paddr;
reg [49:0]  io_writeback_19_bits_debug_vaddr;
reg         io_writeback_19_bits_debugInfo_eliminatedMove;
reg [63:0]  io_writeback_19_bits_debugInfo_renameTime;
reg [63:0]  io_writeback_19_bits_debugInfo_dispatchTime;
reg [63:0]  io_writeback_19_bits_debugInfo_enqRsTime;
reg [63:0]  io_writeback_19_bits_debugInfo_selectTime;
reg [63:0]  io_writeback_19_bits_debugInfo_issueTime;
reg [63:0]  io_writeback_19_bits_debugInfo_writebackTime;
reg [63:0]  io_writeback_19_bits_debugInfo_runahead_checkpoint_id;
reg [63:0]  io_writeback_19_bits_debugInfo_tlbFirstReqTime;
reg [63:0]  io_writeback_19_bits_debugInfo_tlbRespTime;
reg [63:0]  io_writeback_19_bits_debug_seqNum;
reg         io_writeback_18_valid  ;
reg [63:0]  io_writeback_18_bits_data_0;
reg [7:0]   io_writeback_18_bits_pdest;
reg         io_writeback_18_bits_robIdx_flag;
reg [7:0]   io_writeback_18_bits_robIdx_value;
reg         io_writeback_18_bits_intWen;
reg         io_writeback_18_bits_exceptionVec_0;
reg         io_writeback_18_bits_exceptionVec_1;
reg         io_writeback_18_bits_exceptionVec_2;
reg         io_writeback_18_bits_exceptionVec_3;
reg         io_writeback_18_bits_exceptionVec_4;
reg         io_writeback_18_bits_exceptionVec_5;
reg         io_writeback_18_bits_exceptionVec_6;
reg         io_writeback_18_bits_exceptionVec_7;
reg         io_writeback_18_bits_exceptionVec_8;
reg         io_writeback_18_bits_exceptionVec_9;
reg         io_writeback_18_bits_exceptionVec_10;
reg         io_writeback_18_bits_exceptionVec_11;
reg         io_writeback_18_bits_exceptionVec_12;
reg         io_writeback_18_bits_exceptionVec_13;
reg         io_writeback_18_bits_exceptionVec_14;
reg         io_writeback_18_bits_exceptionVec_15;
reg         io_writeback_18_bits_exceptionVec_16;
reg         io_writeback_18_bits_exceptionVec_17;
reg         io_writeback_18_bits_exceptionVec_18;
reg         io_writeback_18_bits_exceptionVec_19;
reg         io_writeback_18_bits_exceptionVec_20;
reg         io_writeback_18_bits_exceptionVec_21;
reg         io_writeback_18_bits_exceptionVec_22;
reg         io_writeback_18_bits_exceptionVec_23;
reg         io_writeback_18_bits_flushPipe;
reg         io_writeback_18_bits_sqIdx_flag;
reg [5:0]   io_writeback_18_bits_sqIdx_value;
reg [3:0]   io_writeback_18_bits_trigger;
reg         io_writeback_18_bits_debug_isMMIO;
reg         io_writeback_18_bits_debug_isNCIO;
reg         io_writeback_18_bits_debug_isPerfCnt;
reg [47:0]  io_writeback_18_bits_debug_paddr;
reg [49:0]  io_writeback_18_bits_debug_vaddr;
reg         io_writeback_18_bits_debugInfo_eliminatedMove;
reg [63:0]  io_writeback_18_bits_debugInfo_renameTime;
reg [63:0]  io_writeback_18_bits_debugInfo_dispatchTime;
reg [63:0]  io_writeback_18_bits_debugInfo_enqRsTime;
reg [63:0]  io_writeback_18_bits_debugInfo_selectTime;
reg [63:0]  io_writeback_18_bits_debugInfo_issueTime;
reg [63:0]  io_writeback_18_bits_debugInfo_writebackTime;
reg [63:0]  io_writeback_18_bits_debugInfo_runahead_checkpoint_id;
reg [63:0]  io_writeback_18_bits_debugInfo_tlbFirstReqTime;
reg [63:0]  io_writeback_18_bits_debugInfo_tlbRespTime;
reg [63:0]  io_writeback_18_bits_debug_seqNum;
reg         io_writeback_17_valid  ;
reg [127:0] io_writeback_17_bits_data_0;
reg [127:0] io_writeback_17_bits_data_1;
reg [127:0] io_writeback_17_bits_data_2;
reg [6:0]   io_writeback_17_bits_pdest;
reg         io_writeback_17_bits_robIdx_flag;
reg [7:0]   io_writeback_17_bits_robIdx_value;
reg         io_writeback_17_bits_vecWen;
reg         io_writeback_17_bits_v0Wen;
reg [4:0]   io_writeback_17_bits_fflags;
reg         io_writeback_17_bits_wflags;
reg         io_writeback_17_bits_debugInfo_eliminatedMove;
reg [63:0]  io_writeback_17_bits_debugInfo_renameTime;
reg [63:0]  io_writeback_17_bits_debugInfo_dispatchTime;
reg [63:0]  io_writeback_17_bits_debugInfo_enqRsTime;
reg [63:0]  io_writeback_17_bits_debugInfo_selectTime;
reg [63:0]  io_writeback_17_bits_debugInfo_issueTime;
reg [63:0]  io_writeback_17_bits_debugInfo_writebackTime;
reg [63:0]  io_writeback_17_bits_debugInfo_runahead_checkpoint_id;
reg [63:0]  io_writeback_17_bits_debugInfo_tlbFirstReqTime;
reg [63:0]  io_writeback_17_bits_debugInfo_tlbRespTime;
reg [63:0]  io_writeback_17_bits_debug_seqNum;
reg         io_writeback_16_valid  ;
reg [127:0] io_writeback_16_bits_data_0;
reg [127:0] io_writeback_16_bits_data_1;
reg [127:0] io_writeback_16_bits_data_2;
reg [127:0] io_writeback_16_bits_data_3;
reg [7:0]   io_writeback_16_bits_pdest;
reg         io_writeback_16_bits_robIdx_flag;
reg [7:0]   io_writeback_16_bits_robIdx_value;
reg         io_writeback_16_bits_fpWen;
reg         io_writeback_16_bits_vecWen;
reg         io_writeback_16_bits_v0Wen;
reg [4:0]   io_writeback_16_bits_fflags;
reg         io_writeback_16_bits_wflags;
reg         io_writeback_16_bits_debugInfo_eliminatedMove;
reg [63:0]  io_writeback_16_bits_debugInfo_renameTime;
reg [63:0]  io_writeback_16_bits_debugInfo_dispatchTime;
reg [63:0]  io_writeback_16_bits_debugInfo_enqRsTime;
reg [63:0]  io_writeback_16_bits_debugInfo_selectTime;
reg [63:0]  io_writeback_16_bits_debugInfo_issueTime;
reg [63:0]  io_writeback_16_bits_debugInfo_writebackTime;
reg [63:0]  io_writeback_16_bits_debugInfo_runahead_checkpoint_id;
reg [63:0]  io_writeback_16_bits_debugInfo_tlbFirstReqTime;
reg [63:0]  io_writeback_16_bits_debugInfo_tlbRespTime;
reg [63:0]  io_writeback_16_bits_debug_seqNum;
reg         io_writeback_15_valid  ;
reg [127:0] io_writeback_15_bits_data_0;
reg [127:0] io_writeback_15_bits_data_1;
reg [127:0] io_writeback_15_bits_data_2;
reg [6:0]   io_writeback_15_bits_pdest;
reg         io_writeback_15_bits_robIdx_flag;
reg [7:0]   io_writeback_15_bits_robIdx_value;
reg         io_writeback_15_bits_vecWen;
reg         io_writeback_15_bits_v0Wen;
reg [4:0]   io_writeback_15_bits_fflags;
reg         io_writeback_15_bits_wflags;
reg         io_writeback_15_bits_vxsat;
reg         io_writeback_15_bits_debugInfo_eliminatedMove;
reg [63:0]  io_writeback_15_bits_debugInfo_renameTime;
reg [63:0]  io_writeback_15_bits_debugInfo_dispatchTime;
reg [63:0]  io_writeback_15_bits_debugInfo_enqRsTime;
reg [63:0]  io_writeback_15_bits_debugInfo_selectTime;
reg [63:0]  io_writeback_15_bits_debugInfo_issueTime;
reg [63:0]  io_writeback_15_bits_debugInfo_writebackTime;
reg [63:0]  io_writeback_15_bits_debugInfo_runahead_checkpoint_id;
reg [63:0]  io_writeback_15_bits_debugInfo_tlbFirstReqTime;
reg [63:0]  io_writeback_15_bits_debugInfo_tlbRespTime;
reg [63:0]  io_writeback_15_bits_debug_seqNum;
reg         io_writeback_14_valid  ;
reg [127:0] io_writeback_14_bits_data_0;
reg [127:0] io_writeback_14_bits_data_1;
reg [127:0] io_writeback_14_bits_data_2;
reg [127:0] io_writeback_14_bits_data_3;
reg [127:0] io_writeback_14_bits_data_4;
reg [127:0] io_writeback_14_bits_data_5;
reg [7:0]   io_writeback_14_bits_pdest;
reg         io_writeback_14_bits_robIdx_flag;
reg [7:0]   io_writeback_14_bits_robIdx_value;
reg         io_writeback_14_bits_intWen;
reg         io_writeback_14_bits_fpWen;
reg         io_writeback_14_bits_vecWen;
reg         io_writeback_14_bits_v0Wen;
reg         io_writeback_14_bits_vlWen;
reg [4:0]   io_writeback_14_bits_fflags;
reg         io_writeback_14_bits_wflags;
reg         io_writeback_14_bits_exceptionVec_2;
reg         io_writeback_14_bits_debugInfo_eliminatedMove;
reg [63:0]  io_writeback_14_bits_debugInfo_renameTime;
reg [63:0]  io_writeback_14_bits_debugInfo_dispatchTime;
reg [63:0]  io_writeback_14_bits_debugInfo_enqRsTime;
reg [63:0]  io_writeback_14_bits_debugInfo_selectTime;
reg [63:0]  io_writeback_14_bits_debugInfo_issueTime;
reg [63:0]  io_writeback_14_bits_debugInfo_writebackTime;
reg [63:0]  io_writeback_14_bits_debugInfo_runahead_checkpoint_id;
reg [63:0]  io_writeback_14_bits_debugInfo_tlbFirstReqTime;
reg [63:0]  io_writeback_14_bits_debugInfo_tlbRespTime;
reg [63:0]  io_writeback_14_bits_debug_seqNum;
reg         io_writeback_13_valid  ;
reg [127:0] io_writeback_13_bits_data_0;
reg [127:0] io_writeback_13_bits_data_1;
reg [127:0] io_writeback_13_bits_data_2;
reg [6:0]   io_writeback_13_bits_pdest;
reg         io_writeback_13_bits_robIdx_flag;
reg [7:0]   io_writeback_13_bits_robIdx_value;
reg         io_writeback_13_bits_vecWen;
reg         io_writeback_13_bits_v0Wen;
reg [4:0]   io_writeback_13_bits_fflags;
reg         io_writeback_13_bits_wflags;
reg         io_writeback_13_bits_vxsat;
reg         io_writeback_13_bits_exceptionVec_2;
reg         io_writeback_13_bits_debugInfo_eliminatedMove;
reg [63:0]  io_writeback_13_bits_debugInfo_renameTime;
reg [63:0]  io_writeback_13_bits_debugInfo_dispatchTime;
reg [63:0]  io_writeback_13_bits_debugInfo_enqRsTime;
reg [63:0]  io_writeback_13_bits_debugInfo_selectTime;
reg [63:0]  io_writeback_13_bits_debugInfo_issueTime;
reg [63:0]  io_writeback_13_bits_debugInfo_writebackTime;
reg [63:0]  io_writeback_13_bits_debugInfo_runahead_checkpoint_id;
reg [63:0]  io_writeback_13_bits_debugInfo_tlbFirstReqTime;
reg [63:0]  io_writeback_13_bits_debugInfo_tlbRespTime;
reg [63:0]  io_writeback_13_bits_debug_seqNum;
reg         io_writeback_7_valid   ;
reg [63:0]  io_writeback_7_bits_data_0;
reg [63:0]  io_writeback_7_bits_data_1;
reg [7:0]   io_writeback_7_bits_pdest;
reg         io_writeback_7_bits_robIdx_flag;
reg [7:0]   io_writeback_7_bits_robIdx_value;
reg         io_writeback_7_bits_intWen;
reg         io_writeback_7_bits_redirect_valid;
reg         io_writeback_7_bits_redirect_bits_isRVC;
reg         io_writeback_7_bits_redirect_bits_robIdx_flag;
reg [7:0]   io_writeback_7_bits_redirect_bits_robIdx_value;
reg         io_writeback_7_bits_redirect_bits_ftqIdx_flag;
reg [5:0]   io_writeback_7_bits_redirect_bits_ftqIdx_value;
reg [3:0]   io_writeback_7_bits_redirect_bits_ftqOffset;
reg         io_writeback_7_bits_redirect_bits_level;
reg         io_writeback_7_bits_redirect_bits_interrupt;
reg [49:0]  io_writeback_7_bits_redirect_bits_cfiUpdate_pc;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC;
reg [1:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet;
reg [3:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_ssp;
reg [2:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_sctr;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag;
reg [4:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag;
reg [4:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag;
reg [4:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value;
reg [49:0]  io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr;
reg [10:0]  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist;
reg [10:0]  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist;
reg [6:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist;
reg [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist;
reg [8:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist;
reg [3:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist;
reg [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist;
reg [8:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist;
reg [6:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist;
reg [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist;
reg [6:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist;
reg [8:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist;
reg [6:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist;
reg [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist;
reg [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist;
reg [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist;
reg [10:0]  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist;
reg [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3;
reg [2:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH;
reg [3:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_ghr;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag;
reg [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value;
reg [9:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0;
reg [9:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken;
reg [49:0]  io_writeback_7_bits_redirect_bits_cfiUpdate_target;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_taken;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred;
reg [1:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_shift;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF;
reg         io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF;
reg [63:0]  io_writeback_7_bits_redirect_bits_fullTarget;
reg         io_writeback_7_bits_redirect_bits_stFtqIdx_flag;
reg [5:0]   io_writeback_7_bits_redirect_bits_stFtqIdx_value;
reg [3:0]   io_writeback_7_bits_redirect_bits_stFtqOffset;
reg [63:0]  io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id;
reg         io_writeback_7_bits_redirect_bits_debugIsCtrl;
reg         io_writeback_7_bits_redirect_bits_debugIsMemVio;
reg         io_writeback_7_bits_exceptionVec_2;
reg         io_writeback_7_bits_exceptionVec_3;
reg         io_writeback_7_bits_exceptionVec_8;
reg         io_writeback_7_bits_exceptionVec_9;
reg         io_writeback_7_bits_exceptionVec_10;
reg         io_writeback_7_bits_exceptionVec_11;
reg         io_writeback_7_bits_exceptionVec_22;
reg         io_writeback_7_bits_flushPipe;
reg         io_writeback_7_bits_predecodeInfo_valid;
reg         io_writeback_7_bits_predecodeInfo_isRVC;
reg [1:0]   io_writeback_7_bits_predecodeInfo_brType;
reg         io_writeback_7_bits_predecodeInfo_isCall;
reg         io_writeback_7_bits_predecodeInfo_isRet;
reg         io_writeback_7_bits_debug_isPerfCnt;
reg         io_writeback_7_bits_debugInfo_eliminatedMove;
reg [63:0]  io_writeback_7_bits_debugInfo_renameTime;
reg [63:0]  io_writeback_7_bits_debugInfo_dispatchTime;
reg [63:0]  io_writeback_7_bits_debugInfo_enqRsTime;
reg [63:0]  io_writeback_7_bits_debugInfo_selectTime;
reg [63:0]  io_writeback_7_bits_debugInfo_issueTime;
reg [63:0]  io_writeback_7_bits_debugInfo_writebackTime;
reg [63:0]  io_writeback_7_bits_debugInfo_runahead_checkpoint_id;
reg [63:0]  io_writeback_7_bits_debugInfo_tlbFirstReqTime;
reg [63:0]  io_writeback_7_bits_debugInfo_tlbRespTime;
reg [63:0]  io_writeback_7_bits_debug_seqNum;
reg         io_writeback_5_valid   ;
reg         io_writeback_5_bits_redirect_valid;
reg         io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred;
reg         io_writeback_3_valid   ;
reg         io_writeback_3_bits_redirect_valid;
reg         io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred;
reg         io_writeback_1_valid   ;
reg         io_writeback_1_bits_redirect_valid;
reg         io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred;
reg         io_exuWriteback_26_valid;
reg [7:0]   io_exuWriteback_26_bits_robIdx_value;
reg         io_exuWriteback_25_valid;
reg [7:0]   io_exuWriteback_25_bits_robIdx_value;
reg         io_exuWriteback_24_valid;
reg [127:0] io_exuWriteback_24_bits_data_0;
reg [6:0]   io_exuWriteback_24_bits_pdest;
reg [7:0]   io_exuWriteback_24_bits_robIdx_value;
reg         io_exuWriteback_24_bits_vecWen;
reg         io_exuWriteback_24_bits_v0Wen;
reg [2:0]   io_exuWriteback_24_bits_vls_vdIdx;
reg         io_exuWriteback_24_bits_debug_isMMIO;
reg         io_exuWriteback_24_bits_debug_isNCIO;
reg         io_exuWriteback_24_bits_debug_isPerfCnt;
reg [47:0]  io_exuWriteback_24_bits_debug_paddr;
reg         io_exuWriteback_23_valid;
reg [127:0] io_exuWriteback_23_bits_data_0;
reg [6:0]   io_exuWriteback_23_bits_pdest;
reg [7:0]   io_exuWriteback_23_bits_robIdx_value;
reg         io_exuWriteback_23_bits_vecWen;
reg         io_exuWriteback_23_bits_v0Wen;
reg [2:0]   io_exuWriteback_23_bits_vls_vdIdx;
reg         io_exuWriteback_23_bits_debug_isMMIO;
reg         io_exuWriteback_23_bits_debug_isNCIO;
reg         io_exuWriteback_23_bits_debug_isPerfCnt;
reg [47:0]  io_exuWriteback_23_bits_debug_paddr;
reg         io_exuWriteback_22_valid;
reg [63:0]  io_exuWriteback_22_bits_data_0;
reg [7:0]   io_exuWriteback_22_bits_robIdx_value;
reg [6:0]   io_exuWriteback_22_bits_lqIdx_value;
reg         io_exuWriteback_22_bits_debug_isMMIO;
reg         io_exuWriteback_22_bits_debug_isNCIO;
reg         io_exuWriteback_22_bits_debug_isPerfCnt;
reg [47:0]  io_exuWriteback_22_bits_debug_paddr;
reg         io_exuWriteback_21_valid;
reg [63:0]  io_exuWriteback_21_bits_data_0;
reg [7:0]   io_exuWriteback_21_bits_robIdx_value;
reg [6:0]   io_exuWriteback_21_bits_lqIdx_value;
reg         io_exuWriteback_21_bits_debug_isMMIO;
reg         io_exuWriteback_21_bits_debug_isNCIO;
reg         io_exuWriteback_21_bits_debug_isPerfCnt;
reg [47:0]  io_exuWriteback_21_bits_debug_paddr;
reg         io_exuWriteback_20_valid;
reg [63:0]  io_exuWriteback_20_bits_data_0;
reg [7:0]   io_exuWriteback_20_bits_robIdx_value;
reg [6:0]   io_exuWriteback_20_bits_lqIdx_value;
reg         io_exuWriteback_20_bits_debug_isMMIO;
reg         io_exuWriteback_20_bits_debug_isNCIO;
reg         io_exuWriteback_20_bits_debug_isPerfCnt;
reg [47:0]  io_exuWriteback_20_bits_debug_paddr;
reg         io_exuWriteback_19_valid;
reg [63:0]  io_exuWriteback_19_bits_data_0;
reg [7:0]   io_exuWriteback_19_bits_robIdx_value;
reg [5:0]   io_exuWriteback_19_bits_sqIdx_value;
reg         io_exuWriteback_19_bits_debug_isMMIO;
reg         io_exuWriteback_19_bits_debug_isNCIO;
reg         io_exuWriteback_19_bits_debug_isPerfCnt;
reg [47:0]  io_exuWriteback_19_bits_debug_paddr;
reg         io_exuWriteback_18_valid;
reg [63:0]  io_exuWriteback_18_bits_data_0;
reg [7:0]   io_exuWriteback_18_bits_robIdx_value;
reg [5:0]   io_exuWriteback_18_bits_sqIdx_value;
reg         io_exuWriteback_18_bits_debug_isMMIO;
reg         io_exuWriteback_18_bits_debug_isNCIO;
reg         io_exuWriteback_18_bits_debug_isPerfCnt;
reg [47:0]  io_exuWriteback_18_bits_debug_paddr;
reg         io_exuWriteback_17_valid;
reg [127:0] io_exuWriteback_17_bits_data_0;
reg [7:0]   io_exuWriteback_17_bits_robIdx_value;
reg [4:0]   io_exuWriteback_17_bits_fflags;
reg         io_exuWriteback_17_bits_wflags;
reg         io_exuWriteback_16_valid;
reg [127:0] io_exuWriteback_16_bits_data_0;
reg [7:0]   io_exuWriteback_16_bits_robIdx_value;
reg [4:0]   io_exuWriteback_16_bits_fflags;
reg         io_exuWriteback_16_bits_wflags;
reg         io_exuWriteback_15_valid;
reg [127:0] io_exuWriteback_15_bits_data_0;
reg [7:0]   io_exuWriteback_15_bits_robIdx_value;
reg [4:0]   io_exuWriteback_15_bits_fflags;
reg         io_exuWriteback_15_bits_wflags;
reg         io_exuWriteback_15_bits_vxsat;
reg         io_exuWriteback_14_valid;
reg [127:0] io_exuWriteback_14_bits_data_0;
reg [7:0]   io_exuWriteback_14_bits_robIdx_value;
reg [4:0]   io_exuWriteback_14_bits_fflags;
reg         io_exuWriteback_14_bits_wflags;
reg         io_exuWriteback_13_valid;
reg [127:0] io_exuWriteback_13_bits_data_0;
reg [7:0]   io_exuWriteback_13_bits_robIdx_value;
reg [4:0]   io_exuWriteback_13_bits_fflags;
reg         io_exuWriteback_13_bits_wflags;
reg         io_exuWriteback_13_bits_vxsat;
reg         io_exuWriteback_12_valid;
reg [63:0]  io_exuWriteback_12_bits_data_0;
reg [7:0]   io_exuWriteback_12_bits_robIdx_value;
reg [4:0]   io_exuWriteback_12_bits_fflags;
reg         io_exuWriteback_12_bits_wflags;
reg         io_exuWriteback_11_valid;
reg [63:0]  io_exuWriteback_11_bits_data_0;
reg [7:0]   io_exuWriteback_11_bits_robIdx_value;
reg [4:0]   io_exuWriteback_11_bits_fflags;
reg         io_exuWriteback_11_bits_wflags;
reg         io_exuWriteback_10_valid;
reg [63:0]  io_exuWriteback_10_bits_data_0;
reg [7:0]   io_exuWriteback_10_bits_robIdx_value;
reg [4:0]   io_exuWriteback_10_bits_fflags;
reg         io_exuWriteback_10_bits_wflags;
reg         io_exuWriteback_9_valid;
reg [63:0]  io_exuWriteback_9_bits_data_0;
reg [7:0]   io_exuWriteback_9_bits_robIdx_value;
reg [4:0]   io_exuWriteback_9_bits_fflags;
reg         io_exuWriteback_9_bits_wflags;
reg         io_exuWriteback_8_valid;
reg [127:0] io_exuWriteback_8_bits_data_0;
reg [7:0]   io_exuWriteback_8_bits_robIdx_value;
reg [4:0]   io_exuWriteback_8_bits_fflags;
reg         io_exuWriteback_8_bits_wflags;
reg         io_exuWriteback_7_valid;
reg [63:0]  io_exuWriteback_7_bits_data_0;
reg [7:0]   io_exuWriteback_7_bits_robIdx_value;
reg         io_exuWriteback_7_bits_debug_isPerfCnt;
reg         io_exuWriteback_6_valid;
reg [63:0]  io_exuWriteback_6_bits_data_0;
reg [7:0]   io_exuWriteback_6_bits_robIdx_value;
reg         io_exuWriteback_5_valid;
reg [127:0] io_exuWriteback_5_bits_data_0;
reg [7:0]   io_exuWriteback_5_bits_robIdx_value;
reg         io_exuWriteback_5_bits_redirect_valid;
reg         io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken;
reg [4:0]   io_exuWriteback_5_bits_fflags;
reg         io_exuWriteback_5_bits_wflags;
reg         io_exuWriteback_4_valid;
reg [63:0]  io_exuWriteback_4_bits_data_0;
reg [7:0]   io_exuWriteback_4_bits_robIdx_value;
reg         io_exuWriteback_3_valid;
reg [63:0]  io_exuWriteback_3_bits_data_0;
reg [7:0]   io_exuWriteback_3_bits_robIdx_value;
reg         io_exuWriteback_3_bits_redirect_valid;
reg         io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken;
reg         io_exuWriteback_2_valid;
reg [63:0]  io_exuWriteback_2_bits_data_0;
reg [7:0]   io_exuWriteback_2_bits_robIdx_value;
reg         io_exuWriteback_1_valid;
reg [63:0]  io_exuWriteback_1_bits_data_0;
reg [7:0]   io_exuWriteback_1_bits_robIdx_value;
reg         io_exuWriteback_1_bits_redirect_valid;
reg         io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken;
reg         io_exuWriteback_0_valid;
reg [63:0]  io_exuWriteback_0_bits_data_0;
reg [7:0]   io_exuWriteback_0_bits_robIdx_value;
reg [4:0]   io_writebackNums_0_bits;
reg [4:0]   io_writebackNums_1_bits;
reg [4:0]   io_writebackNums_2_bits;
reg [4:0]   io_writebackNums_3_bits;
reg [4:0]   io_writebackNums_4_bits;
reg [4:0]   io_writebackNums_5_bits;
reg [4:0]   io_writebackNums_6_bits;
reg [4:0]   io_writebackNums_7_bits;
reg [4:0]   io_writebackNums_8_bits;
reg [4:0]   io_writebackNums_9_bits;
reg [4:0]   io_writebackNums_10_bits;
reg [4:0]   io_writebackNums_11_bits;
reg [4:0]   io_writebackNums_12_bits;
reg [4:0]   io_writebackNums_13_bits;
reg [4:0]   io_writebackNums_14_bits;
reg [4:0]   io_writebackNums_15_bits;
reg [4:0]   io_writebackNums_16_bits;
reg [4:0]   io_writebackNums_17_bits;
reg [4:0]   io_writebackNums_18_bits;
reg [4:0]   io_writebackNums_19_bits;
reg [4:0]   io_writebackNums_20_bits;
reg [4:0]   io_writebackNums_21_bits;
reg [4:0]   io_writebackNums_22_bits;
reg [4:0]   io_writebackNums_23_bits;
reg [4:0]   io_writebackNums_24_bits;
reg         io_writebackNeedFlush_0;
reg         io_writebackNeedFlush_1;
reg         io_writebackNeedFlush_2;
reg         io_writebackNeedFlush_6;
reg         io_writebackNeedFlush_7;
reg         io_writebackNeedFlush_8;
reg         io_writebackNeedFlush_9;
reg         io_writebackNeedFlush_10;
reg         io_writebackNeedFlush_11;
reg         io_writebackNeedFlush_12;
//Redirect_in
reg         io_redirect_valid      ;
reg         io_redirect_bits_robIdx_flag;
reg [7:0]   io_redirect_bits_robIdx_value;
reg         io_redirect_bits_level ;
//CSR_in
reg         io_csr_intrBitSet      ;
reg         io_csr_wfiEvent        ;
reg         io_csr_criticalErrorState;
reg         io_snpt_snptDeq        ;
reg         io_snpt_useSnpt        ;
reg [1:0]   io_snpt_snptSelect     ;
reg         io_snpt_flushVec_0     ;
reg         io_snpt_flushVec_1     ;
reg         io_snpt_flushVec_2     ;
reg         io_snpt_flushVec_3     ;
reg         io_wfi_safeFromMem     ;
reg         io_wfi_safeFromFrontend;
reg         io_wfi_enable          ;
reg         io_fromVecExcpMod_busy ;
reg [55:0]  io_readGPAMemData_gpaddr;
reg         io_readGPAMemData_isForVSnonLeafPTE;
reg         io_vstartIsZero        ;
reg         io_debugEnqLsq_canAccept;
reg [1:0]   io_debugEnqLsq_needAlloc_0;
reg [1:0]   io_debugEnqLsq_needAlloc_1;
reg [1:0]   io_debugEnqLsq_needAlloc_2;
reg [1:0]   io_debugEnqLsq_needAlloc_3;
reg [1:0]   io_debugEnqLsq_needAlloc_4;
reg [1:0]   io_debugEnqLsq_needAlloc_5;
reg         io_debugEnqLsq_req_0_valid;
reg [7:0]   io_debugEnqLsq_req_0_bits_robIdx_value;
reg [6:0]   io_debugEnqLsq_req_0_bits_lqIdx_value;
reg         io_debugEnqLsq_req_1_valid;
reg [7:0]   io_debugEnqLsq_req_1_bits_robIdx_value;
reg [6:0]   io_debugEnqLsq_req_1_bits_lqIdx_value;
reg         io_debugEnqLsq_req_2_valid;
reg [7:0]   io_debugEnqLsq_req_2_bits_robIdx_value;
reg [6:0]   io_debugEnqLsq_req_2_bits_lqIdx_value;
reg         io_debugEnqLsq_req_3_valid;
reg [7:0]   io_debugEnqLsq_req_3_bits_robIdx_value;
reg [6:0]   io_debugEnqLsq_req_3_bits_lqIdx_value;
reg         io_debugEnqLsq_req_4_valid;
reg [7:0]   io_debugEnqLsq_req_4_bits_robIdx_value;
reg [6:0]   io_debugEnqLsq_req_4_bits_lqIdx_value;
reg         io_debugEnqLsq_req_5_valid;
reg [7:0]   io_debugEnqLsq_req_5_bits_robIdx_value;
reg [6:0]   io_debugEnqLsq_req_5_bits_lqIdx_value;
reg         io_debugInstrAddrTransType_bare;
reg         io_debugInstrAddrTransType_sv39;
reg         io_debugInstrAddrTransType_sv39x4;
reg         io_debugInstrAddrTransType_sv48;
reg         io_debugInstrAddrTransType_sv48x4;
reg [7:0]   io_storeDebugInfo_0_robidx_value;
reg [7:0]   io_storeDebugInfo_1_robidx_value;
//Mem_in
reg         io_lsq_mmio_0          ;
reg         io_lsq_mmio_1          ;
reg         io_lsq_mmio_2          ;
reg [7:0]   io_lsq_uop_0_robIdx_value;
reg [7:0]   io_lsq_uop_1_robIdx_value;
reg [7:0]   io_lsq_uop_2_robIdx_value;
//Rob_output
wire         io_enq_canAccept      ;
wire         io_enq_canAcceptForDispatch;
wire         io_enq_isEmpty        ;
wire         io_flushOut_valid     ;
wire         io_flushOut_bits_isRVC;
wire         io_flushOut_bits_robIdx_flag;
wire [7:0]   io_flushOut_bits_robIdx_value;
wire         io_flushOut_bits_ftqIdx_flag;
wire [5:0]   io_flushOut_bits_ftqIdx_value;
wire [3:0]   io_flushOut_bits_ftqOffset;
wire         io_flushOut_bits_level;
wire         io_exception_valid    ;
wire [31:0]  io_exception_bits_instr;
wire [2:0]   io_exception_bits_commitType;
wire         io_exception_bits_exceptionVec_0;
wire         io_exception_bits_exceptionVec_1;
wire         io_exception_bits_exceptionVec_2;
wire         io_exception_bits_exceptionVec_3;
wire         io_exception_bits_exceptionVec_4;
wire         io_exception_bits_exceptionVec_5;
wire         io_exception_bits_exceptionVec_6;
wire         io_exception_bits_exceptionVec_7;
wire         io_exception_bits_exceptionVec_8;
wire         io_exception_bits_exceptionVec_9;
wire         io_exception_bits_exceptionVec_10;
wire         io_exception_bits_exceptionVec_11;
wire         io_exception_bits_exceptionVec_12;
wire         io_exception_bits_exceptionVec_13;
wire         io_exception_bits_exceptionVec_14;
wire         io_exception_bits_exceptionVec_15;
wire         io_exception_bits_exceptionVec_16;
wire         io_exception_bits_exceptionVec_17;
wire         io_exception_bits_exceptionVec_18;
wire         io_exception_bits_exceptionVec_19;
wire         io_exception_bits_exceptionVec_20;
wire         io_exception_bits_exceptionVec_21;
wire         io_exception_bits_exceptionVec_22;
wire         io_exception_bits_exceptionVec_23;
wire         io_exception_bits_isPcBkpt;
wire         io_exception_bits_isFetchMalAddr;
wire [63:0]  io_exception_bits_gpaddr;
wire         io_exception_bits_singleStep;
wire         io_exception_bits_crossPageIPFFix;
wire         io_exception_bits_isInterrupt;
wire         io_exception_bits_isHls;
wire [3:0]   io_exception_bits_trigger;
wire         io_exception_bits_isForVSnonLeafPTE;
wire         io_commits_isCommit   ;
wire         io_commits_commitValid_0;
wire         io_commits_commitValid_1;
wire         io_commits_commitValid_2;
wire         io_commits_commitValid_3;
wire         io_commits_commitValid_4;
wire         io_commits_commitValid_5;
wire         io_commits_commitValid_6;
wire         io_commits_commitValid_7;
wire         io_commits_isWalk     ;
wire         io_commits_walkValid_0;
wire         io_commits_walkValid_1;
wire         io_commits_walkValid_2;
wire         io_commits_walkValid_3;
wire         io_commits_walkValid_4;
wire         io_commits_walkValid_5;
wire         io_commits_walkValid_6;
wire         io_commits_walkValid_7;
wire         io_commits_info_0_walk_v;
wire         io_commits_info_0_commit_v;
wire         io_commits_info_0_commit_w;
wire [6:0]   io_commits_info_0_realDestSize;
wire         io_commits_info_0_interrupt_safe;
wire         io_commits_info_0_wflags;
wire [4:0]   io_commits_info_0_fflags;
wire         io_commits_info_0_vxsat;
wire         io_commits_info_0_isRVC;
wire         io_commits_info_0_isVset;
wire         io_commits_info_0_isHls;
wire         io_commits_info_0_isVls;
wire         io_commits_info_0_vls ;
wire         io_commits_info_0_mmio;
wire [2:0]   io_commits_info_0_commitType;
wire         io_commits_info_0_ftqIdx_flag;
wire [5:0]   io_commits_info_0_ftqIdx_value;
wire [3:0]   io_commits_info_0_ftqOffset;
wire [2:0]   io_commits_info_0_instrSize;
wire         io_commits_info_0_fpWen;
wire         io_commits_info_0_rfWen;
wire         io_commits_info_0_needFlush;
wire [3:0]   io_commits_info_0_traceBlockInPipe_itype;
wire [3:0]   io_commits_info_0_traceBlockInPipe_iretire;
wire         io_commits_info_0_traceBlockInPipe_ilastsize;
wire [49:0]  io_commits_info_0_debug_pc;
wire [31:0]  io_commits_info_0_debug_instr;
wire [5:0]   io_commits_info_0_debug_ldest;
wire [7:0]   io_commits_info_0_debug_pdest;
wire [7:0]   io_commits_info_0_debug_otherPdest_0;
wire [7:0]   io_commits_info_0_debug_otherPdest_1;
wire [7:0]   io_commits_info_0_debug_otherPdest_2;
wire [7:0]   io_commits_info_0_debug_otherPdest_3;
wire [7:0]   io_commits_info_0_debug_otherPdest_4;
wire [7:0]   io_commits_info_0_debug_otherPdest_5;
wire [7:0]   io_commits_info_0_debug_otherPdest_6;
wire [34:0]  io_commits_info_0_debug_fuType;
wire         io_commits_info_0_dirtyFs;
wire         io_commits_info_0_dirtyVs;
wire         io_commits_info_1_walk_v;
wire         io_commits_info_1_commit_v;
wire         io_commits_info_1_commit_w;
wire [6:0]   io_commits_info_1_realDestSize;
wire         io_commits_info_1_interrupt_safe;
wire         io_commits_info_1_wflags;
wire [4:0]   io_commits_info_1_fflags;
wire         io_commits_info_1_vxsat;
wire         io_commits_info_1_isRVC;
wire         io_commits_info_1_isVset;
wire         io_commits_info_1_isHls;
wire         io_commits_info_1_isVls;
wire         io_commits_info_1_vls ;
wire         io_commits_info_1_mmio;
wire [2:0]   io_commits_info_1_commitType;
wire         io_commits_info_1_ftqIdx_flag;
wire [5:0]   io_commits_info_1_ftqIdx_value;
wire [3:0]   io_commits_info_1_ftqOffset;
wire [2:0]   io_commits_info_1_instrSize;
wire         io_commits_info_1_fpWen;
wire         io_commits_info_1_rfWen;
wire         io_commits_info_1_needFlush;
wire [3:0]   io_commits_info_1_traceBlockInPipe_itype;
wire [3:0]   io_commits_info_1_traceBlockInPipe_iretire;
wire         io_commits_info_1_traceBlockInPipe_ilastsize;
wire [49:0]  io_commits_info_1_debug_pc;
wire [31:0]  io_commits_info_1_debug_instr;
wire [5:0]   io_commits_info_1_debug_ldest;
wire [7:0]   io_commits_info_1_debug_pdest;
wire [7:0]   io_commits_info_1_debug_otherPdest_0;
wire [7:0]   io_commits_info_1_debug_otherPdest_1;
wire [7:0]   io_commits_info_1_debug_otherPdest_2;
wire [7:0]   io_commits_info_1_debug_otherPdest_3;
wire [7:0]   io_commits_info_1_debug_otherPdest_4;
wire [7:0]   io_commits_info_1_debug_otherPdest_5;
wire [7:0]   io_commits_info_1_debug_otherPdest_6;
wire [34:0]  io_commits_info_1_debug_fuType;
wire         io_commits_info_1_dirtyFs;
wire         io_commits_info_1_dirtyVs;
wire         io_commits_info_2_walk_v;
wire         io_commits_info_2_commit_v;
wire         io_commits_info_2_commit_w;
wire [6:0]   io_commits_info_2_realDestSize;
wire         io_commits_info_2_interrupt_safe;
wire         io_commits_info_2_wflags;
wire [4:0]   io_commits_info_2_fflags;
wire         io_commits_info_2_vxsat;
wire         io_commits_info_2_isRVC;
wire         io_commits_info_2_isVset;
wire         io_commits_info_2_isHls;
wire         io_commits_info_2_isVls;
wire         io_commits_info_2_vls ;
wire         io_commits_info_2_mmio;
wire [2:0]   io_commits_info_2_commitType;
wire         io_commits_info_2_ftqIdx_flag;
wire [5:0]   io_commits_info_2_ftqIdx_value;
wire [3:0]   io_commits_info_2_ftqOffset;
wire [2:0]   io_commits_info_2_instrSize;
wire         io_commits_info_2_fpWen;
wire         io_commits_info_2_rfWen;
wire         io_commits_info_2_needFlush;
wire [3:0]   io_commits_info_2_traceBlockInPipe_itype;
wire [3:0]   io_commits_info_2_traceBlockInPipe_iretire;
wire         io_commits_info_2_traceBlockInPipe_ilastsize;
wire [49:0]  io_commits_info_2_debug_pc;
wire [31:0]  io_commits_info_2_debug_instr;
wire [5:0]   io_commits_info_2_debug_ldest;
wire [7:0]   io_commits_info_2_debug_pdest;
wire [7:0]   io_commits_info_2_debug_otherPdest_0;
wire [7:0]   io_commits_info_2_debug_otherPdest_1;
wire [7:0]   io_commits_info_2_debug_otherPdest_2;
wire [7:0]   io_commits_info_2_debug_otherPdest_3;
wire [7:0]   io_commits_info_2_debug_otherPdest_4;
wire [7:0]   io_commits_info_2_debug_otherPdest_5;
wire [7:0]   io_commits_info_2_debug_otherPdest_6;
wire [34:0]  io_commits_info_2_debug_fuType;
wire         io_commits_info_2_dirtyFs;
wire         io_commits_info_2_dirtyVs;
wire         io_commits_info_3_walk_v;
wire         io_commits_info_3_commit_v;
wire         io_commits_info_3_commit_w;
wire [6:0]   io_commits_info_3_realDestSize;
wire         io_commits_info_3_interrupt_safe;
wire         io_commits_info_3_wflags;
wire [4:0]   io_commits_info_3_fflags;
wire         io_commits_info_3_vxsat;
wire         io_commits_info_3_isRVC;
wire         io_commits_info_3_isVset;
wire         io_commits_info_3_isHls;
wire         io_commits_info_3_isVls;
wire         io_commits_info_3_vls ;
wire         io_commits_info_3_mmio;
wire [2:0]   io_commits_info_3_commitType;
wire         io_commits_info_3_ftqIdx_flag;
wire [5:0]   io_commits_info_3_ftqIdx_value;
wire [3:0]   io_commits_info_3_ftqOffset;
wire [2:0]   io_commits_info_3_instrSize;
wire         io_commits_info_3_fpWen;
wire         io_commits_info_3_rfWen;
wire         io_commits_info_3_needFlush;
wire [3:0]   io_commits_info_3_traceBlockInPipe_itype;
wire [3:0]   io_commits_info_3_traceBlockInPipe_iretire;
wire         io_commits_info_3_traceBlockInPipe_ilastsize;
wire [49:0]  io_commits_info_3_debug_pc;
wire [31:0]  io_commits_info_3_debug_instr;
wire [5:0]   io_commits_info_3_debug_ldest;
wire [7:0]   io_commits_info_3_debug_pdest;
wire [7:0]   io_commits_info_3_debug_otherPdest_0;
wire [7:0]   io_commits_info_3_debug_otherPdest_1;
wire [7:0]   io_commits_info_3_debug_otherPdest_2;
wire [7:0]   io_commits_info_3_debug_otherPdest_3;
wire [7:0]   io_commits_info_3_debug_otherPdest_4;
wire [7:0]   io_commits_info_3_debug_otherPdest_5;
wire [7:0]   io_commits_info_3_debug_otherPdest_6;
wire [34:0]  io_commits_info_3_debug_fuType;
wire         io_commits_info_3_dirtyFs;
wire         io_commits_info_3_dirtyVs;
wire         io_commits_info_4_walk_v;
wire         io_commits_info_4_commit_v;
wire         io_commits_info_4_commit_w;
wire [6:0]   io_commits_info_4_realDestSize;
wire         io_commits_info_4_interrupt_safe;
wire         io_commits_info_4_wflags;
wire [4:0]   io_commits_info_4_fflags;
wire         io_commits_info_4_vxsat;
wire         io_commits_info_4_isRVC;
wire         io_commits_info_4_isVset;
wire         io_commits_info_4_isHls;
wire         io_commits_info_4_isVls;
wire         io_commits_info_4_vls ;
wire         io_commits_info_4_mmio;
wire [2:0]   io_commits_info_4_commitType;
wire         io_commits_info_4_ftqIdx_flag;
wire [5:0]   io_commits_info_4_ftqIdx_value;
wire [3:0]   io_commits_info_4_ftqOffset;
wire [2:0]   io_commits_info_4_instrSize;
wire         io_commits_info_4_fpWen;
wire         io_commits_info_4_rfWen;
wire         io_commits_info_4_needFlush;
wire [3:0]   io_commits_info_4_traceBlockInPipe_itype;
wire [3:0]   io_commits_info_4_traceBlockInPipe_iretire;
wire         io_commits_info_4_traceBlockInPipe_ilastsize;
wire [49:0]  io_commits_info_4_debug_pc;
wire [31:0]  io_commits_info_4_debug_instr;
wire [5:0]   io_commits_info_4_debug_ldest;
wire [7:0]   io_commits_info_4_debug_pdest;
wire [7:0]   io_commits_info_4_debug_otherPdest_0;
wire [7:0]   io_commits_info_4_debug_otherPdest_1;
wire [7:0]   io_commits_info_4_debug_otherPdest_2;
wire [7:0]   io_commits_info_4_debug_otherPdest_3;
wire [7:0]   io_commits_info_4_debug_otherPdest_4;
wire [7:0]   io_commits_info_4_debug_otherPdest_5;
wire [7:0]   io_commits_info_4_debug_otherPdest_6;
wire [34:0]  io_commits_info_4_debug_fuType;
wire         io_commits_info_4_dirtyFs;
wire         io_commits_info_4_dirtyVs;
wire         io_commits_info_5_walk_v;
wire         io_commits_info_5_commit_v;
wire         io_commits_info_5_commit_w;
wire [6:0]   io_commits_info_5_realDestSize;
wire         io_commits_info_5_interrupt_safe;
wire         io_commits_info_5_wflags;
wire [4:0]   io_commits_info_5_fflags;
wire         io_commits_info_5_vxsat;
wire         io_commits_info_5_isRVC;
wire         io_commits_info_5_isVset;
wire         io_commits_info_5_isHls;
wire         io_commits_info_5_isVls;
wire         io_commits_info_5_vls ;
wire         io_commits_info_5_mmio;
wire [2:0]   io_commits_info_5_commitType;
wire         io_commits_info_5_ftqIdx_flag;
wire [5:0]   io_commits_info_5_ftqIdx_value;
wire [3:0]   io_commits_info_5_ftqOffset;
wire [2:0]   io_commits_info_5_instrSize;
wire         io_commits_info_5_fpWen;
wire         io_commits_info_5_rfWen;
wire         io_commits_info_5_needFlush;
wire [3:0]   io_commits_info_5_traceBlockInPipe_itype;
wire [3:0]   io_commits_info_5_traceBlockInPipe_iretire;
wire         io_commits_info_5_traceBlockInPipe_ilastsize;
wire [49:0]  io_commits_info_5_debug_pc;
wire [31:0]  io_commits_info_5_debug_instr;
wire [5:0]   io_commits_info_5_debug_ldest;
wire [7:0]   io_commits_info_5_debug_pdest;
wire [7:0]   io_commits_info_5_debug_otherPdest_0;
wire [7:0]   io_commits_info_5_debug_otherPdest_1;
wire [7:0]   io_commits_info_5_debug_otherPdest_2;
wire [7:0]   io_commits_info_5_debug_otherPdest_3;
wire [7:0]   io_commits_info_5_debug_otherPdest_4;
wire [7:0]   io_commits_info_5_debug_otherPdest_5;
wire [7:0]   io_commits_info_5_debug_otherPdest_6;
wire [34:0]  io_commits_info_5_debug_fuType;
wire         io_commits_info_5_dirtyFs;
wire         io_commits_info_5_dirtyVs;
wire         io_commits_info_6_walk_v;
wire         io_commits_info_6_commit_v;
wire         io_commits_info_6_commit_w;
wire [6:0]   io_commits_info_6_realDestSize;
wire         io_commits_info_6_interrupt_safe;
wire         io_commits_info_6_wflags;
wire [4:0]   io_commits_info_6_fflags;
wire         io_commits_info_6_vxsat;
wire         io_commits_info_6_isRVC;
wire         io_commits_info_6_isVset;
wire         io_commits_info_6_isHls;
wire         io_commits_info_6_isVls;
wire         io_commits_info_6_vls ;
wire         io_commits_info_6_mmio;
wire [2:0]   io_commits_info_6_commitType;
wire         io_commits_info_6_ftqIdx_flag;
wire [5:0]   io_commits_info_6_ftqIdx_value;
wire [3:0]   io_commits_info_6_ftqOffset;
wire [2:0]   io_commits_info_6_instrSize;
wire         io_commits_info_6_fpWen;
wire         io_commits_info_6_rfWen;
wire         io_commits_info_6_needFlush;
wire [3:0]   io_commits_info_6_traceBlockInPipe_itype;
wire [3:0]   io_commits_info_6_traceBlockInPipe_iretire;
wire         io_commits_info_6_traceBlockInPipe_ilastsize;
wire [49:0]  io_commits_info_6_debug_pc;
wire [31:0]  io_commits_info_6_debug_instr;
wire [5:0]   io_commits_info_6_debug_ldest;
wire [7:0]   io_commits_info_6_debug_pdest;
wire [7:0]   io_commits_info_6_debug_otherPdest_0;
wire [7:0]   io_commits_info_6_debug_otherPdest_1;
wire [7:0]   io_commits_info_6_debug_otherPdest_2;
wire [7:0]   io_commits_info_6_debug_otherPdest_3;
wire [7:0]   io_commits_info_6_debug_otherPdest_4;
wire [7:0]   io_commits_info_6_debug_otherPdest_5;
wire [7:0]   io_commits_info_6_debug_otherPdest_6;
wire [34:0]  io_commits_info_6_debug_fuType;
wire         io_commits_info_6_dirtyFs;
wire         io_commits_info_6_dirtyVs;
wire         io_commits_info_7_walk_v;
wire         io_commits_info_7_commit_v;
wire         io_commits_info_7_commit_w;
wire [6:0]   io_commits_info_7_realDestSize;
wire         io_commits_info_7_interrupt_safe;
wire         io_commits_info_7_wflags;
wire [4:0]   io_commits_info_7_fflags;
wire         io_commits_info_7_vxsat;
wire         io_commits_info_7_isRVC;
wire         io_commits_info_7_isVset;
wire         io_commits_info_7_isHls;
wire         io_commits_info_7_isVls;
wire         io_commits_info_7_vls ;
wire         io_commits_info_7_mmio;
wire [2:0]   io_commits_info_7_commitType;
wire         io_commits_info_7_ftqIdx_flag;
wire [5:0]   io_commits_info_7_ftqIdx_value;
wire [3:0]   io_commits_info_7_ftqOffset;
wire [2:0]   io_commits_info_7_instrSize;
wire         io_commits_info_7_fpWen;
wire         io_commits_info_7_rfWen;
wire         io_commits_info_7_needFlush;
wire [3:0]   io_commits_info_7_traceBlockInPipe_itype;
wire [3:0]   io_commits_info_7_traceBlockInPipe_iretire;
wire         io_commits_info_7_traceBlockInPipe_ilastsize;
wire [49:0]  io_commits_info_7_debug_pc;
wire [31:0]  io_commits_info_7_debug_instr;
wire [5:0]   io_commits_info_7_debug_ldest;
wire [7:0]   io_commits_info_7_debug_pdest;
wire [7:0]   io_commits_info_7_debug_otherPdest_0;
wire [7:0]   io_commits_info_7_debug_otherPdest_1;
wire [7:0]   io_commits_info_7_debug_otherPdest_2;
wire [7:0]   io_commits_info_7_debug_otherPdest_3;
wire [7:0]   io_commits_info_7_debug_otherPdest_4;
wire [7:0]   io_commits_info_7_debug_otherPdest_5;
wire [7:0]   io_commits_info_7_debug_otherPdest_6;
wire [34:0]  io_commits_info_7_debug_fuType;
wire         io_commits_info_7_dirtyFs;
wire         io_commits_info_7_dirtyVs;
wire         io_commits_robIdx_0_flag;
wire [7:0]   io_commits_robIdx_0_value;
wire         io_commits_robIdx_1_flag;
wire [7:0]   io_commits_robIdx_1_value;
wire         io_commits_robIdx_2_flag;
wire [7:0]   io_commits_robIdx_2_value;
wire         io_commits_robIdx_3_flag;
wire [7:0]   io_commits_robIdx_3_value;
wire         io_commits_robIdx_4_flag;
wire [7:0]   io_commits_robIdx_4_value;
wire         io_commits_robIdx_5_flag;
wire [7:0]   io_commits_robIdx_5_value;
wire         io_commits_robIdx_6_flag;
wire [7:0]   io_commits_robIdx_6_value;
wire         io_commits_robIdx_7_flag;
wire [7:0]   io_commits_robIdx_7_value;
reg         io_trace_blockCommit   ;
wire         io_trace_traceCommitInfo_blocks_0_valid;
wire [5:0]   io_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value;
wire [3:0]   io_trace_traceCommitInfo_blocks_0_bits_ftqOffset;
wire [3:0]   io_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype;
wire [3:0]   io_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire;
wire         io_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize;
wire         io_trace_traceCommitInfo_blocks_1_valid;
wire [5:0]   io_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value;
wire [3:0]   io_trace_traceCommitInfo_blocks_1_bits_ftqOffset;
wire [3:0]   io_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype;
wire [3:0]   io_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire;
wire         io_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize;
wire         io_trace_traceCommitInfo_blocks_2_valid;
wire [5:0]   io_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value;
wire [3:0]   io_trace_traceCommitInfo_blocks_2_bits_ftqOffset;
wire [3:0]   io_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype;
wire [3:0]   io_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire;
wire         io_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize;
wire         io_trace_traceCommitInfo_blocks_3_valid;
wire [5:0]   io_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value;
wire [3:0]   io_trace_traceCommitInfo_blocks_3_bits_ftqOffset;
wire [3:0]   io_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype;
wire [3:0]   io_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire;
wire         io_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize;
wire         io_trace_traceCommitInfo_blocks_4_valid;
wire [5:0]   io_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value;
wire [3:0]   io_trace_traceCommitInfo_blocks_4_bits_ftqOffset;
wire [3:0]   io_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype;
wire [3:0]   io_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire;
wire         io_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize;
wire         io_trace_traceCommitInfo_blocks_5_valid;
wire [5:0]   io_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value;
wire [3:0]   io_trace_traceCommitInfo_blocks_5_bits_ftqOffset;
wire [3:0]   io_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype;
wire [3:0]   io_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire;
wire         io_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize;
wire         io_trace_traceCommitInfo_blocks_6_valid;
wire [5:0]   io_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value;
wire [3:0]   io_trace_traceCommitInfo_blocks_6_bits_ftqOffset;
wire [3:0]   io_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype;
wire [3:0]   io_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire;
wire         io_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize;
wire         io_trace_traceCommitInfo_blocks_7_valid;
wire [5:0]   io_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value;
wire [3:0]   io_trace_traceCommitInfo_blocks_7_bits_ftqOffset;
wire [3:0]   io_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype;
wire [3:0]   io_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire;
wire         io_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize;
wire         io_rabCommits_isCommit;
wire         io_rabCommits_commitValid_0;
wire         io_rabCommits_commitValid_1;
wire         io_rabCommits_commitValid_2;
wire         io_rabCommits_commitValid_3;
wire         io_rabCommits_commitValid_4;
wire         io_rabCommits_commitValid_5;
wire         io_rabCommits_isWalk  ;
wire         io_rabCommits_walkValid_0;
wire         io_rabCommits_walkValid_1;
wire         io_rabCommits_walkValid_2;
wire         io_rabCommits_walkValid_3;
wire         io_rabCommits_walkValid_4;
wire         io_rabCommits_walkValid_5;
wire [5:0]   io_rabCommits_info_0_ldest;
wire [7:0]   io_rabCommits_info_0_pdest;
wire         io_rabCommits_info_0_rfWen;
wire         io_rabCommits_info_0_fpWen;
wire         io_rabCommits_info_0_vecWen;
wire         io_rabCommits_info_0_v0Wen;
wire         io_rabCommits_info_0_vlWen;
wire         io_rabCommits_info_0_isMove;
wire [5:0]   io_rabCommits_info_1_ldest;
wire [7:0]   io_rabCommits_info_1_pdest;
wire         io_rabCommits_info_1_rfWen;
wire         io_rabCommits_info_1_fpWen;
wire         io_rabCommits_info_1_vecWen;
wire         io_rabCommits_info_1_v0Wen;
wire         io_rabCommits_info_1_vlWen;
wire         io_rabCommits_info_1_isMove;
wire [5:0]   io_rabCommits_info_2_ldest;
wire [7:0]   io_rabCommits_info_2_pdest;
wire         io_rabCommits_info_2_rfWen;
wire         io_rabCommits_info_2_fpWen;
wire         io_rabCommits_info_2_vecWen;
wire         io_rabCommits_info_2_v0Wen;
wire         io_rabCommits_info_2_vlWen;
wire         io_rabCommits_info_2_isMove;
wire [5:0]   io_rabCommits_info_3_ldest;
wire [7:0]   io_rabCommits_info_3_pdest;
wire         io_rabCommits_info_3_rfWen;
wire         io_rabCommits_info_3_fpWen;
wire         io_rabCommits_info_3_vecWen;
wire         io_rabCommits_info_3_v0Wen;
wire         io_rabCommits_info_3_vlWen;
wire         io_rabCommits_info_3_isMove;
wire [5:0]   io_rabCommits_info_4_ldest;
wire [7:0]   io_rabCommits_info_4_pdest;
wire         io_rabCommits_info_4_rfWen;
wire         io_rabCommits_info_4_fpWen;
wire         io_rabCommits_info_4_vecWen;
wire         io_rabCommits_info_4_v0Wen;
wire         io_rabCommits_info_4_vlWen;
wire         io_rabCommits_info_4_isMove;
wire [5:0]   io_rabCommits_info_5_ldest;
wire [7:0]   io_rabCommits_info_5_pdest;
wire         io_rabCommits_info_5_rfWen;
wire         io_rabCommits_info_5_fpWen;
wire         io_rabCommits_info_5_vecWen;
wire         io_rabCommits_info_5_v0Wen;
wire         io_rabCommits_info_5_vlWen;
wire         io_rabCommits_info_5_isMove;
wire         io_diffCommits_commitValid_0;
wire         io_diffCommits_commitValid_1;
wire         io_diffCommits_commitValid_2;
wire         io_diffCommits_commitValid_3;
wire         io_diffCommits_commitValid_4;
wire         io_diffCommits_commitValid_5;
wire         io_diffCommits_commitValid_6;
wire         io_diffCommits_commitValid_7;
wire         io_diffCommits_commitValid_8;
wire         io_diffCommits_commitValid_9;
wire         io_diffCommits_commitValid_10;
wire         io_diffCommits_commitValid_11;
wire         io_diffCommits_commitValid_12;
wire         io_diffCommits_commitValid_13;
wire         io_diffCommits_commitValid_14;
wire         io_diffCommits_commitValid_15;
wire         io_diffCommits_commitValid_16;
wire         io_diffCommits_commitValid_17;
wire         io_diffCommits_commitValid_18;
wire         io_diffCommits_commitValid_19;
wire         io_diffCommits_commitValid_20;
wire         io_diffCommits_commitValid_21;
wire         io_diffCommits_commitValid_22;
wire         io_diffCommits_commitValid_23;
wire         io_diffCommits_commitValid_24;
wire         io_diffCommits_commitValid_25;
wire         io_diffCommits_commitValid_26;
wire         io_diffCommits_commitValid_27;
wire         io_diffCommits_commitValid_28;
wire         io_diffCommits_commitValid_29;
wire         io_diffCommits_commitValid_30;
wire         io_diffCommits_commitValid_31;
wire         io_diffCommits_commitValid_32;
wire         io_diffCommits_commitValid_33;
wire         io_diffCommits_commitValid_34;
wire         io_diffCommits_commitValid_35;
wire         io_diffCommits_commitValid_36;
wire         io_diffCommits_commitValid_37;
wire         io_diffCommits_commitValid_38;
wire         io_diffCommits_commitValid_39;
wire         io_diffCommits_commitValid_40;
wire         io_diffCommits_commitValid_41;
wire         io_diffCommits_commitValid_42;
wire         io_diffCommits_commitValid_43;
wire         io_diffCommits_commitValid_44;
wire         io_diffCommits_commitValid_45;
wire         io_diffCommits_commitValid_46;
wire         io_diffCommits_commitValid_47;
wire         io_diffCommits_commitValid_48;
wire         io_diffCommits_commitValid_49;
wire         io_diffCommits_commitValid_50;
wire         io_diffCommits_commitValid_51;
wire         io_diffCommits_commitValid_52;
wire         io_diffCommits_commitValid_53;
wire         io_diffCommits_commitValid_54;
wire         io_diffCommits_commitValid_55;
wire         io_diffCommits_commitValid_56;
wire         io_diffCommits_commitValid_57;
wire         io_diffCommits_commitValid_58;
wire         io_diffCommits_commitValid_59;
wire         io_diffCommits_commitValid_60;
wire         io_diffCommits_commitValid_61;
wire         io_diffCommits_commitValid_62;
wire         io_diffCommits_commitValid_63;
wire         io_diffCommits_commitValid_64;
wire         io_diffCommits_commitValid_65;
wire         io_diffCommits_commitValid_66;
wire         io_diffCommits_commitValid_67;
wire         io_diffCommits_commitValid_68;
wire         io_diffCommits_commitValid_69;
wire         io_diffCommits_commitValid_70;
wire         io_diffCommits_commitValid_71;
wire         io_diffCommits_commitValid_72;
wire         io_diffCommits_commitValid_73;
wire         io_diffCommits_commitValid_74;
wire         io_diffCommits_commitValid_75;
wire         io_diffCommits_commitValid_76;
wire         io_diffCommits_commitValid_77;
wire         io_diffCommits_commitValid_78;
wire         io_diffCommits_commitValid_79;
wire         io_diffCommits_commitValid_80;
wire         io_diffCommits_commitValid_81;
wire         io_diffCommits_commitValid_82;
wire         io_diffCommits_commitValid_83;
wire         io_diffCommits_commitValid_84;
wire         io_diffCommits_commitValid_85;
wire         io_diffCommits_commitValid_86;
wire         io_diffCommits_commitValid_87;
wire         io_diffCommits_commitValid_88;
wire         io_diffCommits_commitValid_89;
wire         io_diffCommits_commitValid_90;
wire         io_diffCommits_commitValid_91;
wire         io_diffCommits_commitValid_92;
wire         io_diffCommits_commitValid_93;
wire         io_diffCommits_commitValid_94;
wire         io_diffCommits_commitValid_95;
wire         io_diffCommits_commitValid_96;
wire         io_diffCommits_commitValid_97;
wire         io_diffCommits_commitValid_98;
wire         io_diffCommits_commitValid_99;
wire         io_diffCommits_commitValid_100;
wire         io_diffCommits_commitValid_101;
wire         io_diffCommits_commitValid_102;
wire         io_diffCommits_commitValid_103;
wire         io_diffCommits_commitValid_104;
wire         io_diffCommits_commitValid_105;
wire         io_diffCommits_commitValid_106;
wire         io_diffCommits_commitValid_107;
wire         io_diffCommits_commitValid_108;
wire         io_diffCommits_commitValid_109;
wire         io_diffCommits_commitValid_110;
wire         io_diffCommits_commitValid_111;
wire         io_diffCommits_commitValid_112;
wire         io_diffCommits_commitValid_113;
wire         io_diffCommits_commitValid_114;
wire         io_diffCommits_commitValid_115;
wire         io_diffCommits_commitValid_116;
wire         io_diffCommits_commitValid_117;
wire         io_diffCommits_commitValid_118;
wire         io_diffCommits_commitValid_119;
wire         io_diffCommits_commitValid_120;
wire         io_diffCommits_commitValid_121;
wire         io_diffCommits_commitValid_122;
wire         io_diffCommits_commitValid_123;
wire         io_diffCommits_commitValid_124;
wire         io_diffCommits_commitValid_125;
wire         io_diffCommits_commitValid_126;
wire         io_diffCommits_commitValid_127;
wire         io_diffCommits_commitValid_128;
wire         io_diffCommits_commitValid_129;
wire         io_diffCommits_commitValid_130;
wire         io_diffCommits_commitValid_131;
wire         io_diffCommits_commitValid_132;
wire         io_diffCommits_commitValid_133;
wire         io_diffCommits_commitValid_134;
wire         io_diffCommits_commitValid_135;
wire         io_diffCommits_commitValid_136;
wire         io_diffCommits_commitValid_137;
wire         io_diffCommits_commitValid_138;
wire         io_diffCommits_commitValid_139;
wire         io_diffCommits_commitValid_140;
wire         io_diffCommits_commitValid_141;
wire         io_diffCommits_commitValid_142;
wire         io_diffCommits_commitValid_143;
wire         io_diffCommits_commitValid_144;
wire         io_diffCommits_commitValid_145;
wire         io_diffCommits_commitValid_146;
wire         io_diffCommits_commitValid_147;
wire         io_diffCommits_commitValid_148;
wire         io_diffCommits_commitValid_149;
wire         io_diffCommits_commitValid_150;
wire         io_diffCommits_commitValid_151;
wire         io_diffCommits_commitValid_152;
wire         io_diffCommits_commitValid_153;
wire         io_diffCommits_commitValid_154;
wire         io_diffCommits_commitValid_155;
wire         io_diffCommits_commitValid_156;
wire         io_diffCommits_commitValid_157;
wire         io_diffCommits_commitValid_158;
wire         io_diffCommits_commitValid_159;
wire         io_diffCommits_commitValid_160;
wire         io_diffCommits_commitValid_161;
wire         io_diffCommits_commitValid_162;
wire         io_diffCommits_commitValid_163;
wire         io_diffCommits_commitValid_164;
wire         io_diffCommits_commitValid_165;
wire         io_diffCommits_commitValid_166;
wire         io_diffCommits_commitValid_167;
wire         io_diffCommits_commitValid_168;
wire         io_diffCommits_commitValid_169;
wire         io_diffCommits_commitValid_170;
wire         io_diffCommits_commitValid_171;
wire         io_diffCommits_commitValid_172;
wire         io_diffCommits_commitValid_173;
wire         io_diffCommits_commitValid_174;
wire         io_diffCommits_commitValid_175;
wire         io_diffCommits_commitValid_176;
wire         io_diffCommits_commitValid_177;
wire         io_diffCommits_commitValid_178;
wire         io_diffCommits_commitValid_179;
wire         io_diffCommits_commitValid_180;
wire         io_diffCommits_commitValid_181;
wire         io_diffCommits_commitValid_182;
wire         io_diffCommits_commitValid_183;
wire         io_diffCommits_commitValid_184;
wire         io_diffCommits_commitValid_185;
wire         io_diffCommits_commitValid_186;
wire         io_diffCommits_commitValid_187;
wire         io_diffCommits_commitValid_188;
wire         io_diffCommits_commitValid_189;
wire         io_diffCommits_commitValid_190;
wire         io_diffCommits_commitValid_191;
wire         io_diffCommits_commitValid_192;
wire         io_diffCommits_commitValid_193;
wire         io_diffCommits_commitValid_194;
wire         io_diffCommits_commitValid_195;
wire         io_diffCommits_commitValid_196;
wire         io_diffCommits_commitValid_197;
wire         io_diffCommits_commitValid_198;
wire         io_diffCommits_commitValid_199;
wire         io_diffCommits_commitValid_200;
wire         io_diffCommits_commitValid_201;
wire         io_diffCommits_commitValid_202;
wire         io_diffCommits_commitValid_203;
wire         io_diffCommits_commitValid_204;
wire         io_diffCommits_commitValid_205;
wire         io_diffCommits_commitValid_206;
wire         io_diffCommits_commitValid_207;
wire         io_diffCommits_commitValid_208;
wire         io_diffCommits_commitValid_209;
wire         io_diffCommits_commitValid_210;
wire         io_diffCommits_commitValid_211;
wire         io_diffCommits_commitValid_212;
wire         io_diffCommits_commitValid_213;
wire         io_diffCommits_commitValid_214;
wire         io_diffCommits_commitValid_215;
wire         io_diffCommits_commitValid_216;
wire         io_diffCommits_commitValid_217;
wire         io_diffCommits_commitValid_218;
wire         io_diffCommits_commitValid_219;
wire         io_diffCommits_commitValid_220;
wire         io_diffCommits_commitValid_221;
wire         io_diffCommits_commitValid_222;
wire         io_diffCommits_commitValid_223;
wire         io_diffCommits_commitValid_224;
wire         io_diffCommits_commitValid_225;
wire         io_diffCommits_commitValid_226;
wire         io_diffCommits_commitValid_227;
wire         io_diffCommits_commitValid_228;
wire         io_diffCommits_commitValid_229;
wire         io_diffCommits_commitValid_230;
wire         io_diffCommits_commitValid_231;
wire         io_diffCommits_commitValid_232;
wire         io_diffCommits_commitValid_233;
wire         io_diffCommits_commitValid_234;
wire         io_diffCommits_commitValid_235;
wire         io_diffCommits_commitValid_236;
wire         io_diffCommits_commitValid_237;
wire         io_diffCommits_commitValid_238;
wire         io_diffCommits_commitValid_239;
wire         io_diffCommits_commitValid_240;
wire         io_diffCommits_commitValid_241;
wire         io_diffCommits_commitValid_242;
wire         io_diffCommits_commitValid_243;
wire         io_diffCommits_commitValid_244;
wire         io_diffCommits_commitValid_245;
wire         io_diffCommits_commitValid_246;
wire         io_diffCommits_commitValid_247;
wire         io_diffCommits_commitValid_248;
wire         io_diffCommits_commitValid_249;
wire         io_diffCommits_commitValid_250;
wire         io_diffCommits_commitValid_251;
wire         io_diffCommits_commitValid_252;
wire         io_diffCommits_commitValid_253;
wire         io_diffCommits_commitValid_254;
wire [5:0]   io_diffCommits_info_0_ldest;
wire [7:0]   io_diffCommits_info_0_pdest;
wire         io_diffCommits_info_0_rfWen;
wire         io_diffCommits_info_0_fpWen;
wire         io_diffCommits_info_0_vecWen;
wire         io_diffCommits_info_0_v0Wen;
wire         io_diffCommits_info_0_vlWen;
wire [5:0]   io_diffCommits_info_1_ldest;
wire [7:0]   io_diffCommits_info_1_pdest;
wire         io_diffCommits_info_1_rfWen;
wire         io_diffCommits_info_1_fpWen;
wire         io_diffCommits_info_1_vecWen;
wire         io_diffCommits_info_1_v0Wen;
wire         io_diffCommits_info_1_vlWen;
wire [5:0]   io_diffCommits_info_2_ldest;
wire [7:0]   io_diffCommits_info_2_pdest;
wire         io_diffCommits_info_2_rfWen;
wire         io_diffCommits_info_2_fpWen;
wire         io_diffCommits_info_2_vecWen;
wire         io_diffCommits_info_2_v0Wen;
wire         io_diffCommits_info_2_vlWen;
wire [5:0]   io_diffCommits_info_3_ldest;
wire [7:0]   io_diffCommits_info_3_pdest;
wire         io_diffCommits_info_3_rfWen;
wire         io_diffCommits_info_3_fpWen;
wire         io_diffCommits_info_3_vecWen;
wire         io_diffCommits_info_3_v0Wen;
wire         io_diffCommits_info_3_vlWen;
wire [5:0]   io_diffCommits_info_4_ldest;
wire [7:0]   io_diffCommits_info_4_pdest;
wire         io_diffCommits_info_4_rfWen;
wire         io_diffCommits_info_4_fpWen;
wire         io_diffCommits_info_4_vecWen;
wire         io_diffCommits_info_4_v0Wen;
wire         io_diffCommits_info_4_vlWen;
wire [5:0]   io_diffCommits_info_5_ldest;
wire [7:0]   io_diffCommits_info_5_pdest;
wire         io_diffCommits_info_5_rfWen;
wire         io_diffCommits_info_5_fpWen;
wire         io_diffCommits_info_5_vecWen;
wire         io_diffCommits_info_5_v0Wen;
wire         io_diffCommits_info_5_vlWen;
wire [5:0]   io_diffCommits_info_6_ldest;
wire [7:0]   io_diffCommits_info_6_pdest;
wire         io_diffCommits_info_6_rfWen;
wire         io_diffCommits_info_6_fpWen;
wire         io_diffCommits_info_6_vecWen;
wire         io_diffCommits_info_6_v0Wen;
wire         io_diffCommits_info_6_vlWen;
wire [5:0]   io_diffCommits_info_7_ldest;
wire [7:0]   io_diffCommits_info_7_pdest;
wire         io_diffCommits_info_7_rfWen;
wire         io_diffCommits_info_7_fpWen;
wire         io_diffCommits_info_7_vecWen;
wire         io_diffCommits_info_7_v0Wen;
wire         io_diffCommits_info_7_vlWen;
wire [5:0]   io_diffCommits_info_8_ldest;
wire [7:0]   io_diffCommits_info_8_pdest;
wire         io_diffCommits_info_8_rfWen;
wire         io_diffCommits_info_8_fpWen;
wire         io_diffCommits_info_8_vecWen;
wire         io_diffCommits_info_8_v0Wen;
wire         io_diffCommits_info_8_vlWen;
wire [5:0]   io_diffCommits_info_9_ldest;
wire [7:0]   io_diffCommits_info_9_pdest;
wire         io_diffCommits_info_9_rfWen;
wire         io_diffCommits_info_9_fpWen;
wire         io_diffCommits_info_9_vecWen;
wire         io_diffCommits_info_9_v0Wen;
wire         io_diffCommits_info_9_vlWen;
wire [5:0]   io_diffCommits_info_10_ldest;
wire [7:0]   io_diffCommits_info_10_pdest;
wire         io_diffCommits_info_10_rfWen;
wire         io_diffCommits_info_10_fpWen;
wire         io_diffCommits_info_10_vecWen;
wire         io_diffCommits_info_10_v0Wen;
wire         io_diffCommits_info_10_vlWen;
wire [5:0]   io_diffCommits_info_11_ldest;
wire [7:0]   io_diffCommits_info_11_pdest;
wire         io_diffCommits_info_11_rfWen;
wire         io_diffCommits_info_11_fpWen;
wire         io_diffCommits_info_11_vecWen;
wire         io_diffCommits_info_11_v0Wen;
wire         io_diffCommits_info_11_vlWen;
wire [5:0]   io_diffCommits_info_12_ldest;
wire [7:0]   io_diffCommits_info_12_pdest;
wire         io_diffCommits_info_12_rfWen;
wire         io_diffCommits_info_12_fpWen;
wire         io_diffCommits_info_12_vecWen;
wire         io_diffCommits_info_12_v0Wen;
wire         io_diffCommits_info_12_vlWen;
wire [5:0]   io_diffCommits_info_13_ldest;
wire [7:0]   io_diffCommits_info_13_pdest;
wire         io_diffCommits_info_13_rfWen;
wire         io_diffCommits_info_13_fpWen;
wire         io_diffCommits_info_13_vecWen;
wire         io_diffCommits_info_13_v0Wen;
wire         io_diffCommits_info_13_vlWen;
wire [5:0]   io_diffCommits_info_14_ldest;
wire [7:0]   io_diffCommits_info_14_pdest;
wire         io_diffCommits_info_14_rfWen;
wire         io_diffCommits_info_14_fpWen;
wire         io_diffCommits_info_14_vecWen;
wire         io_diffCommits_info_14_v0Wen;
wire         io_diffCommits_info_14_vlWen;
wire [5:0]   io_diffCommits_info_15_ldest;
wire [7:0]   io_diffCommits_info_15_pdest;
wire         io_diffCommits_info_15_rfWen;
wire         io_diffCommits_info_15_fpWen;
wire         io_diffCommits_info_15_vecWen;
wire         io_diffCommits_info_15_v0Wen;
wire         io_diffCommits_info_15_vlWen;
wire [5:0]   io_diffCommits_info_16_ldest;
wire [7:0]   io_diffCommits_info_16_pdest;
wire         io_diffCommits_info_16_rfWen;
wire         io_diffCommits_info_16_fpWen;
wire         io_diffCommits_info_16_vecWen;
wire         io_diffCommits_info_16_v0Wen;
wire         io_diffCommits_info_16_vlWen;
wire [5:0]   io_diffCommits_info_17_ldest;
wire [7:0]   io_diffCommits_info_17_pdest;
wire         io_diffCommits_info_17_rfWen;
wire         io_diffCommits_info_17_fpWen;
wire         io_diffCommits_info_17_vecWen;
wire         io_diffCommits_info_17_v0Wen;
wire         io_diffCommits_info_17_vlWen;
wire [5:0]   io_diffCommits_info_18_ldest;
wire [7:0]   io_diffCommits_info_18_pdest;
wire         io_diffCommits_info_18_rfWen;
wire         io_diffCommits_info_18_fpWen;
wire         io_diffCommits_info_18_vecWen;
wire         io_diffCommits_info_18_v0Wen;
wire         io_diffCommits_info_18_vlWen;
wire [5:0]   io_diffCommits_info_19_ldest;
wire [7:0]   io_diffCommits_info_19_pdest;
wire         io_diffCommits_info_19_rfWen;
wire         io_diffCommits_info_19_fpWen;
wire         io_diffCommits_info_19_vecWen;
wire         io_diffCommits_info_19_v0Wen;
wire         io_diffCommits_info_19_vlWen;
wire [5:0]   io_diffCommits_info_20_ldest;
wire [7:0]   io_diffCommits_info_20_pdest;
wire         io_diffCommits_info_20_rfWen;
wire         io_diffCommits_info_20_fpWen;
wire         io_diffCommits_info_20_vecWen;
wire         io_diffCommits_info_20_v0Wen;
wire         io_diffCommits_info_20_vlWen;
wire [5:0]   io_diffCommits_info_21_ldest;
wire [7:0]   io_diffCommits_info_21_pdest;
wire         io_diffCommits_info_21_rfWen;
wire         io_diffCommits_info_21_fpWen;
wire         io_diffCommits_info_21_vecWen;
wire         io_diffCommits_info_21_v0Wen;
wire         io_diffCommits_info_21_vlWen;
wire [5:0]   io_diffCommits_info_22_ldest;
wire [7:0]   io_diffCommits_info_22_pdest;
wire         io_diffCommits_info_22_rfWen;
wire         io_diffCommits_info_22_fpWen;
wire         io_diffCommits_info_22_vecWen;
wire         io_diffCommits_info_22_v0Wen;
wire         io_diffCommits_info_22_vlWen;
wire [5:0]   io_diffCommits_info_23_ldest;
wire [7:0]   io_diffCommits_info_23_pdest;
wire         io_diffCommits_info_23_rfWen;
wire         io_diffCommits_info_23_fpWen;
wire         io_diffCommits_info_23_vecWen;
wire         io_diffCommits_info_23_v0Wen;
wire         io_diffCommits_info_23_vlWen;
wire [5:0]   io_diffCommits_info_24_ldest;
wire [7:0]   io_diffCommits_info_24_pdest;
wire         io_diffCommits_info_24_rfWen;
wire         io_diffCommits_info_24_fpWen;
wire         io_diffCommits_info_24_vecWen;
wire         io_diffCommits_info_24_v0Wen;
wire         io_diffCommits_info_24_vlWen;
wire [5:0]   io_diffCommits_info_25_ldest;
wire [7:0]   io_diffCommits_info_25_pdest;
wire         io_diffCommits_info_25_rfWen;
wire         io_diffCommits_info_25_fpWen;
wire         io_diffCommits_info_25_vecWen;
wire         io_diffCommits_info_25_v0Wen;
wire         io_diffCommits_info_25_vlWen;
wire [5:0]   io_diffCommits_info_26_ldest;
wire [7:0]   io_diffCommits_info_26_pdest;
wire         io_diffCommits_info_26_rfWen;
wire         io_diffCommits_info_26_fpWen;
wire         io_diffCommits_info_26_vecWen;
wire         io_diffCommits_info_26_v0Wen;
wire         io_diffCommits_info_26_vlWen;
wire [5:0]   io_diffCommits_info_27_ldest;
wire [7:0]   io_diffCommits_info_27_pdest;
wire         io_diffCommits_info_27_rfWen;
wire         io_diffCommits_info_27_fpWen;
wire         io_diffCommits_info_27_vecWen;
wire         io_diffCommits_info_27_v0Wen;
wire         io_diffCommits_info_27_vlWen;
wire [5:0]   io_diffCommits_info_28_ldest;
wire [7:0]   io_diffCommits_info_28_pdest;
wire         io_diffCommits_info_28_rfWen;
wire         io_diffCommits_info_28_fpWen;
wire         io_diffCommits_info_28_vecWen;
wire         io_diffCommits_info_28_v0Wen;
wire         io_diffCommits_info_28_vlWen;
wire [5:0]   io_diffCommits_info_29_ldest;
wire [7:0]   io_diffCommits_info_29_pdest;
wire         io_diffCommits_info_29_rfWen;
wire         io_diffCommits_info_29_fpWen;
wire         io_diffCommits_info_29_vecWen;
wire         io_diffCommits_info_29_v0Wen;
wire         io_diffCommits_info_29_vlWen;
wire [5:0]   io_diffCommits_info_30_ldest;
wire [7:0]   io_diffCommits_info_30_pdest;
wire         io_diffCommits_info_30_rfWen;
wire         io_diffCommits_info_30_fpWen;
wire         io_diffCommits_info_30_vecWen;
wire         io_diffCommits_info_30_v0Wen;
wire         io_diffCommits_info_30_vlWen;
wire [5:0]   io_diffCommits_info_31_ldest;
wire [7:0]   io_diffCommits_info_31_pdest;
wire         io_diffCommits_info_31_rfWen;
wire         io_diffCommits_info_31_fpWen;
wire         io_diffCommits_info_31_vecWen;
wire         io_diffCommits_info_31_v0Wen;
wire         io_diffCommits_info_31_vlWen;
wire [5:0]   io_diffCommits_info_32_ldest;
wire [7:0]   io_diffCommits_info_32_pdest;
wire         io_diffCommits_info_32_rfWen;
wire         io_diffCommits_info_32_fpWen;
wire         io_diffCommits_info_32_vecWen;
wire         io_diffCommits_info_32_v0Wen;
wire         io_diffCommits_info_32_vlWen;
wire [5:0]   io_diffCommits_info_33_ldest;
wire [7:0]   io_diffCommits_info_33_pdest;
wire         io_diffCommits_info_33_rfWen;
wire         io_diffCommits_info_33_fpWen;
wire         io_diffCommits_info_33_vecWen;
wire         io_diffCommits_info_33_v0Wen;
wire         io_diffCommits_info_33_vlWen;
wire [5:0]   io_diffCommits_info_34_ldest;
wire [7:0]   io_diffCommits_info_34_pdest;
wire         io_diffCommits_info_34_rfWen;
wire         io_diffCommits_info_34_fpWen;
wire         io_diffCommits_info_34_vecWen;
wire         io_diffCommits_info_34_v0Wen;
wire         io_diffCommits_info_34_vlWen;
wire [5:0]   io_diffCommits_info_35_ldest;
wire [7:0]   io_diffCommits_info_35_pdest;
wire         io_diffCommits_info_35_rfWen;
wire         io_diffCommits_info_35_fpWen;
wire         io_diffCommits_info_35_vecWen;
wire         io_diffCommits_info_35_v0Wen;
wire         io_diffCommits_info_35_vlWen;
wire [5:0]   io_diffCommits_info_36_ldest;
wire [7:0]   io_diffCommits_info_36_pdest;
wire         io_diffCommits_info_36_rfWen;
wire         io_diffCommits_info_36_fpWen;
wire         io_diffCommits_info_36_vecWen;
wire         io_diffCommits_info_36_v0Wen;
wire         io_diffCommits_info_36_vlWen;
wire [5:0]   io_diffCommits_info_37_ldest;
wire [7:0]   io_diffCommits_info_37_pdest;
wire         io_diffCommits_info_37_rfWen;
wire         io_diffCommits_info_37_fpWen;
wire         io_diffCommits_info_37_vecWen;
wire         io_diffCommits_info_37_v0Wen;
wire         io_diffCommits_info_37_vlWen;
wire [5:0]   io_diffCommits_info_38_ldest;
wire [7:0]   io_diffCommits_info_38_pdest;
wire         io_diffCommits_info_38_rfWen;
wire         io_diffCommits_info_38_fpWen;
wire         io_diffCommits_info_38_vecWen;
wire         io_diffCommits_info_38_v0Wen;
wire         io_diffCommits_info_38_vlWen;
wire [5:0]   io_diffCommits_info_39_ldest;
wire [7:0]   io_diffCommits_info_39_pdest;
wire         io_diffCommits_info_39_rfWen;
wire         io_diffCommits_info_39_fpWen;
wire         io_diffCommits_info_39_vecWen;
wire         io_diffCommits_info_39_v0Wen;
wire         io_diffCommits_info_39_vlWen;
wire [5:0]   io_diffCommits_info_40_ldest;
wire [7:0]   io_diffCommits_info_40_pdest;
wire         io_diffCommits_info_40_rfWen;
wire         io_diffCommits_info_40_fpWen;
wire         io_diffCommits_info_40_vecWen;
wire         io_diffCommits_info_40_v0Wen;
wire         io_diffCommits_info_40_vlWen;
wire [5:0]   io_diffCommits_info_41_ldest;
wire [7:0]   io_diffCommits_info_41_pdest;
wire         io_diffCommits_info_41_rfWen;
wire         io_diffCommits_info_41_fpWen;
wire         io_diffCommits_info_41_vecWen;
wire         io_diffCommits_info_41_v0Wen;
wire         io_diffCommits_info_41_vlWen;
wire [5:0]   io_diffCommits_info_42_ldest;
wire [7:0]   io_diffCommits_info_42_pdest;
wire         io_diffCommits_info_42_rfWen;
wire         io_diffCommits_info_42_fpWen;
wire         io_diffCommits_info_42_vecWen;
wire         io_diffCommits_info_42_v0Wen;
wire         io_diffCommits_info_42_vlWen;
wire [5:0]   io_diffCommits_info_43_ldest;
wire [7:0]   io_diffCommits_info_43_pdest;
wire         io_diffCommits_info_43_rfWen;
wire         io_diffCommits_info_43_fpWen;
wire         io_diffCommits_info_43_vecWen;
wire         io_diffCommits_info_43_v0Wen;
wire         io_diffCommits_info_43_vlWen;
wire [5:0]   io_diffCommits_info_44_ldest;
wire [7:0]   io_diffCommits_info_44_pdest;
wire         io_diffCommits_info_44_rfWen;
wire         io_diffCommits_info_44_fpWen;
wire         io_diffCommits_info_44_vecWen;
wire         io_diffCommits_info_44_v0Wen;
wire         io_diffCommits_info_44_vlWen;
wire [5:0]   io_diffCommits_info_45_ldest;
wire [7:0]   io_diffCommits_info_45_pdest;
wire         io_diffCommits_info_45_rfWen;
wire         io_diffCommits_info_45_fpWen;
wire         io_diffCommits_info_45_vecWen;
wire         io_diffCommits_info_45_v0Wen;
wire         io_diffCommits_info_45_vlWen;
wire [5:0]   io_diffCommits_info_46_ldest;
wire [7:0]   io_diffCommits_info_46_pdest;
wire         io_diffCommits_info_46_rfWen;
wire         io_diffCommits_info_46_fpWen;
wire         io_diffCommits_info_46_vecWen;
wire         io_diffCommits_info_46_v0Wen;
wire         io_diffCommits_info_46_vlWen;
wire [5:0]   io_diffCommits_info_47_ldest;
wire [7:0]   io_diffCommits_info_47_pdest;
wire         io_diffCommits_info_47_rfWen;
wire         io_diffCommits_info_47_fpWen;
wire         io_diffCommits_info_47_vecWen;
wire         io_diffCommits_info_47_v0Wen;
wire         io_diffCommits_info_47_vlWen;
wire [5:0]   io_diffCommits_info_48_ldest;
wire [7:0]   io_diffCommits_info_48_pdest;
wire         io_diffCommits_info_48_rfWen;
wire         io_diffCommits_info_48_fpWen;
wire         io_diffCommits_info_48_vecWen;
wire         io_diffCommits_info_48_v0Wen;
wire         io_diffCommits_info_48_vlWen;
wire [5:0]   io_diffCommits_info_49_ldest;
wire [7:0]   io_diffCommits_info_49_pdest;
wire         io_diffCommits_info_49_rfWen;
wire         io_diffCommits_info_49_fpWen;
wire         io_diffCommits_info_49_vecWen;
wire         io_diffCommits_info_49_v0Wen;
wire         io_diffCommits_info_49_vlWen;
wire [5:0]   io_diffCommits_info_50_ldest;
wire [7:0]   io_diffCommits_info_50_pdest;
wire         io_diffCommits_info_50_rfWen;
wire         io_diffCommits_info_50_fpWen;
wire         io_diffCommits_info_50_vecWen;
wire         io_diffCommits_info_50_v0Wen;
wire         io_diffCommits_info_50_vlWen;
wire [5:0]   io_diffCommits_info_51_ldest;
wire [7:0]   io_diffCommits_info_51_pdest;
wire         io_diffCommits_info_51_rfWen;
wire         io_diffCommits_info_51_fpWen;
wire         io_diffCommits_info_51_vecWen;
wire         io_diffCommits_info_51_v0Wen;
wire         io_diffCommits_info_51_vlWen;
wire [5:0]   io_diffCommits_info_52_ldest;
wire [7:0]   io_diffCommits_info_52_pdest;
wire         io_diffCommits_info_52_rfWen;
wire         io_diffCommits_info_52_fpWen;
wire         io_diffCommits_info_52_vecWen;
wire         io_diffCommits_info_52_v0Wen;
wire         io_diffCommits_info_52_vlWen;
wire [5:0]   io_diffCommits_info_53_ldest;
wire [7:0]   io_diffCommits_info_53_pdest;
wire         io_diffCommits_info_53_rfWen;
wire         io_diffCommits_info_53_fpWen;
wire         io_diffCommits_info_53_vecWen;
wire         io_diffCommits_info_53_v0Wen;
wire         io_diffCommits_info_53_vlWen;
wire [5:0]   io_diffCommits_info_54_ldest;
wire [7:0]   io_diffCommits_info_54_pdest;
wire         io_diffCommits_info_54_rfWen;
wire         io_diffCommits_info_54_fpWen;
wire         io_diffCommits_info_54_vecWen;
wire         io_diffCommits_info_54_v0Wen;
wire         io_diffCommits_info_54_vlWen;
wire [5:0]   io_diffCommits_info_55_ldest;
wire [7:0]   io_diffCommits_info_55_pdest;
wire         io_diffCommits_info_55_rfWen;
wire         io_diffCommits_info_55_fpWen;
wire         io_diffCommits_info_55_vecWen;
wire         io_diffCommits_info_55_v0Wen;
wire         io_diffCommits_info_55_vlWen;
wire [5:0]   io_diffCommits_info_56_ldest;
wire [7:0]   io_diffCommits_info_56_pdest;
wire         io_diffCommits_info_56_rfWen;
wire         io_diffCommits_info_56_fpWen;
wire         io_diffCommits_info_56_vecWen;
wire         io_diffCommits_info_56_v0Wen;
wire         io_diffCommits_info_56_vlWen;
wire [5:0]   io_diffCommits_info_57_ldest;
wire [7:0]   io_diffCommits_info_57_pdest;
wire         io_diffCommits_info_57_rfWen;
wire         io_diffCommits_info_57_fpWen;
wire         io_diffCommits_info_57_vecWen;
wire         io_diffCommits_info_57_v0Wen;
wire         io_diffCommits_info_57_vlWen;
wire [5:0]   io_diffCommits_info_58_ldest;
wire [7:0]   io_diffCommits_info_58_pdest;
wire         io_diffCommits_info_58_rfWen;
wire         io_diffCommits_info_58_fpWen;
wire         io_diffCommits_info_58_vecWen;
wire         io_diffCommits_info_58_v0Wen;
wire         io_diffCommits_info_58_vlWen;
wire [5:0]   io_diffCommits_info_59_ldest;
wire [7:0]   io_diffCommits_info_59_pdest;
wire         io_diffCommits_info_59_rfWen;
wire         io_diffCommits_info_59_fpWen;
wire         io_diffCommits_info_59_vecWen;
wire         io_diffCommits_info_59_v0Wen;
wire         io_diffCommits_info_59_vlWen;
wire [5:0]   io_diffCommits_info_60_ldest;
wire [7:0]   io_diffCommits_info_60_pdest;
wire         io_diffCommits_info_60_rfWen;
wire         io_diffCommits_info_60_fpWen;
wire         io_diffCommits_info_60_vecWen;
wire         io_diffCommits_info_60_v0Wen;
wire         io_diffCommits_info_60_vlWen;
wire [5:0]   io_diffCommits_info_61_ldest;
wire [7:0]   io_diffCommits_info_61_pdest;
wire         io_diffCommits_info_61_rfWen;
wire         io_diffCommits_info_61_fpWen;
wire         io_diffCommits_info_61_vecWen;
wire         io_diffCommits_info_61_v0Wen;
wire         io_diffCommits_info_61_vlWen;
wire [5:0]   io_diffCommits_info_62_ldest;
wire [7:0]   io_diffCommits_info_62_pdest;
wire         io_diffCommits_info_62_rfWen;
wire         io_diffCommits_info_62_fpWen;
wire         io_diffCommits_info_62_vecWen;
wire         io_diffCommits_info_62_v0Wen;
wire         io_diffCommits_info_62_vlWen;
wire [5:0]   io_diffCommits_info_63_ldest;
wire [7:0]   io_diffCommits_info_63_pdest;
wire         io_diffCommits_info_63_rfWen;
wire         io_diffCommits_info_63_fpWen;
wire         io_diffCommits_info_63_vecWen;
wire         io_diffCommits_info_63_v0Wen;
wire         io_diffCommits_info_63_vlWen;
wire [5:0]   io_diffCommits_info_64_ldest;
wire [7:0]   io_diffCommits_info_64_pdest;
wire         io_diffCommits_info_64_rfWen;
wire         io_diffCommits_info_64_fpWen;
wire         io_diffCommits_info_64_vecWen;
wire         io_diffCommits_info_64_v0Wen;
wire         io_diffCommits_info_64_vlWen;
wire [5:0]   io_diffCommits_info_65_ldest;
wire [7:0]   io_diffCommits_info_65_pdest;
wire         io_diffCommits_info_65_rfWen;
wire         io_diffCommits_info_65_fpWen;
wire         io_diffCommits_info_65_vecWen;
wire         io_diffCommits_info_65_v0Wen;
wire         io_diffCommits_info_65_vlWen;
wire [5:0]   io_diffCommits_info_66_ldest;
wire [7:0]   io_diffCommits_info_66_pdest;
wire         io_diffCommits_info_66_rfWen;
wire         io_diffCommits_info_66_fpWen;
wire         io_diffCommits_info_66_vecWen;
wire         io_diffCommits_info_66_v0Wen;
wire         io_diffCommits_info_66_vlWen;
wire [5:0]   io_diffCommits_info_67_ldest;
wire [7:0]   io_diffCommits_info_67_pdest;
wire         io_diffCommits_info_67_rfWen;
wire         io_diffCommits_info_67_fpWen;
wire         io_diffCommits_info_67_vecWen;
wire         io_diffCommits_info_67_v0Wen;
wire         io_diffCommits_info_67_vlWen;
wire [5:0]   io_diffCommits_info_68_ldest;
wire [7:0]   io_diffCommits_info_68_pdest;
wire         io_diffCommits_info_68_rfWen;
wire         io_diffCommits_info_68_fpWen;
wire         io_diffCommits_info_68_vecWen;
wire         io_diffCommits_info_68_v0Wen;
wire         io_diffCommits_info_68_vlWen;
wire [5:0]   io_diffCommits_info_69_ldest;
wire [7:0]   io_diffCommits_info_69_pdest;
wire         io_diffCommits_info_69_rfWen;
wire         io_diffCommits_info_69_fpWen;
wire         io_diffCommits_info_69_vecWen;
wire         io_diffCommits_info_69_v0Wen;
wire         io_diffCommits_info_69_vlWen;
wire [5:0]   io_diffCommits_info_70_ldest;
wire [7:0]   io_diffCommits_info_70_pdest;
wire         io_diffCommits_info_70_rfWen;
wire         io_diffCommits_info_70_fpWen;
wire         io_diffCommits_info_70_vecWen;
wire         io_diffCommits_info_70_v0Wen;
wire         io_diffCommits_info_70_vlWen;
wire [5:0]   io_diffCommits_info_71_ldest;
wire [7:0]   io_diffCommits_info_71_pdest;
wire         io_diffCommits_info_71_rfWen;
wire         io_diffCommits_info_71_fpWen;
wire         io_diffCommits_info_71_vecWen;
wire         io_diffCommits_info_71_v0Wen;
wire         io_diffCommits_info_71_vlWen;
wire [5:0]   io_diffCommits_info_72_ldest;
wire [7:0]   io_diffCommits_info_72_pdest;
wire         io_diffCommits_info_72_rfWen;
wire         io_diffCommits_info_72_fpWen;
wire         io_diffCommits_info_72_vecWen;
wire         io_diffCommits_info_72_v0Wen;
wire         io_diffCommits_info_72_vlWen;
wire [5:0]   io_diffCommits_info_73_ldest;
wire [7:0]   io_diffCommits_info_73_pdest;
wire         io_diffCommits_info_73_rfWen;
wire         io_diffCommits_info_73_fpWen;
wire         io_diffCommits_info_73_vecWen;
wire         io_diffCommits_info_73_v0Wen;
wire         io_diffCommits_info_73_vlWen;
wire [5:0]   io_diffCommits_info_74_ldest;
wire [7:0]   io_diffCommits_info_74_pdest;
wire         io_diffCommits_info_74_rfWen;
wire         io_diffCommits_info_74_fpWen;
wire         io_diffCommits_info_74_vecWen;
wire         io_diffCommits_info_74_v0Wen;
wire         io_diffCommits_info_74_vlWen;
wire [5:0]   io_diffCommits_info_75_ldest;
wire [7:0]   io_diffCommits_info_75_pdest;
wire         io_diffCommits_info_75_rfWen;
wire         io_diffCommits_info_75_fpWen;
wire         io_diffCommits_info_75_vecWen;
wire         io_diffCommits_info_75_v0Wen;
wire         io_diffCommits_info_75_vlWen;
wire [5:0]   io_diffCommits_info_76_ldest;
wire [7:0]   io_diffCommits_info_76_pdest;
wire         io_diffCommits_info_76_rfWen;
wire         io_diffCommits_info_76_fpWen;
wire         io_diffCommits_info_76_vecWen;
wire         io_diffCommits_info_76_v0Wen;
wire         io_diffCommits_info_76_vlWen;
wire [5:0]   io_diffCommits_info_77_ldest;
wire [7:0]   io_diffCommits_info_77_pdest;
wire         io_diffCommits_info_77_rfWen;
wire         io_diffCommits_info_77_fpWen;
wire         io_diffCommits_info_77_vecWen;
wire         io_diffCommits_info_77_v0Wen;
wire         io_diffCommits_info_77_vlWen;
wire [5:0]   io_diffCommits_info_78_ldest;
wire [7:0]   io_diffCommits_info_78_pdest;
wire         io_diffCommits_info_78_rfWen;
wire         io_diffCommits_info_78_fpWen;
wire         io_diffCommits_info_78_vecWen;
wire         io_diffCommits_info_78_v0Wen;
wire         io_diffCommits_info_78_vlWen;
wire [5:0]   io_diffCommits_info_79_ldest;
wire [7:0]   io_diffCommits_info_79_pdest;
wire         io_diffCommits_info_79_rfWen;
wire         io_diffCommits_info_79_fpWen;
wire         io_diffCommits_info_79_vecWen;
wire         io_diffCommits_info_79_v0Wen;
wire         io_diffCommits_info_79_vlWen;
wire [5:0]   io_diffCommits_info_80_ldest;
wire [7:0]   io_diffCommits_info_80_pdest;
wire         io_diffCommits_info_80_rfWen;
wire         io_diffCommits_info_80_fpWen;
wire         io_diffCommits_info_80_vecWen;
wire         io_diffCommits_info_80_v0Wen;
wire         io_diffCommits_info_80_vlWen;
wire [5:0]   io_diffCommits_info_81_ldest;
wire [7:0]   io_diffCommits_info_81_pdest;
wire         io_diffCommits_info_81_rfWen;
wire         io_diffCommits_info_81_fpWen;
wire         io_diffCommits_info_81_vecWen;
wire         io_diffCommits_info_81_v0Wen;
wire         io_diffCommits_info_81_vlWen;
wire [5:0]   io_diffCommits_info_82_ldest;
wire [7:0]   io_diffCommits_info_82_pdest;
wire         io_diffCommits_info_82_rfWen;
wire         io_diffCommits_info_82_fpWen;
wire         io_diffCommits_info_82_vecWen;
wire         io_diffCommits_info_82_v0Wen;
wire         io_diffCommits_info_82_vlWen;
wire [5:0]   io_diffCommits_info_83_ldest;
wire [7:0]   io_diffCommits_info_83_pdest;
wire         io_diffCommits_info_83_rfWen;
wire         io_diffCommits_info_83_fpWen;
wire         io_diffCommits_info_83_vecWen;
wire         io_diffCommits_info_83_v0Wen;
wire         io_diffCommits_info_83_vlWen;
wire [5:0]   io_diffCommits_info_84_ldest;
wire [7:0]   io_diffCommits_info_84_pdest;
wire         io_diffCommits_info_84_rfWen;
wire         io_diffCommits_info_84_fpWen;
wire         io_diffCommits_info_84_vecWen;
wire         io_diffCommits_info_84_v0Wen;
wire         io_diffCommits_info_84_vlWen;
wire [5:0]   io_diffCommits_info_85_ldest;
wire [7:0]   io_diffCommits_info_85_pdest;
wire         io_diffCommits_info_85_rfWen;
wire         io_diffCommits_info_85_fpWen;
wire         io_diffCommits_info_85_vecWen;
wire         io_diffCommits_info_85_v0Wen;
wire         io_diffCommits_info_85_vlWen;
wire [5:0]   io_diffCommits_info_86_ldest;
wire [7:0]   io_diffCommits_info_86_pdest;
wire         io_diffCommits_info_86_rfWen;
wire         io_diffCommits_info_86_fpWen;
wire         io_diffCommits_info_86_vecWen;
wire         io_diffCommits_info_86_v0Wen;
wire         io_diffCommits_info_86_vlWen;
wire [5:0]   io_diffCommits_info_87_ldest;
wire [7:0]   io_diffCommits_info_87_pdest;
wire         io_diffCommits_info_87_rfWen;
wire         io_diffCommits_info_87_fpWen;
wire         io_diffCommits_info_87_vecWen;
wire         io_diffCommits_info_87_v0Wen;
wire         io_diffCommits_info_87_vlWen;
wire [5:0]   io_diffCommits_info_88_ldest;
wire [7:0]   io_diffCommits_info_88_pdest;
wire         io_diffCommits_info_88_rfWen;
wire         io_diffCommits_info_88_fpWen;
wire         io_diffCommits_info_88_vecWen;
wire         io_diffCommits_info_88_v0Wen;
wire         io_diffCommits_info_88_vlWen;
wire [5:0]   io_diffCommits_info_89_ldest;
wire [7:0]   io_diffCommits_info_89_pdest;
wire         io_diffCommits_info_89_rfWen;
wire         io_diffCommits_info_89_fpWen;
wire         io_diffCommits_info_89_vecWen;
wire         io_diffCommits_info_89_v0Wen;
wire         io_diffCommits_info_89_vlWen;
wire [5:0]   io_diffCommits_info_90_ldest;
wire [7:0]   io_diffCommits_info_90_pdest;
wire         io_diffCommits_info_90_rfWen;
wire         io_diffCommits_info_90_fpWen;
wire         io_diffCommits_info_90_vecWen;
wire         io_diffCommits_info_90_v0Wen;
wire         io_diffCommits_info_90_vlWen;
wire [5:0]   io_diffCommits_info_91_ldest;
wire [7:0]   io_diffCommits_info_91_pdest;
wire         io_diffCommits_info_91_rfWen;
wire         io_diffCommits_info_91_fpWen;
wire         io_diffCommits_info_91_vecWen;
wire         io_diffCommits_info_91_v0Wen;
wire         io_diffCommits_info_91_vlWen;
wire [5:0]   io_diffCommits_info_92_ldest;
wire [7:0]   io_diffCommits_info_92_pdest;
wire         io_diffCommits_info_92_rfWen;
wire         io_diffCommits_info_92_fpWen;
wire         io_diffCommits_info_92_vecWen;
wire         io_diffCommits_info_92_v0Wen;
wire         io_diffCommits_info_92_vlWen;
wire [5:0]   io_diffCommits_info_93_ldest;
wire [7:0]   io_diffCommits_info_93_pdest;
wire         io_diffCommits_info_93_rfWen;
wire         io_diffCommits_info_93_fpWen;
wire         io_diffCommits_info_93_vecWen;
wire         io_diffCommits_info_93_v0Wen;
wire         io_diffCommits_info_93_vlWen;
wire [5:0]   io_diffCommits_info_94_ldest;
wire [7:0]   io_diffCommits_info_94_pdest;
wire         io_diffCommits_info_94_rfWen;
wire         io_diffCommits_info_94_fpWen;
wire         io_diffCommits_info_94_vecWen;
wire         io_diffCommits_info_94_v0Wen;
wire         io_diffCommits_info_94_vlWen;
wire [5:0]   io_diffCommits_info_95_ldest;
wire [7:0]   io_diffCommits_info_95_pdest;
wire         io_diffCommits_info_95_rfWen;
wire         io_diffCommits_info_95_fpWen;
wire         io_diffCommits_info_95_vecWen;
wire         io_diffCommits_info_95_v0Wen;
wire         io_diffCommits_info_95_vlWen;
wire [5:0]   io_diffCommits_info_96_ldest;
wire [7:0]   io_diffCommits_info_96_pdest;
wire         io_diffCommits_info_96_rfWen;
wire         io_diffCommits_info_96_fpWen;
wire         io_diffCommits_info_96_vecWen;
wire         io_diffCommits_info_96_v0Wen;
wire         io_diffCommits_info_96_vlWen;
wire [5:0]   io_diffCommits_info_97_ldest;
wire [7:0]   io_diffCommits_info_97_pdest;
wire         io_diffCommits_info_97_rfWen;
wire         io_diffCommits_info_97_fpWen;
wire         io_diffCommits_info_97_vecWen;
wire         io_diffCommits_info_97_v0Wen;
wire         io_diffCommits_info_97_vlWen;
wire [5:0]   io_diffCommits_info_98_ldest;
wire [7:0]   io_diffCommits_info_98_pdest;
wire         io_diffCommits_info_98_rfWen;
wire         io_diffCommits_info_98_fpWen;
wire         io_diffCommits_info_98_vecWen;
wire         io_diffCommits_info_98_v0Wen;
wire         io_diffCommits_info_98_vlWen;
wire [5:0]   io_diffCommits_info_99_ldest;
wire [7:0]   io_diffCommits_info_99_pdest;
wire         io_diffCommits_info_99_rfWen;
wire         io_diffCommits_info_99_fpWen;
wire         io_diffCommits_info_99_vecWen;
wire         io_diffCommits_info_99_v0Wen;
wire         io_diffCommits_info_99_vlWen;
wire [5:0]   io_diffCommits_info_100_ldest;
wire [7:0]   io_diffCommits_info_100_pdest;
wire         io_diffCommits_info_100_rfWen;
wire         io_diffCommits_info_100_fpWen;
wire         io_diffCommits_info_100_vecWen;
wire         io_diffCommits_info_100_v0Wen;
wire         io_diffCommits_info_100_vlWen;
wire [5:0]   io_diffCommits_info_101_ldest;
wire [7:0]   io_diffCommits_info_101_pdest;
wire         io_diffCommits_info_101_rfWen;
wire         io_diffCommits_info_101_fpWen;
wire         io_diffCommits_info_101_vecWen;
wire         io_diffCommits_info_101_v0Wen;
wire         io_diffCommits_info_101_vlWen;
wire [5:0]   io_diffCommits_info_102_ldest;
wire [7:0]   io_diffCommits_info_102_pdest;
wire         io_diffCommits_info_102_rfWen;
wire         io_diffCommits_info_102_fpWen;
wire         io_diffCommits_info_102_vecWen;
wire         io_diffCommits_info_102_v0Wen;
wire         io_diffCommits_info_102_vlWen;
wire [5:0]   io_diffCommits_info_103_ldest;
wire [7:0]   io_diffCommits_info_103_pdest;
wire         io_diffCommits_info_103_rfWen;
wire         io_diffCommits_info_103_fpWen;
wire         io_diffCommits_info_103_vecWen;
wire         io_diffCommits_info_103_v0Wen;
wire         io_diffCommits_info_103_vlWen;
wire [5:0]   io_diffCommits_info_104_ldest;
wire [7:0]   io_diffCommits_info_104_pdest;
wire         io_diffCommits_info_104_rfWen;
wire         io_diffCommits_info_104_fpWen;
wire         io_diffCommits_info_104_vecWen;
wire         io_diffCommits_info_104_v0Wen;
wire         io_diffCommits_info_104_vlWen;
wire [5:0]   io_diffCommits_info_105_ldest;
wire [7:0]   io_diffCommits_info_105_pdest;
wire         io_diffCommits_info_105_rfWen;
wire         io_diffCommits_info_105_fpWen;
wire         io_diffCommits_info_105_vecWen;
wire         io_diffCommits_info_105_v0Wen;
wire         io_diffCommits_info_105_vlWen;
wire [5:0]   io_diffCommits_info_106_ldest;
wire [7:0]   io_diffCommits_info_106_pdest;
wire         io_diffCommits_info_106_rfWen;
wire         io_diffCommits_info_106_fpWen;
wire         io_diffCommits_info_106_vecWen;
wire         io_diffCommits_info_106_v0Wen;
wire         io_diffCommits_info_106_vlWen;
wire [5:0]   io_diffCommits_info_107_ldest;
wire [7:0]   io_diffCommits_info_107_pdest;
wire         io_diffCommits_info_107_rfWen;
wire         io_diffCommits_info_107_fpWen;
wire         io_diffCommits_info_107_vecWen;
wire         io_diffCommits_info_107_v0Wen;
wire         io_diffCommits_info_107_vlWen;
wire [5:0]   io_diffCommits_info_108_ldest;
wire [7:0]   io_diffCommits_info_108_pdest;
wire         io_diffCommits_info_108_rfWen;
wire         io_diffCommits_info_108_fpWen;
wire         io_diffCommits_info_108_vecWen;
wire         io_diffCommits_info_108_v0Wen;
wire         io_diffCommits_info_108_vlWen;
wire [5:0]   io_diffCommits_info_109_ldest;
wire [7:0]   io_diffCommits_info_109_pdest;
wire         io_diffCommits_info_109_rfWen;
wire         io_diffCommits_info_109_fpWen;
wire         io_diffCommits_info_109_vecWen;
wire         io_diffCommits_info_109_v0Wen;
wire         io_diffCommits_info_109_vlWen;
wire [5:0]   io_diffCommits_info_110_ldest;
wire [7:0]   io_diffCommits_info_110_pdest;
wire         io_diffCommits_info_110_rfWen;
wire         io_diffCommits_info_110_fpWen;
wire         io_diffCommits_info_110_vecWen;
wire         io_diffCommits_info_110_v0Wen;
wire         io_diffCommits_info_110_vlWen;
wire [5:0]   io_diffCommits_info_111_ldest;
wire [7:0]   io_diffCommits_info_111_pdest;
wire         io_diffCommits_info_111_rfWen;
wire         io_diffCommits_info_111_fpWen;
wire         io_diffCommits_info_111_vecWen;
wire         io_diffCommits_info_111_v0Wen;
wire         io_diffCommits_info_111_vlWen;
wire [5:0]   io_diffCommits_info_112_ldest;
wire [7:0]   io_diffCommits_info_112_pdest;
wire         io_diffCommits_info_112_rfWen;
wire         io_diffCommits_info_112_fpWen;
wire         io_diffCommits_info_112_vecWen;
wire         io_diffCommits_info_112_v0Wen;
wire         io_diffCommits_info_112_vlWen;
wire [5:0]   io_diffCommits_info_113_ldest;
wire [7:0]   io_diffCommits_info_113_pdest;
wire         io_diffCommits_info_113_rfWen;
wire         io_diffCommits_info_113_fpWen;
wire         io_diffCommits_info_113_vecWen;
wire         io_diffCommits_info_113_v0Wen;
wire         io_diffCommits_info_113_vlWen;
wire [5:0]   io_diffCommits_info_114_ldest;
wire [7:0]   io_diffCommits_info_114_pdest;
wire         io_diffCommits_info_114_rfWen;
wire         io_diffCommits_info_114_fpWen;
wire         io_diffCommits_info_114_vecWen;
wire         io_diffCommits_info_114_v0Wen;
wire         io_diffCommits_info_114_vlWen;
wire [5:0]   io_diffCommits_info_115_ldest;
wire [7:0]   io_diffCommits_info_115_pdest;
wire         io_diffCommits_info_115_rfWen;
wire         io_diffCommits_info_115_fpWen;
wire         io_diffCommits_info_115_vecWen;
wire         io_diffCommits_info_115_v0Wen;
wire         io_diffCommits_info_115_vlWen;
wire [5:0]   io_diffCommits_info_116_ldest;
wire [7:0]   io_diffCommits_info_116_pdest;
wire         io_diffCommits_info_116_rfWen;
wire         io_diffCommits_info_116_fpWen;
wire         io_diffCommits_info_116_vecWen;
wire         io_diffCommits_info_116_v0Wen;
wire         io_diffCommits_info_116_vlWen;
wire [5:0]   io_diffCommits_info_117_ldest;
wire [7:0]   io_diffCommits_info_117_pdest;
wire         io_diffCommits_info_117_rfWen;
wire         io_diffCommits_info_117_fpWen;
wire         io_diffCommits_info_117_vecWen;
wire         io_diffCommits_info_117_v0Wen;
wire         io_diffCommits_info_117_vlWen;
wire [5:0]   io_diffCommits_info_118_ldest;
wire [7:0]   io_diffCommits_info_118_pdest;
wire         io_diffCommits_info_118_rfWen;
wire         io_diffCommits_info_118_fpWen;
wire         io_diffCommits_info_118_vecWen;
wire         io_diffCommits_info_118_v0Wen;
wire         io_diffCommits_info_118_vlWen;
wire [5:0]   io_diffCommits_info_119_ldest;
wire [7:0]   io_diffCommits_info_119_pdest;
wire         io_diffCommits_info_119_rfWen;
wire         io_diffCommits_info_119_fpWen;
wire         io_diffCommits_info_119_vecWen;
wire         io_diffCommits_info_119_v0Wen;
wire         io_diffCommits_info_119_vlWen;
wire [5:0]   io_diffCommits_info_120_ldest;
wire [7:0]   io_diffCommits_info_120_pdest;
wire         io_diffCommits_info_120_rfWen;
wire         io_diffCommits_info_120_fpWen;
wire         io_diffCommits_info_120_vecWen;
wire         io_diffCommits_info_120_v0Wen;
wire         io_diffCommits_info_120_vlWen;
wire [5:0]   io_diffCommits_info_121_ldest;
wire [7:0]   io_diffCommits_info_121_pdest;
wire         io_diffCommits_info_121_rfWen;
wire         io_diffCommits_info_121_fpWen;
wire         io_diffCommits_info_121_vecWen;
wire         io_diffCommits_info_121_v0Wen;
wire         io_diffCommits_info_121_vlWen;
wire [5:0]   io_diffCommits_info_122_ldest;
wire [7:0]   io_diffCommits_info_122_pdest;
wire         io_diffCommits_info_122_rfWen;
wire         io_diffCommits_info_122_fpWen;
wire         io_diffCommits_info_122_vecWen;
wire         io_diffCommits_info_122_v0Wen;
wire         io_diffCommits_info_122_vlWen;
wire [5:0]   io_diffCommits_info_123_ldest;
wire [7:0]   io_diffCommits_info_123_pdest;
wire         io_diffCommits_info_123_rfWen;
wire         io_diffCommits_info_123_fpWen;
wire         io_diffCommits_info_123_vecWen;
wire         io_diffCommits_info_123_v0Wen;
wire         io_diffCommits_info_123_vlWen;
wire [5:0]   io_diffCommits_info_124_ldest;
wire [7:0]   io_diffCommits_info_124_pdest;
wire         io_diffCommits_info_124_rfWen;
wire         io_diffCommits_info_124_fpWen;
wire         io_diffCommits_info_124_vecWen;
wire         io_diffCommits_info_124_v0Wen;
wire         io_diffCommits_info_124_vlWen;
wire [5:0]   io_diffCommits_info_125_ldest;
wire [7:0]   io_diffCommits_info_125_pdest;
wire         io_diffCommits_info_125_rfWen;
wire         io_diffCommits_info_125_fpWen;
wire         io_diffCommits_info_125_vecWen;
wire         io_diffCommits_info_125_v0Wen;
wire         io_diffCommits_info_125_vlWen;
wire [5:0]   io_diffCommits_info_126_ldest;
wire [7:0]   io_diffCommits_info_126_pdest;
wire         io_diffCommits_info_126_rfWen;
wire         io_diffCommits_info_126_fpWen;
wire         io_diffCommits_info_126_vecWen;
wire         io_diffCommits_info_126_v0Wen;
wire         io_diffCommits_info_126_vlWen;
wire [5:0]   io_diffCommits_info_127_ldest;
wire [7:0]   io_diffCommits_info_127_pdest;
wire         io_diffCommits_info_127_rfWen;
wire         io_diffCommits_info_127_fpWen;
wire         io_diffCommits_info_127_vecWen;
wire         io_diffCommits_info_127_v0Wen;
wire         io_diffCommits_info_127_vlWen;
wire [5:0]   io_diffCommits_info_128_ldest;
wire [7:0]   io_diffCommits_info_128_pdest;
wire         io_diffCommits_info_128_rfWen;
wire         io_diffCommits_info_128_fpWen;
wire         io_diffCommits_info_128_vecWen;
wire         io_diffCommits_info_128_v0Wen;
wire         io_diffCommits_info_128_vlWen;
wire [5:0]   io_diffCommits_info_129_ldest;
wire [7:0]   io_diffCommits_info_129_pdest;
wire         io_diffCommits_info_129_rfWen;
wire         io_diffCommits_info_129_fpWen;
wire         io_diffCommits_info_129_vecWen;
wire         io_diffCommits_info_129_v0Wen;
wire         io_diffCommits_info_129_vlWen;
wire [5:0]   io_diffCommits_info_130_ldest;
wire [7:0]   io_diffCommits_info_130_pdest;
wire         io_diffCommits_info_130_rfWen;
wire         io_diffCommits_info_130_fpWen;
wire         io_diffCommits_info_130_vecWen;
wire         io_diffCommits_info_130_v0Wen;
wire         io_diffCommits_info_130_vlWen;
wire [5:0]   io_diffCommits_info_131_ldest;
wire [7:0]   io_diffCommits_info_131_pdest;
wire         io_diffCommits_info_131_rfWen;
wire         io_diffCommits_info_131_fpWen;
wire         io_diffCommits_info_131_vecWen;
wire         io_diffCommits_info_131_v0Wen;
wire         io_diffCommits_info_131_vlWen;
wire [5:0]   io_diffCommits_info_132_ldest;
wire [7:0]   io_diffCommits_info_132_pdest;
wire         io_diffCommits_info_132_rfWen;
wire         io_diffCommits_info_132_fpWen;
wire         io_diffCommits_info_132_vecWen;
wire         io_diffCommits_info_132_v0Wen;
wire         io_diffCommits_info_132_vlWen;
wire [5:0]   io_diffCommits_info_133_ldest;
wire [7:0]   io_diffCommits_info_133_pdest;
wire         io_diffCommits_info_133_rfWen;
wire         io_diffCommits_info_133_fpWen;
wire         io_diffCommits_info_133_vecWen;
wire         io_diffCommits_info_133_v0Wen;
wire         io_diffCommits_info_133_vlWen;
wire [5:0]   io_diffCommits_info_134_ldest;
wire [7:0]   io_diffCommits_info_134_pdest;
wire         io_diffCommits_info_134_rfWen;
wire         io_diffCommits_info_134_fpWen;
wire         io_diffCommits_info_134_vecWen;
wire         io_diffCommits_info_134_v0Wen;
wire         io_diffCommits_info_134_vlWen;
wire [5:0]   io_diffCommits_info_135_ldest;
wire [7:0]   io_diffCommits_info_135_pdest;
wire         io_diffCommits_info_135_rfWen;
wire         io_diffCommits_info_135_fpWen;
wire         io_diffCommits_info_135_vecWen;
wire         io_diffCommits_info_135_v0Wen;
wire         io_diffCommits_info_135_vlWen;
wire [5:0]   io_diffCommits_info_136_ldest;
wire [7:0]   io_diffCommits_info_136_pdest;
wire         io_diffCommits_info_136_rfWen;
wire         io_diffCommits_info_136_fpWen;
wire         io_diffCommits_info_136_vecWen;
wire         io_diffCommits_info_136_v0Wen;
wire         io_diffCommits_info_136_vlWen;
wire [5:0]   io_diffCommits_info_137_ldest;
wire [7:0]   io_diffCommits_info_137_pdest;
wire         io_diffCommits_info_137_rfWen;
wire         io_diffCommits_info_137_fpWen;
wire         io_diffCommits_info_137_vecWen;
wire         io_diffCommits_info_137_v0Wen;
wire         io_diffCommits_info_137_vlWen;
wire [5:0]   io_diffCommits_info_138_ldest;
wire [7:0]   io_diffCommits_info_138_pdest;
wire         io_diffCommits_info_138_rfWen;
wire         io_diffCommits_info_138_fpWen;
wire         io_diffCommits_info_138_vecWen;
wire         io_diffCommits_info_138_v0Wen;
wire         io_diffCommits_info_138_vlWen;
wire [5:0]   io_diffCommits_info_139_ldest;
wire [7:0]   io_diffCommits_info_139_pdest;
wire         io_diffCommits_info_139_rfWen;
wire         io_diffCommits_info_139_fpWen;
wire         io_diffCommits_info_139_vecWen;
wire         io_diffCommits_info_139_v0Wen;
wire         io_diffCommits_info_139_vlWen;
wire [5:0]   io_diffCommits_info_140_ldest;
wire [7:0]   io_diffCommits_info_140_pdest;
wire         io_diffCommits_info_140_rfWen;
wire         io_diffCommits_info_140_fpWen;
wire         io_diffCommits_info_140_vecWen;
wire         io_diffCommits_info_140_v0Wen;
wire         io_diffCommits_info_140_vlWen;
wire [5:0]   io_diffCommits_info_141_ldest;
wire [7:0]   io_diffCommits_info_141_pdest;
wire         io_diffCommits_info_141_rfWen;
wire         io_diffCommits_info_141_fpWen;
wire         io_diffCommits_info_141_vecWen;
wire         io_diffCommits_info_141_v0Wen;
wire         io_diffCommits_info_141_vlWen;
wire [5:0]   io_diffCommits_info_142_ldest;
wire [7:0]   io_diffCommits_info_142_pdest;
wire         io_diffCommits_info_142_rfWen;
wire         io_diffCommits_info_142_fpWen;
wire         io_diffCommits_info_142_vecWen;
wire         io_diffCommits_info_142_v0Wen;
wire         io_diffCommits_info_142_vlWen;
wire [5:0]   io_diffCommits_info_143_ldest;
wire [7:0]   io_diffCommits_info_143_pdest;
wire         io_diffCommits_info_143_rfWen;
wire         io_diffCommits_info_143_fpWen;
wire         io_diffCommits_info_143_vecWen;
wire         io_diffCommits_info_143_v0Wen;
wire         io_diffCommits_info_143_vlWen;
wire [5:0]   io_diffCommits_info_144_ldest;
wire [7:0]   io_diffCommits_info_144_pdest;
wire         io_diffCommits_info_144_rfWen;
wire         io_diffCommits_info_144_fpWen;
wire         io_diffCommits_info_144_vecWen;
wire         io_diffCommits_info_144_v0Wen;
wire         io_diffCommits_info_144_vlWen;
wire [5:0]   io_diffCommits_info_145_ldest;
wire [7:0]   io_diffCommits_info_145_pdest;
wire         io_diffCommits_info_145_rfWen;
wire         io_diffCommits_info_145_fpWen;
wire         io_diffCommits_info_145_vecWen;
wire         io_diffCommits_info_145_v0Wen;
wire         io_diffCommits_info_145_vlWen;
wire [5:0]   io_diffCommits_info_146_ldest;
wire [7:0]   io_diffCommits_info_146_pdest;
wire         io_diffCommits_info_146_rfWen;
wire         io_diffCommits_info_146_fpWen;
wire         io_diffCommits_info_146_vecWen;
wire         io_diffCommits_info_146_v0Wen;
wire         io_diffCommits_info_146_vlWen;
wire [5:0]   io_diffCommits_info_147_ldest;
wire [7:0]   io_diffCommits_info_147_pdest;
wire         io_diffCommits_info_147_rfWen;
wire         io_diffCommits_info_147_fpWen;
wire         io_diffCommits_info_147_vecWen;
wire         io_diffCommits_info_147_v0Wen;
wire         io_diffCommits_info_147_vlWen;
wire [5:0]   io_diffCommits_info_148_ldest;
wire [7:0]   io_diffCommits_info_148_pdest;
wire         io_diffCommits_info_148_rfWen;
wire         io_diffCommits_info_148_fpWen;
wire         io_diffCommits_info_148_vecWen;
wire         io_diffCommits_info_148_v0Wen;
wire         io_diffCommits_info_148_vlWen;
wire [5:0]   io_diffCommits_info_149_ldest;
wire [7:0]   io_diffCommits_info_149_pdest;
wire         io_diffCommits_info_149_rfWen;
wire         io_diffCommits_info_149_fpWen;
wire         io_diffCommits_info_149_vecWen;
wire         io_diffCommits_info_149_v0Wen;
wire         io_diffCommits_info_149_vlWen;
wire [5:0]   io_diffCommits_info_150_ldest;
wire [7:0]   io_diffCommits_info_150_pdest;
wire         io_diffCommits_info_150_rfWen;
wire         io_diffCommits_info_150_fpWen;
wire         io_diffCommits_info_150_vecWen;
wire         io_diffCommits_info_150_v0Wen;
wire         io_diffCommits_info_150_vlWen;
wire [5:0]   io_diffCommits_info_151_ldest;
wire [7:0]   io_diffCommits_info_151_pdest;
wire         io_diffCommits_info_151_rfWen;
wire         io_diffCommits_info_151_fpWen;
wire         io_diffCommits_info_151_vecWen;
wire         io_diffCommits_info_151_v0Wen;
wire         io_diffCommits_info_151_vlWen;
wire [5:0]   io_diffCommits_info_152_ldest;
wire [7:0]   io_diffCommits_info_152_pdest;
wire         io_diffCommits_info_152_rfWen;
wire         io_diffCommits_info_152_fpWen;
wire         io_diffCommits_info_152_vecWen;
wire         io_diffCommits_info_152_v0Wen;
wire         io_diffCommits_info_152_vlWen;
wire [5:0]   io_diffCommits_info_153_ldest;
wire [7:0]   io_diffCommits_info_153_pdest;
wire         io_diffCommits_info_153_rfWen;
wire         io_diffCommits_info_153_fpWen;
wire         io_diffCommits_info_153_vecWen;
wire         io_diffCommits_info_153_v0Wen;
wire         io_diffCommits_info_153_vlWen;
wire [5:0]   io_diffCommits_info_154_ldest;
wire [7:0]   io_diffCommits_info_154_pdest;
wire         io_diffCommits_info_154_rfWen;
wire         io_diffCommits_info_154_fpWen;
wire         io_diffCommits_info_154_vecWen;
wire         io_diffCommits_info_154_v0Wen;
wire         io_diffCommits_info_154_vlWen;
wire [5:0]   io_diffCommits_info_155_ldest;
wire [7:0]   io_diffCommits_info_155_pdest;
wire         io_diffCommits_info_155_rfWen;
wire         io_diffCommits_info_155_fpWen;
wire         io_diffCommits_info_155_vecWen;
wire         io_diffCommits_info_155_v0Wen;
wire         io_diffCommits_info_155_vlWen;
wire [5:0]   io_diffCommits_info_156_ldest;
wire [7:0]   io_diffCommits_info_156_pdest;
wire         io_diffCommits_info_156_rfWen;
wire         io_diffCommits_info_156_fpWen;
wire         io_diffCommits_info_156_vecWen;
wire         io_diffCommits_info_156_v0Wen;
wire         io_diffCommits_info_156_vlWen;
wire [5:0]   io_diffCommits_info_157_ldest;
wire [7:0]   io_diffCommits_info_157_pdest;
wire         io_diffCommits_info_157_rfWen;
wire         io_diffCommits_info_157_fpWen;
wire         io_diffCommits_info_157_vecWen;
wire         io_diffCommits_info_157_v0Wen;
wire         io_diffCommits_info_157_vlWen;
wire [5:0]   io_diffCommits_info_158_ldest;
wire [7:0]   io_diffCommits_info_158_pdest;
wire         io_diffCommits_info_158_rfWen;
wire         io_diffCommits_info_158_fpWen;
wire         io_diffCommits_info_158_vecWen;
wire         io_diffCommits_info_158_v0Wen;
wire         io_diffCommits_info_158_vlWen;
wire [5:0]   io_diffCommits_info_159_ldest;
wire [7:0]   io_diffCommits_info_159_pdest;
wire         io_diffCommits_info_159_rfWen;
wire         io_diffCommits_info_159_fpWen;
wire         io_diffCommits_info_159_vecWen;
wire         io_diffCommits_info_159_v0Wen;
wire         io_diffCommits_info_159_vlWen;
wire [5:0]   io_diffCommits_info_160_ldest;
wire [7:0]   io_diffCommits_info_160_pdest;
wire         io_diffCommits_info_160_rfWen;
wire         io_diffCommits_info_160_fpWen;
wire         io_diffCommits_info_160_vecWen;
wire         io_diffCommits_info_160_v0Wen;
wire         io_diffCommits_info_160_vlWen;
wire [5:0]   io_diffCommits_info_161_ldest;
wire [7:0]   io_diffCommits_info_161_pdest;
wire         io_diffCommits_info_161_rfWen;
wire         io_diffCommits_info_161_fpWen;
wire         io_diffCommits_info_161_vecWen;
wire         io_diffCommits_info_161_v0Wen;
wire         io_diffCommits_info_161_vlWen;
wire [5:0]   io_diffCommits_info_162_ldest;
wire [7:0]   io_diffCommits_info_162_pdest;
wire         io_diffCommits_info_162_rfWen;
wire         io_diffCommits_info_162_fpWen;
wire         io_diffCommits_info_162_vecWen;
wire         io_diffCommits_info_162_v0Wen;
wire         io_diffCommits_info_162_vlWen;
wire [5:0]   io_diffCommits_info_163_ldest;
wire [7:0]   io_diffCommits_info_163_pdest;
wire         io_diffCommits_info_163_rfWen;
wire         io_diffCommits_info_163_fpWen;
wire         io_diffCommits_info_163_vecWen;
wire         io_diffCommits_info_163_v0Wen;
wire         io_diffCommits_info_163_vlWen;
wire [5:0]   io_diffCommits_info_164_ldest;
wire [7:0]   io_diffCommits_info_164_pdest;
wire         io_diffCommits_info_164_rfWen;
wire         io_diffCommits_info_164_fpWen;
wire         io_diffCommits_info_164_vecWen;
wire         io_diffCommits_info_164_v0Wen;
wire         io_diffCommits_info_164_vlWen;
wire [5:0]   io_diffCommits_info_165_ldest;
wire [7:0]   io_diffCommits_info_165_pdest;
wire         io_diffCommits_info_165_rfWen;
wire         io_diffCommits_info_165_fpWen;
wire         io_diffCommits_info_165_vecWen;
wire         io_diffCommits_info_165_v0Wen;
wire         io_diffCommits_info_165_vlWen;
wire [5:0]   io_diffCommits_info_166_ldest;
wire [7:0]   io_diffCommits_info_166_pdest;
wire         io_diffCommits_info_166_rfWen;
wire         io_diffCommits_info_166_fpWen;
wire         io_diffCommits_info_166_vecWen;
wire         io_diffCommits_info_166_v0Wen;
wire         io_diffCommits_info_166_vlWen;
wire [5:0]   io_diffCommits_info_167_ldest;
wire [7:0]   io_diffCommits_info_167_pdest;
wire         io_diffCommits_info_167_rfWen;
wire         io_diffCommits_info_167_fpWen;
wire         io_diffCommits_info_167_vecWen;
wire         io_diffCommits_info_167_v0Wen;
wire         io_diffCommits_info_167_vlWen;
wire [5:0]   io_diffCommits_info_168_ldest;
wire [7:0]   io_diffCommits_info_168_pdest;
wire         io_diffCommits_info_168_rfWen;
wire         io_diffCommits_info_168_fpWen;
wire         io_diffCommits_info_168_vecWen;
wire         io_diffCommits_info_168_v0Wen;
wire         io_diffCommits_info_168_vlWen;
wire [5:0]   io_diffCommits_info_169_ldest;
wire [7:0]   io_diffCommits_info_169_pdest;
wire         io_diffCommits_info_169_rfWen;
wire         io_diffCommits_info_169_fpWen;
wire         io_diffCommits_info_169_vecWen;
wire         io_diffCommits_info_169_v0Wen;
wire         io_diffCommits_info_169_vlWen;
wire [5:0]   io_diffCommits_info_170_ldest;
wire [7:0]   io_diffCommits_info_170_pdest;
wire         io_diffCommits_info_170_rfWen;
wire         io_diffCommits_info_170_fpWen;
wire         io_diffCommits_info_170_vecWen;
wire         io_diffCommits_info_170_v0Wen;
wire         io_diffCommits_info_170_vlWen;
wire [5:0]   io_diffCommits_info_171_ldest;
wire [7:0]   io_diffCommits_info_171_pdest;
wire         io_diffCommits_info_171_rfWen;
wire         io_diffCommits_info_171_fpWen;
wire         io_diffCommits_info_171_vecWen;
wire         io_diffCommits_info_171_v0Wen;
wire         io_diffCommits_info_171_vlWen;
wire [5:0]   io_diffCommits_info_172_ldest;
wire [7:0]   io_diffCommits_info_172_pdest;
wire         io_diffCommits_info_172_rfWen;
wire         io_diffCommits_info_172_fpWen;
wire         io_diffCommits_info_172_vecWen;
wire         io_diffCommits_info_172_v0Wen;
wire         io_diffCommits_info_172_vlWen;
wire [5:0]   io_diffCommits_info_173_ldest;
wire [7:0]   io_diffCommits_info_173_pdest;
wire         io_diffCommits_info_173_rfWen;
wire         io_diffCommits_info_173_fpWen;
wire         io_diffCommits_info_173_vecWen;
wire         io_diffCommits_info_173_v0Wen;
wire         io_diffCommits_info_173_vlWen;
wire [5:0]   io_diffCommits_info_174_ldest;
wire [7:0]   io_diffCommits_info_174_pdest;
wire         io_diffCommits_info_174_rfWen;
wire         io_diffCommits_info_174_fpWen;
wire         io_diffCommits_info_174_vecWen;
wire         io_diffCommits_info_174_v0Wen;
wire         io_diffCommits_info_174_vlWen;
wire [5:0]   io_diffCommits_info_175_ldest;
wire [7:0]   io_diffCommits_info_175_pdest;
wire         io_diffCommits_info_175_rfWen;
wire         io_diffCommits_info_175_fpWen;
wire         io_diffCommits_info_175_vecWen;
wire         io_diffCommits_info_175_v0Wen;
wire         io_diffCommits_info_175_vlWen;
wire [5:0]   io_diffCommits_info_176_ldest;
wire [7:0]   io_diffCommits_info_176_pdest;
wire         io_diffCommits_info_176_rfWen;
wire         io_diffCommits_info_176_fpWen;
wire         io_diffCommits_info_176_vecWen;
wire         io_diffCommits_info_176_v0Wen;
wire         io_diffCommits_info_176_vlWen;
wire [5:0]   io_diffCommits_info_177_ldest;
wire [7:0]   io_diffCommits_info_177_pdest;
wire         io_diffCommits_info_177_rfWen;
wire         io_diffCommits_info_177_fpWen;
wire         io_diffCommits_info_177_vecWen;
wire         io_diffCommits_info_177_v0Wen;
wire         io_diffCommits_info_177_vlWen;
wire [5:0]   io_diffCommits_info_178_ldest;
wire [7:0]   io_diffCommits_info_178_pdest;
wire         io_diffCommits_info_178_rfWen;
wire         io_diffCommits_info_178_fpWen;
wire         io_diffCommits_info_178_vecWen;
wire         io_diffCommits_info_178_v0Wen;
wire         io_diffCommits_info_178_vlWen;
wire [5:0]   io_diffCommits_info_179_ldest;
wire [7:0]   io_diffCommits_info_179_pdest;
wire         io_diffCommits_info_179_rfWen;
wire         io_diffCommits_info_179_fpWen;
wire         io_diffCommits_info_179_vecWen;
wire         io_diffCommits_info_179_v0Wen;
wire         io_diffCommits_info_179_vlWen;
wire [5:0]   io_diffCommits_info_180_ldest;
wire [7:0]   io_diffCommits_info_180_pdest;
wire         io_diffCommits_info_180_rfWen;
wire         io_diffCommits_info_180_fpWen;
wire         io_diffCommits_info_180_vecWen;
wire         io_diffCommits_info_180_v0Wen;
wire         io_diffCommits_info_180_vlWen;
wire [5:0]   io_diffCommits_info_181_ldest;
wire [7:0]   io_diffCommits_info_181_pdest;
wire         io_diffCommits_info_181_rfWen;
wire         io_diffCommits_info_181_fpWen;
wire         io_diffCommits_info_181_vecWen;
wire         io_diffCommits_info_181_v0Wen;
wire         io_diffCommits_info_181_vlWen;
wire [5:0]   io_diffCommits_info_182_ldest;
wire [7:0]   io_diffCommits_info_182_pdest;
wire         io_diffCommits_info_182_rfWen;
wire         io_diffCommits_info_182_fpWen;
wire         io_diffCommits_info_182_vecWen;
wire         io_diffCommits_info_182_v0Wen;
wire         io_diffCommits_info_182_vlWen;
wire [5:0]   io_diffCommits_info_183_ldest;
wire [7:0]   io_diffCommits_info_183_pdest;
wire         io_diffCommits_info_183_rfWen;
wire         io_diffCommits_info_183_fpWen;
wire         io_diffCommits_info_183_vecWen;
wire         io_diffCommits_info_183_v0Wen;
wire         io_diffCommits_info_183_vlWen;
wire [5:0]   io_diffCommits_info_184_ldest;
wire [7:0]   io_diffCommits_info_184_pdest;
wire         io_diffCommits_info_184_rfWen;
wire         io_diffCommits_info_184_fpWen;
wire         io_diffCommits_info_184_vecWen;
wire         io_diffCommits_info_184_v0Wen;
wire         io_diffCommits_info_184_vlWen;
wire [5:0]   io_diffCommits_info_185_ldest;
wire [7:0]   io_diffCommits_info_185_pdest;
wire         io_diffCommits_info_185_rfWen;
wire         io_diffCommits_info_185_fpWen;
wire         io_diffCommits_info_185_vecWen;
wire         io_diffCommits_info_185_v0Wen;
wire         io_diffCommits_info_185_vlWen;
wire [5:0]   io_diffCommits_info_186_ldest;
wire [7:0]   io_diffCommits_info_186_pdest;
wire         io_diffCommits_info_186_rfWen;
wire         io_diffCommits_info_186_fpWen;
wire         io_diffCommits_info_186_vecWen;
wire         io_diffCommits_info_186_v0Wen;
wire         io_diffCommits_info_186_vlWen;
wire [5:0]   io_diffCommits_info_187_ldest;
wire [7:0]   io_diffCommits_info_187_pdest;
wire         io_diffCommits_info_187_rfWen;
wire         io_diffCommits_info_187_fpWen;
wire         io_diffCommits_info_187_vecWen;
wire         io_diffCommits_info_187_v0Wen;
wire         io_diffCommits_info_187_vlWen;
wire [5:0]   io_diffCommits_info_188_ldest;
wire [7:0]   io_diffCommits_info_188_pdest;
wire         io_diffCommits_info_188_rfWen;
wire         io_diffCommits_info_188_fpWen;
wire         io_diffCommits_info_188_vecWen;
wire         io_diffCommits_info_188_v0Wen;
wire         io_diffCommits_info_188_vlWen;
wire [5:0]   io_diffCommits_info_189_ldest;
wire [7:0]   io_diffCommits_info_189_pdest;
wire         io_diffCommits_info_189_rfWen;
wire         io_diffCommits_info_189_fpWen;
wire         io_diffCommits_info_189_vecWen;
wire         io_diffCommits_info_189_v0Wen;
wire         io_diffCommits_info_189_vlWen;
wire [5:0]   io_diffCommits_info_190_ldest;
wire [7:0]   io_diffCommits_info_190_pdest;
wire         io_diffCommits_info_190_rfWen;
wire         io_diffCommits_info_190_fpWen;
wire         io_diffCommits_info_190_vecWen;
wire         io_diffCommits_info_190_v0Wen;
wire         io_diffCommits_info_190_vlWen;
wire [5:0]   io_diffCommits_info_191_ldest;
wire [7:0]   io_diffCommits_info_191_pdest;
wire         io_diffCommits_info_191_rfWen;
wire         io_diffCommits_info_191_fpWen;
wire         io_diffCommits_info_191_vecWen;
wire         io_diffCommits_info_191_v0Wen;
wire         io_diffCommits_info_191_vlWen;
wire [5:0]   io_diffCommits_info_192_ldest;
wire [7:0]   io_diffCommits_info_192_pdest;
wire         io_diffCommits_info_192_rfWen;
wire         io_diffCommits_info_192_fpWen;
wire         io_diffCommits_info_192_vecWen;
wire         io_diffCommits_info_192_v0Wen;
wire         io_diffCommits_info_192_vlWen;
wire [5:0]   io_diffCommits_info_193_ldest;
wire [7:0]   io_diffCommits_info_193_pdest;
wire         io_diffCommits_info_193_rfWen;
wire         io_diffCommits_info_193_fpWen;
wire         io_diffCommits_info_193_vecWen;
wire         io_diffCommits_info_193_v0Wen;
wire         io_diffCommits_info_193_vlWen;
wire [5:0]   io_diffCommits_info_194_ldest;
wire [7:0]   io_diffCommits_info_194_pdest;
wire         io_diffCommits_info_194_rfWen;
wire         io_diffCommits_info_194_fpWen;
wire         io_diffCommits_info_194_vecWen;
wire         io_diffCommits_info_194_v0Wen;
wire         io_diffCommits_info_194_vlWen;
wire [5:0]   io_diffCommits_info_195_ldest;
wire [7:0]   io_diffCommits_info_195_pdest;
wire         io_diffCommits_info_195_rfWen;
wire         io_diffCommits_info_195_fpWen;
wire         io_diffCommits_info_195_vecWen;
wire         io_diffCommits_info_195_v0Wen;
wire         io_diffCommits_info_195_vlWen;
wire [5:0]   io_diffCommits_info_196_ldest;
wire [7:0]   io_diffCommits_info_196_pdest;
wire         io_diffCommits_info_196_rfWen;
wire         io_diffCommits_info_196_fpWen;
wire         io_diffCommits_info_196_vecWen;
wire         io_diffCommits_info_196_v0Wen;
wire         io_diffCommits_info_196_vlWen;
wire [5:0]   io_diffCommits_info_197_ldest;
wire [7:0]   io_diffCommits_info_197_pdest;
wire         io_diffCommits_info_197_rfWen;
wire         io_diffCommits_info_197_fpWen;
wire         io_diffCommits_info_197_vecWen;
wire         io_diffCommits_info_197_v0Wen;
wire         io_diffCommits_info_197_vlWen;
wire [5:0]   io_diffCommits_info_198_ldest;
wire [7:0]   io_diffCommits_info_198_pdest;
wire         io_diffCommits_info_198_rfWen;
wire         io_diffCommits_info_198_fpWen;
wire         io_diffCommits_info_198_vecWen;
wire         io_diffCommits_info_198_v0Wen;
wire         io_diffCommits_info_198_vlWen;
wire [5:0]   io_diffCommits_info_199_ldest;
wire [7:0]   io_diffCommits_info_199_pdest;
wire         io_diffCommits_info_199_rfWen;
wire         io_diffCommits_info_199_fpWen;
wire         io_diffCommits_info_199_vecWen;
wire         io_diffCommits_info_199_v0Wen;
wire         io_diffCommits_info_199_vlWen;
wire [5:0]   io_diffCommits_info_200_ldest;
wire [7:0]   io_diffCommits_info_200_pdest;
wire         io_diffCommits_info_200_rfWen;
wire         io_diffCommits_info_200_fpWen;
wire         io_diffCommits_info_200_vecWen;
wire         io_diffCommits_info_200_v0Wen;
wire         io_diffCommits_info_200_vlWen;
wire [5:0]   io_diffCommits_info_201_ldest;
wire [7:0]   io_diffCommits_info_201_pdest;
wire         io_diffCommits_info_201_rfWen;
wire         io_diffCommits_info_201_fpWen;
wire         io_diffCommits_info_201_vecWen;
wire         io_diffCommits_info_201_v0Wen;
wire         io_diffCommits_info_201_vlWen;
wire [5:0]   io_diffCommits_info_202_ldest;
wire [7:0]   io_diffCommits_info_202_pdest;
wire         io_diffCommits_info_202_rfWen;
wire         io_diffCommits_info_202_fpWen;
wire         io_diffCommits_info_202_vecWen;
wire         io_diffCommits_info_202_v0Wen;
wire         io_diffCommits_info_202_vlWen;
wire [5:0]   io_diffCommits_info_203_ldest;
wire [7:0]   io_diffCommits_info_203_pdest;
wire         io_diffCommits_info_203_rfWen;
wire         io_diffCommits_info_203_fpWen;
wire         io_diffCommits_info_203_vecWen;
wire         io_diffCommits_info_203_v0Wen;
wire         io_diffCommits_info_203_vlWen;
wire [5:0]   io_diffCommits_info_204_ldest;
wire [7:0]   io_diffCommits_info_204_pdest;
wire         io_diffCommits_info_204_rfWen;
wire         io_diffCommits_info_204_fpWen;
wire         io_diffCommits_info_204_vecWen;
wire         io_diffCommits_info_204_v0Wen;
wire         io_diffCommits_info_204_vlWen;
wire [5:0]   io_diffCommits_info_205_ldest;
wire [7:0]   io_diffCommits_info_205_pdest;
wire         io_diffCommits_info_205_rfWen;
wire         io_diffCommits_info_205_fpWen;
wire         io_diffCommits_info_205_vecWen;
wire         io_diffCommits_info_205_v0Wen;
wire         io_diffCommits_info_205_vlWen;
wire [5:0]   io_diffCommits_info_206_ldest;
wire [7:0]   io_diffCommits_info_206_pdest;
wire         io_diffCommits_info_206_rfWen;
wire         io_diffCommits_info_206_fpWen;
wire         io_diffCommits_info_206_vecWen;
wire         io_diffCommits_info_206_v0Wen;
wire         io_diffCommits_info_206_vlWen;
wire [5:0]   io_diffCommits_info_207_ldest;
wire [7:0]   io_diffCommits_info_207_pdest;
wire         io_diffCommits_info_207_rfWen;
wire         io_diffCommits_info_207_fpWen;
wire         io_diffCommits_info_207_vecWen;
wire         io_diffCommits_info_207_v0Wen;
wire         io_diffCommits_info_207_vlWen;
wire [5:0]   io_diffCommits_info_208_ldest;
wire [7:0]   io_diffCommits_info_208_pdest;
wire         io_diffCommits_info_208_rfWen;
wire         io_diffCommits_info_208_fpWen;
wire         io_diffCommits_info_208_vecWen;
wire         io_diffCommits_info_208_v0Wen;
wire         io_diffCommits_info_208_vlWen;
wire [5:0]   io_diffCommits_info_209_ldest;
wire [7:0]   io_diffCommits_info_209_pdest;
wire         io_diffCommits_info_209_rfWen;
wire         io_diffCommits_info_209_fpWen;
wire         io_diffCommits_info_209_vecWen;
wire         io_diffCommits_info_209_v0Wen;
wire         io_diffCommits_info_209_vlWen;
wire [5:0]   io_diffCommits_info_210_ldest;
wire [7:0]   io_diffCommits_info_210_pdest;
wire         io_diffCommits_info_210_rfWen;
wire         io_diffCommits_info_210_fpWen;
wire         io_diffCommits_info_210_vecWen;
wire         io_diffCommits_info_210_v0Wen;
wire         io_diffCommits_info_210_vlWen;
wire [5:0]   io_diffCommits_info_211_ldest;
wire [7:0]   io_diffCommits_info_211_pdest;
wire         io_diffCommits_info_211_rfWen;
wire         io_diffCommits_info_211_fpWen;
wire         io_diffCommits_info_211_vecWen;
wire         io_diffCommits_info_211_v0Wen;
wire         io_diffCommits_info_211_vlWen;
wire [5:0]   io_diffCommits_info_212_ldest;
wire [7:0]   io_diffCommits_info_212_pdest;
wire         io_diffCommits_info_212_rfWen;
wire         io_diffCommits_info_212_fpWen;
wire         io_diffCommits_info_212_vecWen;
wire         io_diffCommits_info_212_v0Wen;
wire         io_diffCommits_info_212_vlWen;
wire [5:0]   io_diffCommits_info_213_ldest;
wire [7:0]   io_diffCommits_info_213_pdest;
wire         io_diffCommits_info_213_rfWen;
wire         io_diffCommits_info_213_fpWen;
wire         io_diffCommits_info_213_vecWen;
wire         io_diffCommits_info_213_v0Wen;
wire         io_diffCommits_info_213_vlWen;
wire [5:0]   io_diffCommits_info_214_ldest;
wire [7:0]   io_diffCommits_info_214_pdest;
wire         io_diffCommits_info_214_rfWen;
wire         io_diffCommits_info_214_fpWen;
wire         io_diffCommits_info_214_vecWen;
wire         io_diffCommits_info_214_v0Wen;
wire         io_diffCommits_info_214_vlWen;
wire [5:0]   io_diffCommits_info_215_ldest;
wire [7:0]   io_diffCommits_info_215_pdest;
wire         io_diffCommits_info_215_rfWen;
wire         io_diffCommits_info_215_fpWen;
wire         io_diffCommits_info_215_vecWen;
wire         io_diffCommits_info_215_v0Wen;
wire         io_diffCommits_info_215_vlWen;
wire [5:0]   io_diffCommits_info_216_ldest;
wire [7:0]   io_diffCommits_info_216_pdest;
wire         io_diffCommits_info_216_rfWen;
wire         io_diffCommits_info_216_fpWen;
wire         io_diffCommits_info_216_vecWen;
wire         io_diffCommits_info_216_v0Wen;
wire         io_diffCommits_info_216_vlWen;
wire [5:0]   io_diffCommits_info_217_ldest;
wire [7:0]   io_diffCommits_info_217_pdest;
wire         io_diffCommits_info_217_rfWen;
wire         io_diffCommits_info_217_fpWen;
wire         io_diffCommits_info_217_vecWen;
wire         io_diffCommits_info_217_v0Wen;
wire         io_diffCommits_info_217_vlWen;
wire [5:0]   io_diffCommits_info_218_ldest;
wire [7:0]   io_diffCommits_info_218_pdest;
wire         io_diffCommits_info_218_rfWen;
wire         io_diffCommits_info_218_fpWen;
wire         io_diffCommits_info_218_vecWen;
wire         io_diffCommits_info_218_v0Wen;
wire         io_diffCommits_info_218_vlWen;
wire [5:0]   io_diffCommits_info_219_ldest;
wire [7:0]   io_diffCommits_info_219_pdest;
wire         io_diffCommits_info_219_rfWen;
wire         io_diffCommits_info_219_fpWen;
wire         io_diffCommits_info_219_vecWen;
wire         io_diffCommits_info_219_v0Wen;
wire         io_diffCommits_info_219_vlWen;
wire [5:0]   io_diffCommits_info_220_ldest;
wire [7:0]   io_diffCommits_info_220_pdest;
wire         io_diffCommits_info_220_rfWen;
wire         io_diffCommits_info_220_fpWen;
wire         io_diffCommits_info_220_vecWen;
wire         io_diffCommits_info_220_v0Wen;
wire         io_diffCommits_info_220_vlWen;
wire [5:0]   io_diffCommits_info_221_ldest;
wire [7:0]   io_diffCommits_info_221_pdest;
wire         io_diffCommits_info_221_rfWen;
wire         io_diffCommits_info_221_fpWen;
wire         io_diffCommits_info_221_vecWen;
wire         io_diffCommits_info_221_v0Wen;
wire         io_diffCommits_info_221_vlWen;
wire [5:0]   io_diffCommits_info_222_ldest;
wire [7:0]   io_diffCommits_info_222_pdest;
wire         io_diffCommits_info_222_rfWen;
wire         io_diffCommits_info_222_fpWen;
wire         io_diffCommits_info_222_vecWen;
wire         io_diffCommits_info_222_v0Wen;
wire         io_diffCommits_info_222_vlWen;
wire [5:0]   io_diffCommits_info_223_ldest;
wire [7:0]   io_diffCommits_info_223_pdest;
wire         io_diffCommits_info_223_rfWen;
wire         io_diffCommits_info_223_fpWen;
wire         io_diffCommits_info_223_vecWen;
wire         io_diffCommits_info_223_v0Wen;
wire         io_diffCommits_info_223_vlWen;
wire [5:0]   io_diffCommits_info_224_ldest;
wire [7:0]   io_diffCommits_info_224_pdest;
wire         io_diffCommits_info_224_rfWen;
wire         io_diffCommits_info_224_fpWen;
wire         io_diffCommits_info_224_vecWen;
wire         io_diffCommits_info_224_v0Wen;
wire         io_diffCommits_info_224_vlWen;
wire [5:0]   io_diffCommits_info_225_ldest;
wire [7:0]   io_diffCommits_info_225_pdest;
wire         io_diffCommits_info_225_rfWen;
wire         io_diffCommits_info_225_fpWen;
wire         io_diffCommits_info_225_vecWen;
wire         io_diffCommits_info_225_v0Wen;
wire         io_diffCommits_info_225_vlWen;
wire [5:0]   io_diffCommits_info_226_ldest;
wire [7:0]   io_diffCommits_info_226_pdest;
wire         io_diffCommits_info_226_rfWen;
wire         io_diffCommits_info_226_fpWen;
wire         io_diffCommits_info_226_vecWen;
wire         io_diffCommits_info_226_v0Wen;
wire         io_diffCommits_info_226_vlWen;
wire [5:0]   io_diffCommits_info_227_ldest;
wire [7:0]   io_diffCommits_info_227_pdest;
wire         io_diffCommits_info_227_rfWen;
wire         io_diffCommits_info_227_fpWen;
wire         io_diffCommits_info_227_vecWen;
wire         io_diffCommits_info_227_v0Wen;
wire         io_diffCommits_info_227_vlWen;
wire [5:0]   io_diffCommits_info_228_ldest;
wire [7:0]   io_diffCommits_info_228_pdest;
wire         io_diffCommits_info_228_rfWen;
wire         io_diffCommits_info_228_fpWen;
wire         io_diffCommits_info_228_vecWen;
wire         io_diffCommits_info_228_v0Wen;
wire         io_diffCommits_info_228_vlWen;
wire [5:0]   io_diffCommits_info_229_ldest;
wire [7:0]   io_diffCommits_info_229_pdest;
wire         io_diffCommits_info_229_rfWen;
wire         io_diffCommits_info_229_fpWen;
wire         io_diffCommits_info_229_vecWen;
wire         io_diffCommits_info_229_v0Wen;
wire         io_diffCommits_info_229_vlWen;
wire [5:0]   io_diffCommits_info_230_ldest;
wire [7:0]   io_diffCommits_info_230_pdest;
wire         io_diffCommits_info_230_rfWen;
wire         io_diffCommits_info_230_fpWen;
wire         io_diffCommits_info_230_vecWen;
wire         io_diffCommits_info_230_v0Wen;
wire         io_diffCommits_info_230_vlWen;
wire [5:0]   io_diffCommits_info_231_ldest;
wire [7:0]   io_diffCommits_info_231_pdest;
wire         io_diffCommits_info_231_rfWen;
wire         io_diffCommits_info_231_fpWen;
wire         io_diffCommits_info_231_vecWen;
wire         io_diffCommits_info_231_v0Wen;
wire         io_diffCommits_info_231_vlWen;
wire [5:0]   io_diffCommits_info_232_ldest;
wire [7:0]   io_diffCommits_info_232_pdest;
wire         io_diffCommits_info_232_rfWen;
wire         io_diffCommits_info_232_fpWen;
wire         io_diffCommits_info_232_vecWen;
wire         io_diffCommits_info_232_v0Wen;
wire         io_diffCommits_info_232_vlWen;
wire [5:0]   io_diffCommits_info_233_ldest;
wire [7:0]   io_diffCommits_info_233_pdest;
wire         io_diffCommits_info_233_rfWen;
wire         io_diffCommits_info_233_fpWen;
wire         io_diffCommits_info_233_vecWen;
wire         io_diffCommits_info_233_v0Wen;
wire         io_diffCommits_info_233_vlWen;
wire [5:0]   io_diffCommits_info_234_ldest;
wire [7:0]   io_diffCommits_info_234_pdest;
wire         io_diffCommits_info_234_rfWen;
wire         io_diffCommits_info_234_fpWen;
wire         io_diffCommits_info_234_vecWen;
wire         io_diffCommits_info_234_v0Wen;
wire         io_diffCommits_info_234_vlWen;
wire [5:0]   io_diffCommits_info_235_ldest;
wire [7:0]   io_diffCommits_info_235_pdest;
wire         io_diffCommits_info_235_rfWen;
wire         io_diffCommits_info_235_fpWen;
wire         io_diffCommits_info_235_vecWen;
wire         io_diffCommits_info_235_v0Wen;
wire         io_diffCommits_info_235_vlWen;
wire [5:0]   io_diffCommits_info_236_ldest;
wire [7:0]   io_diffCommits_info_236_pdest;
wire         io_diffCommits_info_236_rfWen;
wire         io_diffCommits_info_236_fpWen;
wire         io_diffCommits_info_236_vecWen;
wire         io_diffCommits_info_236_v0Wen;
wire         io_diffCommits_info_236_vlWen;
wire [5:0]   io_diffCommits_info_237_ldest;
wire [7:0]   io_diffCommits_info_237_pdest;
wire         io_diffCommits_info_237_rfWen;
wire         io_diffCommits_info_237_fpWen;
wire         io_diffCommits_info_237_vecWen;
wire         io_diffCommits_info_237_v0Wen;
wire         io_diffCommits_info_237_vlWen;
wire [5:0]   io_diffCommits_info_238_ldest;
wire [7:0]   io_diffCommits_info_238_pdest;
wire         io_diffCommits_info_238_rfWen;
wire         io_diffCommits_info_238_fpWen;
wire         io_diffCommits_info_238_vecWen;
wire         io_diffCommits_info_238_v0Wen;
wire         io_diffCommits_info_238_vlWen;
wire [5:0]   io_diffCommits_info_239_ldest;
wire [7:0]   io_diffCommits_info_239_pdest;
wire         io_diffCommits_info_239_rfWen;
wire         io_diffCommits_info_239_fpWen;
wire         io_diffCommits_info_239_vecWen;
wire         io_diffCommits_info_239_v0Wen;
wire         io_diffCommits_info_239_vlWen;
wire [5:0]   io_diffCommits_info_240_ldest;
wire [7:0]   io_diffCommits_info_240_pdest;
wire         io_diffCommits_info_240_rfWen;
wire         io_diffCommits_info_240_fpWen;
wire         io_diffCommits_info_240_vecWen;
wire         io_diffCommits_info_240_v0Wen;
wire         io_diffCommits_info_240_vlWen;
wire [5:0]   io_diffCommits_info_241_ldest;
wire [7:0]   io_diffCommits_info_241_pdest;
wire         io_diffCommits_info_241_rfWen;
wire         io_diffCommits_info_241_fpWen;
wire         io_diffCommits_info_241_vecWen;
wire         io_diffCommits_info_241_v0Wen;
wire         io_diffCommits_info_241_vlWen;
wire [5:0]   io_diffCommits_info_242_ldest;
wire [7:0]   io_diffCommits_info_242_pdest;
wire         io_diffCommits_info_242_rfWen;
wire         io_diffCommits_info_242_fpWen;
wire         io_diffCommits_info_242_vecWen;
wire         io_diffCommits_info_242_v0Wen;
wire         io_diffCommits_info_242_vlWen;
wire [5:0]   io_diffCommits_info_243_ldest;
wire [7:0]   io_diffCommits_info_243_pdest;
wire         io_diffCommits_info_243_rfWen;
wire         io_diffCommits_info_243_fpWen;
wire         io_diffCommits_info_243_vecWen;
wire         io_diffCommits_info_243_v0Wen;
wire         io_diffCommits_info_243_vlWen;
wire [5:0]   io_diffCommits_info_244_ldest;
wire [7:0]   io_diffCommits_info_244_pdest;
wire         io_diffCommits_info_244_rfWen;
wire         io_diffCommits_info_244_fpWen;
wire         io_diffCommits_info_244_vecWen;
wire         io_diffCommits_info_244_v0Wen;
wire         io_diffCommits_info_244_vlWen;
wire [5:0]   io_diffCommits_info_245_ldest;
wire [7:0]   io_diffCommits_info_245_pdest;
wire         io_diffCommits_info_245_rfWen;
wire         io_diffCommits_info_245_fpWen;
wire         io_diffCommits_info_245_vecWen;
wire         io_diffCommits_info_245_v0Wen;
wire         io_diffCommits_info_245_vlWen;
wire [5:0]   io_diffCommits_info_246_ldest;
wire [7:0]   io_diffCommits_info_246_pdest;
wire         io_diffCommits_info_246_rfWen;
wire         io_diffCommits_info_246_fpWen;
wire         io_diffCommits_info_246_vecWen;
wire         io_diffCommits_info_246_v0Wen;
wire         io_diffCommits_info_246_vlWen;
wire [5:0]   io_diffCommits_info_247_ldest;
wire [7:0]   io_diffCommits_info_247_pdest;
wire         io_diffCommits_info_247_rfWen;
wire         io_diffCommits_info_247_fpWen;
wire         io_diffCommits_info_247_vecWen;
wire         io_diffCommits_info_247_v0Wen;
wire         io_diffCommits_info_247_vlWen;
wire [5:0]   io_diffCommits_info_248_ldest;
wire [7:0]   io_diffCommits_info_248_pdest;
wire         io_diffCommits_info_248_rfWen;
wire         io_diffCommits_info_248_fpWen;
wire         io_diffCommits_info_248_vecWen;
wire         io_diffCommits_info_248_v0Wen;
wire         io_diffCommits_info_248_vlWen;
wire [5:0]   io_diffCommits_info_249_ldest;
wire [7:0]   io_diffCommits_info_249_pdest;
wire         io_diffCommits_info_249_rfWen;
wire         io_diffCommits_info_249_fpWen;
wire         io_diffCommits_info_249_vecWen;
wire         io_diffCommits_info_249_v0Wen;
wire         io_diffCommits_info_249_vlWen;
wire [5:0]   io_diffCommits_info_250_ldest;
wire [7:0]   io_diffCommits_info_250_pdest;
wire         io_diffCommits_info_250_rfWen;
wire         io_diffCommits_info_250_fpWen;
wire         io_diffCommits_info_250_vecWen;
wire         io_diffCommits_info_250_v0Wen;
wire         io_diffCommits_info_250_vlWen;
wire [5:0]   io_diffCommits_info_251_ldest;
wire [7:0]   io_diffCommits_info_251_pdest;
wire         io_diffCommits_info_251_rfWen;
wire         io_diffCommits_info_251_fpWen;
wire         io_diffCommits_info_251_vecWen;
wire         io_diffCommits_info_251_v0Wen;
wire         io_diffCommits_info_251_vlWen;
wire [5:0]   io_diffCommits_info_252_ldest;
wire [7:0]   io_diffCommits_info_252_pdest;
wire         io_diffCommits_info_252_rfWen;
wire         io_diffCommits_info_252_fpWen;
wire         io_diffCommits_info_252_vecWen;
wire         io_diffCommits_info_252_v0Wen;
wire         io_diffCommits_info_252_vlWen;
wire [5:0]   io_diffCommits_info_253_ldest;
wire [7:0]   io_diffCommits_info_253_pdest;
wire         io_diffCommits_info_253_rfWen;
wire         io_diffCommits_info_253_fpWen;
wire         io_diffCommits_info_253_vecWen;
wire         io_diffCommits_info_253_v0Wen;
wire         io_diffCommits_info_253_vlWen;
wire [5:0]   io_diffCommits_info_254_ldest;
wire [7:0]   io_diffCommits_info_254_pdest;
wire         io_diffCommits_info_254_rfWen;
wire         io_diffCommits_info_254_fpWen;
wire         io_diffCommits_info_254_vecWen;
wire         io_diffCommits_info_254_v0Wen;
wire         io_diffCommits_info_254_vlWen;
wire [5:0]   io_diffCommits_info_255_ldest;
wire [7:0]   io_diffCommits_info_255_pdest;
wire [5:0]   io_diffCommits_info_256_ldest;
wire [7:0]   io_diffCommits_info_256_pdest;
wire [5:0]   io_diffCommits_info_257_ldest;
wire [7:0]   io_diffCommits_info_257_pdest;
wire [5:0]   io_diffCommits_info_258_ldest;
wire [7:0]   io_diffCommits_info_258_pdest;
wire [5:0]   io_diffCommits_info_259_ldest;
wire [7:0]   io_diffCommits_info_259_pdest;
wire [5:0]   io_diffCommits_info_260_ldest;
wire [7:0]   io_diffCommits_info_260_pdest;
wire [5:0]   io_diffCommits_info_261_ldest;
wire [7:0]   io_diffCommits_info_261_pdest;
wire [5:0]   io_diffCommits_info_262_ldest;
wire [7:0]   io_diffCommits_info_262_pdest;
wire [5:0]   io_diffCommits_info_263_ldest;
wire [7:0]   io_diffCommits_info_263_pdest;
wire [5:0]   io_diffCommits_info_264_ldest;
wire [7:0]   io_diffCommits_info_264_pdest;
wire [5:0]   io_diffCommits_info_265_ldest;
wire [7:0]   io_diffCommits_info_265_pdest;
wire [5:0]   io_diffCommits_info_266_ldest;
wire [7:0]   io_diffCommits_info_266_pdest;
wire [5:0]   io_diffCommits_info_267_ldest;
wire [7:0]   io_diffCommits_info_267_pdest;
wire [5:0]   io_diffCommits_info_268_ldest;
wire [7:0]   io_diffCommits_info_268_pdest;
wire [5:0]   io_diffCommits_info_269_ldest;
wire [7:0]   io_diffCommits_info_269_pdest;
wire [5:0]   io_diffCommits_info_270_ldest;
wire [7:0]   io_diffCommits_info_270_pdest;
wire [5:0]   io_diffCommits_info_271_ldest;
wire [7:0]   io_diffCommits_info_271_pdest;
wire [5:0]   io_diffCommits_info_272_ldest;
wire [7:0]   io_diffCommits_info_272_pdest;
wire [5:0]   io_diffCommits_info_273_ldest;
wire [7:0]   io_diffCommits_info_273_pdest;
wire [5:0]   io_diffCommits_info_274_ldest;
wire [7:0]   io_diffCommits_info_274_pdest;
wire [5:0]   io_diffCommits_info_275_ldest;
wire [7:0]   io_diffCommits_info_275_pdest;
wire [5:0]   io_diffCommits_info_276_ldest;
wire [7:0]   io_diffCommits_info_276_pdest;
wire [5:0]   io_diffCommits_info_277_ldest;
wire [7:0]   io_diffCommits_info_277_pdest;
wire [5:0]   io_diffCommits_info_278_ldest;
wire [7:0]   io_diffCommits_info_278_pdest;
wire [5:0]   io_diffCommits_info_279_ldest;
wire [7:0]   io_diffCommits_info_279_pdest;
wire [5:0]   io_diffCommits_info_280_ldest;
wire [7:0]   io_diffCommits_info_280_pdest;
wire [5:0]   io_diffCommits_info_281_ldest;
wire [7:0]   io_diffCommits_info_281_pdest;
wire [5:0]   io_diffCommits_info_282_ldest;
wire [7:0]   io_diffCommits_info_282_pdest;
wire [5:0]   io_diffCommits_info_283_ldest;
wire [7:0]   io_diffCommits_info_283_pdest;
wire [5:0]   io_diffCommits_info_284_ldest;
wire [7:0]   io_diffCommits_info_284_pdest;
wire [5:0]   io_diffCommits_info_285_ldest;
wire [7:0]   io_diffCommits_info_285_pdest;
wire [5:0]   io_diffCommits_info_286_ldest;
wire [7:0]   io_diffCommits_info_286_pdest;
wire [5:0]   io_diffCommits_info_287_ldest;
wire [7:0]   io_diffCommits_info_287_pdest;
wire [5:0]   io_diffCommits_info_288_ldest;
wire [7:0]   io_diffCommits_info_288_pdest;
wire [5:0]   io_diffCommits_info_289_ldest;
wire [7:0]   io_diffCommits_info_289_pdest;
wire [5:0]   io_diffCommits_info_290_ldest;
wire [7:0]   io_diffCommits_info_290_pdest;
wire [5:0]   io_diffCommits_info_291_ldest;
wire [7:0]   io_diffCommits_info_291_pdest;
wire [5:0]   io_diffCommits_info_292_ldest;
wire [7:0]   io_diffCommits_info_292_pdest;
wire [5:0]   io_diffCommits_info_293_ldest;
wire [7:0]   io_diffCommits_info_293_pdest;
wire [5:0]   io_diffCommits_info_294_ldest;
wire [7:0]   io_diffCommits_info_294_pdest;
wire [5:0]   io_diffCommits_info_295_ldest;
wire [7:0]   io_diffCommits_info_295_pdest;
wire [5:0]   io_diffCommits_info_296_ldest;
wire [7:0]   io_diffCommits_info_296_pdest;
wire [5:0]   io_diffCommits_info_297_ldest;
wire [7:0]   io_diffCommits_info_297_pdest;
wire [5:0]   io_diffCommits_info_298_ldest;
wire [7:0]   io_diffCommits_info_298_pdest;
wire [5:0]   io_diffCommits_info_299_ldest;
wire [7:0]   io_diffCommits_info_299_pdest;
wire [5:0]   io_diffCommits_info_300_ldest;
wire [7:0]   io_diffCommits_info_300_pdest;
wire [5:0]   io_diffCommits_info_301_ldest;
wire [7:0]   io_diffCommits_info_301_pdest;
wire [5:0]   io_diffCommits_info_302_ldest;
wire [7:0]   io_diffCommits_info_302_pdest;
wire [5:0]   io_diffCommits_info_303_ldest;
wire [7:0]   io_diffCommits_info_303_pdest;
wire [5:0]   io_diffCommits_info_304_ldest;
wire [7:0]   io_diffCommits_info_304_pdest;
wire [5:0]   io_diffCommits_info_305_ldest;
wire [7:0]   io_diffCommits_info_305_pdest;
wire [5:0]   io_diffCommits_info_306_ldest;
wire [7:0]   io_diffCommits_info_306_pdest;
wire [5:0]   io_diffCommits_info_307_ldest;
wire [7:0]   io_diffCommits_info_307_pdest;
wire [5:0]   io_diffCommits_info_308_ldest;
wire [7:0]   io_diffCommits_info_308_pdest;
wire [5:0]   io_diffCommits_info_309_ldest;
wire [7:0]   io_diffCommits_info_309_pdest;
wire [5:0]   io_diffCommits_info_310_ldest;
wire [7:0]   io_diffCommits_info_310_pdest;
wire [5:0]   io_diffCommits_info_311_ldest;
wire [7:0]   io_diffCommits_info_311_pdest;
wire [5:0]   io_diffCommits_info_312_ldest;
wire [7:0]   io_diffCommits_info_312_pdest;
wire [5:0]   io_diffCommits_info_313_ldest;
wire [7:0]   io_diffCommits_info_313_pdest;
wire [5:0]   io_diffCommits_info_314_ldest;
wire [7:0]   io_diffCommits_info_314_pdest;
wire [5:0]   io_diffCommits_info_315_ldest;
wire [7:0]   io_diffCommits_info_315_pdest;
wire [5:0]   io_diffCommits_info_316_ldest;
wire [7:0]   io_diffCommits_info_316_pdest;
wire [5:0]   io_diffCommits_info_317_ldest;
wire [7:0]   io_diffCommits_info_317_pdest;
wire [5:0]   io_diffCommits_info_318_ldest;
wire [7:0]   io_diffCommits_info_318_pdest;
wire [5:0]   io_diffCommits_info_319_ldest;
wire [7:0]   io_diffCommits_info_319_pdest;
wire [5:0]   io_diffCommits_info_320_ldest;
wire [7:0]   io_diffCommits_info_320_pdest;
wire [5:0]   io_diffCommits_info_321_ldest;
wire [7:0]   io_diffCommits_info_321_pdest;
wire [5:0]   io_diffCommits_info_322_ldest;
wire [7:0]   io_diffCommits_info_322_pdest;
wire [5:0]   io_diffCommits_info_323_ldest;
wire [7:0]   io_diffCommits_info_323_pdest;
wire [5:0]   io_diffCommits_info_324_ldest;
wire [7:0]   io_diffCommits_info_324_pdest;
wire [5:0]   io_diffCommits_info_325_ldest;
wire [7:0]   io_diffCommits_info_325_pdest;
wire [5:0]   io_diffCommits_info_326_ldest;
wire [7:0]   io_diffCommits_info_326_pdest;
wire [5:0]   io_diffCommits_info_327_ldest;
wire [7:0]   io_diffCommits_info_327_pdest;
wire [5:0]   io_diffCommits_info_328_ldest;
wire [7:0]   io_diffCommits_info_328_pdest;
wire [5:0]   io_diffCommits_info_329_ldest;
wire [7:0]   io_diffCommits_info_329_pdest;
wire [5:0]   io_diffCommits_info_330_ldest;
wire [7:0]   io_diffCommits_info_330_pdest;
wire [5:0]   io_diffCommits_info_331_ldest;
wire [7:0]   io_diffCommits_info_331_pdest;
wire [5:0]   io_diffCommits_info_332_ldest;
wire [7:0]   io_diffCommits_info_332_pdest;
wire [5:0]   io_diffCommits_info_333_ldest;
wire [7:0]   io_diffCommits_info_333_pdest;
wire [5:0]   io_diffCommits_info_334_ldest;
wire [7:0]   io_diffCommits_info_334_pdest;
wire [5:0]   io_diffCommits_info_335_ldest;
wire [7:0]   io_diffCommits_info_335_pdest;
wire [5:0]   io_diffCommits_info_336_ldest;
wire [7:0]   io_diffCommits_info_336_pdest;
wire [5:0]   io_diffCommits_info_337_ldest;
wire [7:0]   io_diffCommits_info_337_pdest;
wire [5:0]   io_diffCommits_info_338_ldest;
wire [7:0]   io_diffCommits_info_338_pdest;
wire [5:0]   io_diffCommits_info_339_ldest;
wire [7:0]   io_diffCommits_info_339_pdest;
wire [5:0]   io_diffCommits_info_340_ldest;
wire [7:0]   io_diffCommits_info_340_pdest;
wire [5:0]   io_diffCommits_info_341_ldest;
wire [7:0]   io_diffCommits_info_341_pdest;
wire [5:0]   io_diffCommits_info_342_ldest;
wire [7:0]   io_diffCommits_info_342_pdest;
wire [5:0]   io_diffCommits_info_343_ldest;
wire [7:0]   io_diffCommits_info_343_pdest;
wire [5:0]   io_diffCommits_info_344_ldest;
wire [7:0]   io_diffCommits_info_344_pdest;
wire [5:0]   io_diffCommits_info_345_ldest;
wire [7:0]   io_diffCommits_info_345_pdest;
wire [5:0]   io_diffCommits_info_346_ldest;
wire [7:0]   io_diffCommits_info_346_pdest;
wire [5:0]   io_diffCommits_info_347_ldest;
wire [7:0]   io_diffCommits_info_347_pdest;
wire [5:0]   io_diffCommits_info_348_ldest;
wire [7:0]   io_diffCommits_info_348_pdest;
wire [5:0]   io_diffCommits_info_349_ldest;
wire [7:0]   io_diffCommits_info_349_pdest;
wire [5:0]   io_diffCommits_info_350_ldest;
wire [7:0]   io_diffCommits_info_350_pdest;
wire [5:0]   io_diffCommits_info_351_ldest;
wire [7:0]   io_diffCommits_info_351_pdest;
wire [5:0]   io_diffCommits_info_352_ldest;
wire [7:0]   io_diffCommits_info_352_pdest;
wire [5:0]   io_diffCommits_info_353_ldest;
wire [7:0]   io_diffCommits_info_353_pdest;
wire [5:0]   io_diffCommits_info_354_ldest;
wire [7:0]   io_diffCommits_info_354_pdest;
wire [5:0]   io_diffCommits_info_355_ldest;
wire [7:0]   io_diffCommits_info_355_pdest;
wire [5:0]   io_diffCommits_info_356_ldest;
wire [7:0]   io_diffCommits_info_356_pdest;
wire [5:0]   io_diffCommits_info_357_ldest;
wire [7:0]   io_diffCommits_info_357_pdest;
wire [5:0]   io_diffCommits_info_358_ldest;
wire [7:0]   io_diffCommits_info_358_pdest;
wire [5:0]   io_diffCommits_info_359_ldest;
wire [7:0]   io_diffCommits_info_359_pdest;
wire [5:0]   io_diffCommits_info_360_ldest;
wire [7:0]   io_diffCommits_info_360_pdest;
wire [5:0]   io_diffCommits_info_361_ldest;
wire [7:0]   io_diffCommits_info_361_pdest;
wire [5:0]   io_diffCommits_info_362_ldest;
wire [7:0]   io_diffCommits_info_362_pdest;
wire [5:0]   io_diffCommits_info_363_ldest;
wire [7:0]   io_diffCommits_info_363_pdest;
wire [5:0]   io_diffCommits_info_364_ldest;
wire [7:0]   io_diffCommits_info_364_pdest;
wire [5:0]   io_diffCommits_info_365_ldest;
wire [7:0]   io_diffCommits_info_365_pdest;
wire [5:0]   io_diffCommits_info_366_ldest;
wire [7:0]   io_diffCommits_info_366_pdest;
wire [5:0]   io_diffCommits_info_367_ldest;
wire [7:0]   io_diffCommits_info_367_pdest;
wire [5:0]   io_diffCommits_info_368_ldest;
wire [7:0]   io_diffCommits_info_368_pdest;
wire [5:0]   io_diffCommits_info_369_ldest;
wire [7:0]   io_diffCommits_info_369_pdest;
wire [5:0]   io_diffCommits_info_370_ldest;
wire [7:0]   io_diffCommits_info_370_pdest;
wire [5:0]   io_diffCommits_info_371_ldest;
wire [7:0]   io_diffCommits_info_371_pdest;
wire [5:0]   io_diffCommits_info_372_ldest;
wire [7:0]   io_diffCommits_info_372_pdest;
wire [5:0]   io_diffCommits_info_373_ldest;
wire [7:0]   io_diffCommits_info_373_pdest;
wire [5:0]   io_diffCommits_info_374_ldest;
wire [7:0]   io_diffCommits_info_374_pdest;
wire [5:0]   io_diffCommits_info_375_ldest;
wire [7:0]   io_diffCommits_info_375_pdest;
wire [5:0]   io_diffCommits_info_376_ldest;
wire [7:0]   io_diffCommits_info_376_pdest;
wire [5:0]   io_diffCommits_info_377_ldest;
wire [7:0]   io_diffCommits_info_377_pdest;
wire [5:0]   io_diffCommits_info_378_ldest;
wire [7:0]   io_diffCommits_info_378_pdest;
wire [5:0]   io_diffCommits_info_379_ldest;
wire [7:0]   io_diffCommits_info_379_pdest;
wire [5:0]   io_diffCommits_info_380_ldest;
wire [7:0]   io_diffCommits_info_380_pdest;
wire [5:0]   io_diffCommits_info_381_ldest;
wire [7:0]   io_diffCommits_info_381_pdest;
wire [5:0]   io_diffCommits_info_382_ldest;
wire [7:0]   io_diffCommits_info_382_pdest;
wire [5:0]   io_diffCommits_info_383_ldest;
wire [7:0]   io_diffCommits_info_383_pdest;
wire [5:0]   io_diffCommits_info_384_ldest;
wire [7:0]   io_diffCommits_info_384_pdest;
wire [5:0]   io_diffCommits_info_385_ldest;
wire [7:0]   io_diffCommits_info_385_pdest;
wire [5:0]   io_diffCommits_info_386_ldest;
wire [7:0]   io_diffCommits_info_386_pdest;
wire [5:0]   io_diffCommits_info_387_ldest;
wire [7:0]   io_diffCommits_info_387_pdest;
wire [5:0]   io_diffCommits_info_388_ldest;
wire [7:0]   io_diffCommits_info_388_pdest;
wire [5:0]   io_diffCommits_info_389_ldest;
wire [7:0]   io_diffCommits_info_389_pdest;
wire [3:0]   io_lsq_scommit        ;
wire         io_lsq_pendingMMIOld  ;
wire         io_lsq_pendingst      ;
wire         io_lsq_pendingPtr_flag;
wire [7:0]   io_lsq_pendingPtr_value;
wire         io_robDeqPtr_flag     ;
wire [7:0]   io_robDeqPtr_value    ;
wire         io_csr_fflags_valid   ;
wire [4:0]   io_csr_fflags_bits    ;
wire         io_csr_vxsat_valid    ;
wire         io_csr_vxsat_bits     ;
wire         io_csr_vstart_valid   ;
wire [63:0]  io_csr_vstart_bits    ;
wire         io_csr_dirty_fs       ;
wire         io_csr_dirty_vs       ;
wire [6:0]   io_csr_perfinfo_retiredInstr;
wire         io_cpu_halt           ;
wire         io_wfi_wfiReq         ;
wire         io_toDecode_isResumeVType;
wire         io_toDecode_walkToArchVType;
wire         io_toDecode_walkVType_valid;
wire         io_toDecode_walkVType_bits_illegal;
wire         io_toDecode_walkVType_bits_vma;
wire         io_toDecode_walkVType_bits_vta;
wire [1:0]   io_toDecode_walkVType_bits_vsew;
wire [2:0]   io_toDecode_walkVType_bits_vlmul;
wire         io_toDecode_commitVType_vtype_valid;
wire         io_toDecode_commitVType_vtype_bits_illegal;
wire         io_toDecode_commitVType_vtype_bits_vma;
wire         io_toDecode_commitVType_vtype_bits_vta;
wire [1:0]   io_toDecode_commitVType_vtype_bits_vsew;
wire [2:0]   io_toDecode_commitVType_vtype_bits_vlmul;
wire         io_toDecode_commitVType_hasVsetvl;
wire         io_readGPAMemAddr_valid;
wire [5:0]   io_readGPAMemAddr_bits_ftqPtr_value;
wire [3:0]   io_readGPAMemAddr_bits_ftqOffset;
wire         io_toVecExcpMod_logicPhyRegMap_0_valid;
wire [5:0]   io_toVecExcpMod_logicPhyRegMap_0_bits_lreg;
wire [6:0]   io_toVecExcpMod_logicPhyRegMap_0_bits_preg;
wire         io_toVecExcpMod_logicPhyRegMap_1_valid;
wire [5:0]   io_toVecExcpMod_logicPhyRegMap_1_bits_lreg;
wire [6:0]   io_toVecExcpMod_logicPhyRegMap_1_bits_preg;
wire         io_toVecExcpMod_logicPhyRegMap_2_valid;
wire [5:0]   io_toVecExcpMod_logicPhyRegMap_2_bits_lreg;
wire [6:0]   io_toVecExcpMod_logicPhyRegMap_2_bits_preg;
wire         io_toVecExcpMod_logicPhyRegMap_3_valid;
wire [5:0]   io_toVecExcpMod_logicPhyRegMap_3_bits_lreg;
wire [6:0]   io_toVecExcpMod_logicPhyRegMap_3_bits_preg;
wire         io_toVecExcpMod_logicPhyRegMap_4_valid;
wire [5:0]   io_toVecExcpMod_logicPhyRegMap_4_bits_lreg;
wire [6:0]   io_toVecExcpMod_logicPhyRegMap_4_bits_preg;
wire         io_toVecExcpMod_logicPhyRegMap_5_valid;
wire [5:0]   io_toVecExcpMod_logicPhyRegMap_5_bits_lreg;
wire [6:0]   io_toVecExcpMod_logicPhyRegMap_5_bits_preg;
wire         io_toVecExcpMod_excpInfo_valid;
wire [6:0]   io_toVecExcpMod_excpInfo_bits_vstart;
wire [1:0]   io_toVecExcpMod_excpInfo_bits_vsew;
wire [1:0]   io_toVecExcpMod_excpInfo_bits_veew;
wire [2:0]   io_toVecExcpMod_excpInfo_bits_vlmul;
wire [2:0]   io_toVecExcpMod_excpInfo_bits_nf;
wire         io_toVecExcpMod_excpInfo_bits_isStride;
wire         io_toVecExcpMod_excpInfo_bits_isIndexed;
wire         io_toVecExcpMod_excpInfo_bits_isWhole;
wire         io_toVecExcpMod_excpInfo_bits_isVlm;
wire [49:0]  io_storeDebugInfo_1_pc;
wire [5:0]   io_perf_0_value       ;
wire [5:0]   io_perf_1_value       ;
wire [5:0]   io_perf_2_value       ;
wire [5:0]   io_perf_3_value       ;
wire [5:0]   io_perf_4_value       ;
wire [5:0]   io_perf_5_value       ;
wire [5:0]   io_perf_6_value       ;
wire [5:0]   io_perf_7_value       ;
wire [5:0]   io_perf_8_value       ;
wire [5:0]   io_perf_9_value       ;
wire [5:0]   io_perf_10_value      ;
wire [5:0]   io_perf_11_value      ;
wire [5:0]   io_perf_12_value      ;
wire [5:0]   io_perf_13_value      ;
wire [5:0]   io_perf_14_value      ;
wire [5:0]   io_perf_15_value      ;
wire [5:0]   io_perf_16_value      ;
wire [5:0]   io_perf_17_value      ;
wire         io_error_0            ;

bosc_Rob U_Rob (
    //clock & reset
    .clock                  ( clk                  ),
    .reset                ( ~tc_if.rst_n          ),
    //rename_in
    // .clock                ( clock                ),
    // .reset                ( reset                ),
    .io_hartId            ( io_hartId            ),
    .io_enq_req_0_valid   ( io_enq_req_0_valid   ),
    .io_enq_req_0_bits_instr ( io_enq_req_0_bits_instr ),
    .io_enq_req_0_bits_pc ( io_enq_req_0_bits_pc ),
    .io_enq_req_0_bits_exceptionVec_0 ( io_enq_req_0_bits_exceptionVec_0 ),
    .io_enq_req_0_bits_exceptionVec_1 ( io_enq_req_0_bits_exceptionVec_1 ),
    .io_enq_req_0_bits_exceptionVec_2 ( io_enq_req_0_bits_exceptionVec_2 ),
    .io_enq_req_0_bits_exceptionVec_3 ( io_enq_req_0_bits_exceptionVec_3 ),
    .io_enq_req_0_bits_exceptionVec_12 ( io_enq_req_0_bits_exceptionVec_12 ),
    .io_enq_req_0_bits_exceptionVec_20 ( io_enq_req_0_bits_exceptionVec_20 ),
    .io_enq_req_0_bits_exceptionVec_22 ( io_enq_req_0_bits_exceptionVec_22 ),
    .io_enq_req_0_bits_isFetchMalAddr ( io_enq_req_0_bits_isFetchMalAddr ),
    .io_enq_req_0_bits_hasException ( io_enq_req_0_bits_hasException ),
    .io_enq_req_0_bits_trigger ( io_enq_req_0_bits_trigger ),
    .io_enq_req_0_bits_preDecodeInfo_isRVC ( io_enq_req_0_bits_preDecodeInfo_isRVC ),
    .io_enq_req_0_bits_crossPageIPFFix ( io_enq_req_0_bits_crossPageIPFFix ),
    .io_enq_req_0_bits_ftqPtr_flag ( io_enq_req_0_bits_ftqPtr_flag ),
    .io_enq_req_0_bits_ftqPtr_value ( io_enq_req_0_bits_ftqPtr_value ),
    .io_enq_req_0_bits_ftqOffset ( io_enq_req_0_bits_ftqOffset ),
    .io_enq_req_0_bits_ldest ( io_enq_req_0_bits_ldest ),
    .io_enq_req_0_bits_fuType ( io_enq_req_0_bits_fuType ),
    .io_enq_req_0_bits_fuOpType ( io_enq_req_0_bits_fuOpType ),
    .io_enq_req_0_bits_rfWen ( io_enq_req_0_bits_rfWen ),
    .io_enq_req_0_bits_fpWen ( io_enq_req_0_bits_fpWen ),
    .io_enq_req_0_bits_vecWen ( io_enq_req_0_bits_vecWen ),
    .io_enq_req_0_bits_v0Wen ( io_enq_req_0_bits_v0Wen ),
    .io_enq_req_0_bits_vlWen ( io_enq_req_0_bits_vlWen ),
    .io_enq_req_0_bits_isXSTrap ( io_enq_req_0_bits_isXSTrap ),
    .io_enq_req_0_bits_waitForward ( io_enq_req_0_bits_waitForward ),
    .io_enq_req_0_bits_blockBackward ( io_enq_req_0_bits_blockBackward ),
    .io_enq_req_0_bits_flushPipe ( io_enq_req_0_bits_flushPipe ),
    .io_enq_req_0_bits_vpu_vill ( io_enq_req_0_bits_vpu_vill ),
    .io_enq_req_0_bits_vpu_vma ( io_enq_req_0_bits_vpu_vma ),
    .io_enq_req_0_bits_vpu_vta ( io_enq_req_0_bits_vpu_vta ),
    .io_enq_req_0_bits_vpu_vsew ( io_enq_req_0_bits_vpu_vsew ),
    .io_enq_req_0_bits_vpu_vlmul ( io_enq_req_0_bits_vpu_vlmul ),
    .io_enq_req_0_bits_vpu_specVill ( io_enq_req_0_bits_vpu_specVill ),
    .io_enq_req_0_bits_vpu_specVma ( io_enq_req_0_bits_vpu_specVma ),
    .io_enq_req_0_bits_vpu_specVta ( io_enq_req_0_bits_vpu_specVta ),
    .io_enq_req_0_bits_vpu_specVsew ( io_enq_req_0_bits_vpu_specVsew ),
    .io_enq_req_0_bits_vpu_specVlmul ( io_enq_req_0_bits_vpu_specVlmul ),
    .io_enq_req_0_bits_vlsInstr ( io_enq_req_0_bits_vlsInstr ),
    .io_enq_req_0_bits_wfflags ( io_enq_req_0_bits_wfflags ),
    .io_enq_req_0_bits_isMove ( io_enq_req_0_bits_isMove ),
    .io_enq_req_0_bits_isVset ( io_enq_req_0_bits_isVset ),
    .io_enq_req_0_bits_firstUop ( io_enq_req_0_bits_firstUop ),
    .io_enq_req_0_bits_lastUop ( io_enq_req_0_bits_lastUop ),
    .io_enq_req_0_bits_numWB ( io_enq_req_0_bits_numWB ),
    .io_enq_req_0_bits_commitType ( io_enq_req_0_bits_commitType ),
    .io_enq_req_0_bits_pdest ( io_enq_req_0_bits_pdest ),
    .io_enq_req_0_bits_robIdx_flag ( io_enq_req_0_bits_robIdx_flag ),
    .io_enq_req_0_bits_robIdx_value ( io_enq_req_0_bits_robIdx_value ),
    .io_enq_req_0_bits_instrSize ( io_enq_req_0_bits_instrSize ),
    .io_enq_req_0_bits_dirtyFs ( io_enq_req_0_bits_dirtyFs ),
    .io_enq_req_0_bits_dirtyVs ( io_enq_req_0_bits_dirtyVs ),
    .io_enq_req_0_bits_traceBlockInPipe_itype ( io_enq_req_0_bits_traceBlockInPipe_itype ),
    .io_enq_req_0_bits_traceBlockInPipe_iretire ( io_enq_req_0_bits_traceBlockInPipe_iretire ),
    .io_enq_req_0_bits_traceBlockInPipe_ilastsize ( io_enq_req_0_bits_traceBlockInPipe_ilastsize ),
    .io_enq_req_0_bits_eliminatedMove ( io_enq_req_0_bits_eliminatedMove ),
    .io_enq_req_0_bits_snapshot ( io_enq_req_0_bits_snapshot ),
    .io_enq_req_0_bits_lqIdx_value ( io_enq_req_0_bits_lqIdx_value ),
    .io_enq_req_0_bits_sqIdx_value ( io_enq_req_0_bits_sqIdx_value ),
    .io_enq_req_0_bits_singleStep ( io_enq_req_0_bits_singleStep ),
    .io_enq_req_0_bits_debug_sim_trig ( io_enq_req_0_bits_debug_sim_trig ),
    .io_enq_req_1_valid   ( io_enq_req_1_valid   ),
    .io_enq_req_1_bits_instr ( io_enq_req_1_bits_instr ),
    .io_enq_req_1_bits_pc ( io_enq_req_1_bits_pc ),
    .io_enq_req_1_bits_exceptionVec_0 ( io_enq_req_1_bits_exceptionVec_0 ),
    .io_enq_req_1_bits_exceptionVec_1 ( io_enq_req_1_bits_exceptionVec_1 ),
    .io_enq_req_1_bits_exceptionVec_2 ( io_enq_req_1_bits_exceptionVec_2 ),
    .io_enq_req_1_bits_exceptionVec_3 ( io_enq_req_1_bits_exceptionVec_3 ),
    .io_enq_req_1_bits_exceptionVec_12 ( io_enq_req_1_bits_exceptionVec_12 ),
    .io_enq_req_1_bits_exceptionVec_20 ( io_enq_req_1_bits_exceptionVec_20 ),
    .io_enq_req_1_bits_exceptionVec_22 ( io_enq_req_1_bits_exceptionVec_22 ),
    .io_enq_req_1_bits_isFetchMalAddr ( io_enq_req_1_bits_isFetchMalAddr ),
    .io_enq_req_1_bits_hasException ( io_enq_req_1_bits_hasException ),
    .io_enq_req_1_bits_trigger ( io_enq_req_1_bits_trigger ),
    .io_enq_req_1_bits_preDecodeInfo_isRVC ( io_enq_req_1_bits_preDecodeInfo_isRVC ),
    .io_enq_req_1_bits_crossPageIPFFix ( io_enq_req_1_bits_crossPageIPFFix ),
    .io_enq_req_1_bits_ftqPtr_flag ( io_enq_req_1_bits_ftqPtr_flag ),
    .io_enq_req_1_bits_ftqPtr_value ( io_enq_req_1_bits_ftqPtr_value ),
    .io_enq_req_1_bits_ftqOffset ( io_enq_req_1_bits_ftqOffset ),
    .io_enq_req_1_bits_ldest ( io_enq_req_1_bits_ldest ),
    .io_enq_req_1_bits_fuType ( io_enq_req_1_bits_fuType ),
    .io_enq_req_1_bits_fuOpType ( io_enq_req_1_bits_fuOpType ),
    .io_enq_req_1_bits_rfWen ( io_enq_req_1_bits_rfWen ),
    .io_enq_req_1_bits_fpWen ( io_enq_req_1_bits_fpWen ),
    .io_enq_req_1_bits_vecWen ( io_enq_req_1_bits_vecWen ),
    .io_enq_req_1_bits_v0Wen ( io_enq_req_1_bits_v0Wen ),
    .io_enq_req_1_bits_vlWen ( io_enq_req_1_bits_vlWen ),
    .io_enq_req_1_bits_isXSTrap ( io_enq_req_1_bits_isXSTrap ),
    .io_enq_req_1_bits_waitForward ( io_enq_req_1_bits_waitForward ),
    .io_enq_req_1_bits_blockBackward ( io_enq_req_1_bits_blockBackward ),
    .io_enq_req_1_bits_flushPipe ( io_enq_req_1_bits_flushPipe ),
    .io_enq_req_1_bits_vpu_vill ( io_enq_req_1_bits_vpu_vill ),
    .io_enq_req_1_bits_vpu_vma ( io_enq_req_1_bits_vpu_vma ),
    .io_enq_req_1_bits_vpu_vta ( io_enq_req_1_bits_vpu_vta ),
    .io_enq_req_1_bits_vpu_vsew ( io_enq_req_1_bits_vpu_vsew ),
    .io_enq_req_1_bits_vpu_vlmul ( io_enq_req_1_bits_vpu_vlmul ),
    .io_enq_req_1_bits_vpu_specVill ( io_enq_req_1_bits_vpu_specVill ),
    .io_enq_req_1_bits_vpu_specVma ( io_enq_req_1_bits_vpu_specVma ),
    .io_enq_req_1_bits_vpu_specVta ( io_enq_req_1_bits_vpu_specVta ),
    .io_enq_req_1_bits_vpu_specVsew ( io_enq_req_1_bits_vpu_specVsew ),
    .io_enq_req_1_bits_vpu_specVlmul ( io_enq_req_1_bits_vpu_specVlmul ),
    .io_enq_req_1_bits_vlsInstr ( io_enq_req_1_bits_vlsInstr ),
    .io_enq_req_1_bits_wfflags ( io_enq_req_1_bits_wfflags ),
    .io_enq_req_1_bits_isMove ( io_enq_req_1_bits_isMove ),
    .io_enq_req_1_bits_isVset ( io_enq_req_1_bits_isVset ),
    .io_enq_req_1_bits_firstUop ( io_enq_req_1_bits_firstUop ),
    .io_enq_req_1_bits_lastUop ( io_enq_req_1_bits_lastUop ),
    .io_enq_req_1_bits_numWB ( io_enq_req_1_bits_numWB ),
    .io_enq_req_1_bits_commitType ( io_enq_req_1_bits_commitType ),
    .io_enq_req_1_bits_pdest ( io_enq_req_1_bits_pdest ),
    .io_enq_req_1_bits_robIdx_flag ( io_enq_req_1_bits_robIdx_flag ),
    .io_enq_req_1_bits_robIdx_value ( io_enq_req_1_bits_robIdx_value ),
    .io_enq_req_1_bits_instrSize ( io_enq_req_1_bits_instrSize ),
    .io_enq_req_1_bits_dirtyFs ( io_enq_req_1_bits_dirtyFs ),
    .io_enq_req_1_bits_dirtyVs ( io_enq_req_1_bits_dirtyVs ),
    .io_enq_req_1_bits_traceBlockInPipe_itype ( io_enq_req_1_bits_traceBlockInPipe_itype ),
    .io_enq_req_1_bits_traceBlockInPipe_iretire ( io_enq_req_1_bits_traceBlockInPipe_iretire ),
    .io_enq_req_1_bits_traceBlockInPipe_ilastsize ( io_enq_req_1_bits_traceBlockInPipe_ilastsize ),
    .io_enq_req_1_bits_eliminatedMove ( io_enq_req_1_bits_eliminatedMove ),
    .io_enq_req_1_bits_snapshot ( io_enq_req_1_bits_snapshot ),
    .io_enq_req_1_bits_lqIdx_value ( io_enq_req_1_bits_lqIdx_value ),
    .io_enq_req_1_bits_sqIdx_value ( io_enq_req_1_bits_sqIdx_value ),
    .io_enq_req_1_bits_singleStep ( io_enq_req_1_bits_singleStep ),
    .io_enq_req_1_bits_debug_sim_trig ( io_enq_req_1_bits_debug_sim_trig ),
    .io_enq_req_2_valid   ( io_enq_req_2_valid   ),
    .io_enq_req_2_bits_instr ( io_enq_req_2_bits_instr ),
    .io_enq_req_2_bits_pc ( io_enq_req_2_bits_pc ),
    .io_enq_req_2_bits_exceptionVec_0 ( io_enq_req_2_bits_exceptionVec_0 ),
    .io_enq_req_2_bits_exceptionVec_1 ( io_enq_req_2_bits_exceptionVec_1 ),
    .io_enq_req_2_bits_exceptionVec_2 ( io_enq_req_2_bits_exceptionVec_2 ),
    .io_enq_req_2_bits_exceptionVec_3 ( io_enq_req_2_bits_exceptionVec_3 ),
    .io_enq_req_2_bits_exceptionVec_12 ( io_enq_req_2_bits_exceptionVec_12 ),
    .io_enq_req_2_bits_exceptionVec_20 ( io_enq_req_2_bits_exceptionVec_20 ),
    .io_enq_req_2_bits_exceptionVec_22 ( io_enq_req_2_bits_exceptionVec_22 ),
    .io_enq_req_2_bits_isFetchMalAddr ( io_enq_req_2_bits_isFetchMalAddr ),
    .io_enq_req_2_bits_hasException ( io_enq_req_2_bits_hasException ),
    .io_enq_req_2_bits_trigger ( io_enq_req_2_bits_trigger ),
    .io_enq_req_2_bits_preDecodeInfo_isRVC ( io_enq_req_2_bits_preDecodeInfo_isRVC ),
    .io_enq_req_2_bits_crossPageIPFFix ( io_enq_req_2_bits_crossPageIPFFix ),
    .io_enq_req_2_bits_ftqPtr_flag ( io_enq_req_2_bits_ftqPtr_flag ),
    .io_enq_req_2_bits_ftqPtr_value ( io_enq_req_2_bits_ftqPtr_value ),
    .io_enq_req_2_bits_ftqOffset ( io_enq_req_2_bits_ftqOffset ),
    .io_enq_req_2_bits_ldest ( io_enq_req_2_bits_ldest ),
    .io_enq_req_2_bits_fuType ( io_enq_req_2_bits_fuType ),
    .io_enq_req_2_bits_fuOpType ( io_enq_req_2_bits_fuOpType ),
    .io_enq_req_2_bits_rfWen ( io_enq_req_2_bits_rfWen ),
    .io_enq_req_2_bits_fpWen ( io_enq_req_2_bits_fpWen ),
    .io_enq_req_2_bits_vecWen ( io_enq_req_2_bits_vecWen ),
    .io_enq_req_2_bits_v0Wen ( io_enq_req_2_bits_v0Wen ),
    .io_enq_req_2_bits_vlWen ( io_enq_req_2_bits_vlWen ),
    .io_enq_req_2_bits_isXSTrap ( io_enq_req_2_bits_isXSTrap ),
    .io_enq_req_2_bits_waitForward ( io_enq_req_2_bits_waitForward ),
    .io_enq_req_2_bits_blockBackward ( io_enq_req_2_bits_blockBackward ),
    .io_enq_req_2_bits_flushPipe ( io_enq_req_2_bits_flushPipe ),
    .io_enq_req_2_bits_vpu_vill ( io_enq_req_2_bits_vpu_vill ),
    .io_enq_req_2_bits_vpu_vma ( io_enq_req_2_bits_vpu_vma ),
    .io_enq_req_2_bits_vpu_vta ( io_enq_req_2_bits_vpu_vta ),
    .io_enq_req_2_bits_vpu_vsew ( io_enq_req_2_bits_vpu_vsew ),
    .io_enq_req_2_bits_vpu_vlmul ( io_enq_req_2_bits_vpu_vlmul ),
    .io_enq_req_2_bits_vpu_specVill ( io_enq_req_2_bits_vpu_specVill ),
    .io_enq_req_2_bits_vpu_specVma ( io_enq_req_2_bits_vpu_specVma ),
    .io_enq_req_2_bits_vpu_specVta ( io_enq_req_2_bits_vpu_specVta ),
    .io_enq_req_2_bits_vpu_specVsew ( io_enq_req_2_bits_vpu_specVsew ),
    .io_enq_req_2_bits_vpu_specVlmul ( io_enq_req_2_bits_vpu_specVlmul ),
    .io_enq_req_2_bits_vlsInstr ( io_enq_req_2_bits_vlsInstr ),
    .io_enq_req_2_bits_wfflags ( io_enq_req_2_bits_wfflags ),
    .io_enq_req_2_bits_isMove ( io_enq_req_2_bits_isMove ),
    .io_enq_req_2_bits_isVset ( io_enq_req_2_bits_isVset ),
    .io_enq_req_2_bits_firstUop ( io_enq_req_2_bits_firstUop ),
    .io_enq_req_2_bits_lastUop ( io_enq_req_2_bits_lastUop ),
    .io_enq_req_2_bits_numWB ( io_enq_req_2_bits_numWB ),
    .io_enq_req_2_bits_commitType ( io_enq_req_2_bits_commitType ),
    .io_enq_req_2_bits_pdest ( io_enq_req_2_bits_pdest ),
    .io_enq_req_2_bits_robIdx_flag ( io_enq_req_2_bits_robIdx_flag ),
    .io_enq_req_2_bits_robIdx_value ( io_enq_req_2_bits_robIdx_value ),
    .io_enq_req_2_bits_instrSize ( io_enq_req_2_bits_instrSize ),
    .io_enq_req_2_bits_dirtyFs ( io_enq_req_2_bits_dirtyFs ),
    .io_enq_req_2_bits_dirtyVs ( io_enq_req_2_bits_dirtyVs ),
    .io_enq_req_2_bits_traceBlockInPipe_itype ( io_enq_req_2_bits_traceBlockInPipe_itype ),
    .io_enq_req_2_bits_traceBlockInPipe_iretire ( io_enq_req_2_bits_traceBlockInPipe_iretire ),
    .io_enq_req_2_bits_traceBlockInPipe_ilastsize ( io_enq_req_2_bits_traceBlockInPipe_ilastsize ),
    .io_enq_req_2_bits_eliminatedMove ( io_enq_req_2_bits_eliminatedMove ),
    .io_enq_req_2_bits_snapshot ( io_enq_req_2_bits_snapshot ),
    .io_enq_req_2_bits_lqIdx_value ( io_enq_req_2_bits_lqIdx_value ),
    .io_enq_req_2_bits_sqIdx_value ( io_enq_req_2_bits_sqIdx_value ),
    .io_enq_req_2_bits_singleStep ( io_enq_req_2_bits_singleStep ),
    .io_enq_req_2_bits_debug_sim_trig ( io_enq_req_2_bits_debug_sim_trig ),
    .io_enq_req_3_valid   ( io_enq_req_3_valid   ),
    .io_enq_req_3_bits_instr ( io_enq_req_3_bits_instr ),
    .io_enq_req_3_bits_pc ( io_enq_req_3_bits_pc ),
    .io_enq_req_3_bits_exceptionVec_0 ( io_enq_req_3_bits_exceptionVec_0 ),
    .io_enq_req_3_bits_exceptionVec_1 ( io_enq_req_3_bits_exceptionVec_1 ),
    .io_enq_req_3_bits_exceptionVec_2 ( io_enq_req_3_bits_exceptionVec_2 ),
    .io_enq_req_3_bits_exceptionVec_3 ( io_enq_req_3_bits_exceptionVec_3 ),
    .io_enq_req_3_bits_exceptionVec_12 ( io_enq_req_3_bits_exceptionVec_12 ),
    .io_enq_req_3_bits_exceptionVec_20 ( io_enq_req_3_bits_exceptionVec_20 ),
    .io_enq_req_3_bits_exceptionVec_22 ( io_enq_req_3_bits_exceptionVec_22 ),
    .io_enq_req_3_bits_isFetchMalAddr ( io_enq_req_3_bits_isFetchMalAddr ),
    .io_enq_req_3_bits_hasException ( io_enq_req_3_bits_hasException ),
    .io_enq_req_3_bits_trigger ( io_enq_req_3_bits_trigger ),
    .io_enq_req_3_bits_preDecodeInfo_isRVC ( io_enq_req_3_bits_preDecodeInfo_isRVC ),
    .io_enq_req_3_bits_crossPageIPFFix ( io_enq_req_3_bits_crossPageIPFFix ),
    .io_enq_req_3_bits_ftqPtr_flag ( io_enq_req_3_bits_ftqPtr_flag ),
    .io_enq_req_3_bits_ftqPtr_value ( io_enq_req_3_bits_ftqPtr_value ),
    .io_enq_req_3_bits_ftqOffset ( io_enq_req_3_bits_ftqOffset ),
    .io_enq_req_3_bits_ldest ( io_enq_req_3_bits_ldest ),
    .io_enq_req_3_bits_fuType ( io_enq_req_3_bits_fuType ),
    .io_enq_req_3_bits_fuOpType ( io_enq_req_3_bits_fuOpType ),
    .io_enq_req_3_bits_rfWen ( io_enq_req_3_bits_rfWen ),
    .io_enq_req_3_bits_fpWen ( io_enq_req_3_bits_fpWen ),
    .io_enq_req_3_bits_vecWen ( io_enq_req_3_bits_vecWen ),
    .io_enq_req_3_bits_v0Wen ( io_enq_req_3_bits_v0Wen ),
    .io_enq_req_3_bits_vlWen ( io_enq_req_3_bits_vlWen ),
    .io_enq_req_3_bits_isXSTrap ( io_enq_req_3_bits_isXSTrap ),
    .io_enq_req_3_bits_waitForward ( io_enq_req_3_bits_waitForward ),
    .io_enq_req_3_bits_blockBackward ( io_enq_req_3_bits_blockBackward ),
    .io_enq_req_3_bits_flushPipe ( io_enq_req_3_bits_flushPipe ),
    .io_enq_req_3_bits_vpu_vill ( io_enq_req_3_bits_vpu_vill ),
    .io_enq_req_3_bits_vpu_vma ( io_enq_req_3_bits_vpu_vma ),
    .io_enq_req_3_bits_vpu_vta ( io_enq_req_3_bits_vpu_vta ),
    .io_enq_req_3_bits_vpu_vsew ( io_enq_req_3_bits_vpu_vsew ),
    .io_enq_req_3_bits_vpu_vlmul ( io_enq_req_3_bits_vpu_vlmul ),
    .io_enq_req_3_bits_vpu_specVill ( io_enq_req_3_bits_vpu_specVill ),
    .io_enq_req_3_bits_vpu_specVma ( io_enq_req_3_bits_vpu_specVma ),
    .io_enq_req_3_bits_vpu_specVta ( io_enq_req_3_bits_vpu_specVta ),
    .io_enq_req_3_bits_vpu_specVsew ( io_enq_req_3_bits_vpu_specVsew ),
    .io_enq_req_3_bits_vpu_specVlmul ( io_enq_req_3_bits_vpu_specVlmul ),
    .io_enq_req_3_bits_vlsInstr ( io_enq_req_3_bits_vlsInstr ),
    .io_enq_req_3_bits_wfflags ( io_enq_req_3_bits_wfflags ),
    .io_enq_req_3_bits_isMove ( io_enq_req_3_bits_isMove ),
    .io_enq_req_3_bits_isVset ( io_enq_req_3_bits_isVset ),
    .io_enq_req_3_bits_firstUop ( io_enq_req_3_bits_firstUop ),
    .io_enq_req_3_bits_lastUop ( io_enq_req_3_bits_lastUop ),
    .io_enq_req_3_bits_numWB ( io_enq_req_3_bits_numWB ),
    .io_enq_req_3_bits_commitType ( io_enq_req_3_bits_commitType ),
    .io_enq_req_3_bits_pdest ( io_enq_req_3_bits_pdest ),
    .io_enq_req_3_bits_robIdx_flag ( io_enq_req_3_bits_robIdx_flag ),
    .io_enq_req_3_bits_robIdx_value ( io_enq_req_3_bits_robIdx_value ),
    .io_enq_req_3_bits_instrSize ( io_enq_req_3_bits_instrSize ),
    .io_enq_req_3_bits_dirtyFs ( io_enq_req_3_bits_dirtyFs ),
    .io_enq_req_3_bits_dirtyVs ( io_enq_req_3_bits_dirtyVs ),
    .io_enq_req_3_bits_traceBlockInPipe_itype ( io_enq_req_3_bits_traceBlockInPipe_itype ),
    .io_enq_req_3_bits_traceBlockInPipe_iretire ( io_enq_req_3_bits_traceBlockInPipe_iretire ),
    .io_enq_req_3_bits_traceBlockInPipe_ilastsize ( io_enq_req_3_bits_traceBlockInPipe_ilastsize ),
    .io_enq_req_3_bits_eliminatedMove ( io_enq_req_3_bits_eliminatedMove ),
    .io_enq_req_3_bits_snapshot ( io_enq_req_3_bits_snapshot ),
    .io_enq_req_3_bits_lqIdx_value ( io_enq_req_3_bits_lqIdx_value ),
    .io_enq_req_3_bits_sqIdx_value ( io_enq_req_3_bits_sqIdx_value ),
    .io_enq_req_3_bits_singleStep ( io_enq_req_3_bits_singleStep ),
    .io_enq_req_3_bits_debug_sim_trig ( io_enq_req_3_bits_debug_sim_trig ),
    .io_enq_req_4_valid   ( io_enq_req_4_valid   ),
    .io_enq_req_4_bits_instr ( io_enq_req_4_bits_instr ),
    .io_enq_req_4_bits_pc ( io_enq_req_4_bits_pc ),
    .io_enq_req_4_bits_exceptionVec_0 ( io_enq_req_4_bits_exceptionVec_0 ),
    .io_enq_req_4_bits_exceptionVec_1 ( io_enq_req_4_bits_exceptionVec_1 ),
    .io_enq_req_4_bits_exceptionVec_2 ( io_enq_req_4_bits_exceptionVec_2 ),
    .io_enq_req_4_bits_exceptionVec_3 ( io_enq_req_4_bits_exceptionVec_3 ),
    .io_enq_req_4_bits_exceptionVec_12 ( io_enq_req_4_bits_exceptionVec_12 ),
    .io_enq_req_4_bits_exceptionVec_20 ( io_enq_req_4_bits_exceptionVec_20 ),
    .io_enq_req_4_bits_exceptionVec_22 ( io_enq_req_4_bits_exceptionVec_22 ),
    .io_enq_req_4_bits_isFetchMalAddr ( io_enq_req_4_bits_isFetchMalAddr ),
    .io_enq_req_4_bits_hasException ( io_enq_req_4_bits_hasException ),
    .io_enq_req_4_bits_trigger ( io_enq_req_4_bits_trigger ),
    .io_enq_req_4_bits_preDecodeInfo_isRVC ( io_enq_req_4_bits_preDecodeInfo_isRVC ),
    .io_enq_req_4_bits_crossPageIPFFix ( io_enq_req_4_bits_crossPageIPFFix ),
    .io_enq_req_4_bits_ftqPtr_flag ( io_enq_req_4_bits_ftqPtr_flag ),
    .io_enq_req_4_bits_ftqPtr_value ( io_enq_req_4_bits_ftqPtr_value ),
    .io_enq_req_4_bits_ftqOffset ( io_enq_req_4_bits_ftqOffset ),
    .io_enq_req_4_bits_ldest ( io_enq_req_4_bits_ldest ),
    .io_enq_req_4_bits_fuType ( io_enq_req_4_bits_fuType ),
    .io_enq_req_4_bits_fuOpType ( io_enq_req_4_bits_fuOpType ),
    .io_enq_req_4_bits_rfWen ( io_enq_req_4_bits_rfWen ),
    .io_enq_req_4_bits_fpWen ( io_enq_req_4_bits_fpWen ),
    .io_enq_req_4_bits_vecWen ( io_enq_req_4_bits_vecWen ),
    .io_enq_req_4_bits_v0Wen ( io_enq_req_4_bits_v0Wen ),
    .io_enq_req_4_bits_vlWen ( io_enq_req_4_bits_vlWen ),
    .io_enq_req_4_bits_isXSTrap ( io_enq_req_4_bits_isXSTrap ),
    .io_enq_req_4_bits_waitForward ( io_enq_req_4_bits_waitForward ),
    .io_enq_req_4_bits_blockBackward ( io_enq_req_4_bits_blockBackward ),
    .io_enq_req_4_bits_flushPipe ( io_enq_req_4_bits_flushPipe ),
    .io_enq_req_4_bits_vpu_vill ( io_enq_req_4_bits_vpu_vill ),
    .io_enq_req_4_bits_vpu_vma ( io_enq_req_4_bits_vpu_vma ),
    .io_enq_req_4_bits_vpu_vta ( io_enq_req_4_bits_vpu_vta ),
    .io_enq_req_4_bits_vpu_vsew ( io_enq_req_4_bits_vpu_vsew ),
    .io_enq_req_4_bits_vpu_vlmul ( io_enq_req_4_bits_vpu_vlmul ),
    .io_enq_req_4_bits_vpu_specVill ( io_enq_req_4_bits_vpu_specVill ),
    .io_enq_req_4_bits_vpu_specVma ( io_enq_req_4_bits_vpu_specVma ),
    .io_enq_req_4_bits_vpu_specVta ( io_enq_req_4_bits_vpu_specVta ),
    .io_enq_req_4_bits_vpu_specVsew ( io_enq_req_4_bits_vpu_specVsew ),
    .io_enq_req_4_bits_vpu_specVlmul ( io_enq_req_4_bits_vpu_specVlmul ),
    .io_enq_req_4_bits_vlsInstr ( io_enq_req_4_bits_vlsInstr ),
    .io_enq_req_4_bits_wfflags ( io_enq_req_4_bits_wfflags ),
    .io_enq_req_4_bits_isMove ( io_enq_req_4_bits_isMove ),
    .io_enq_req_4_bits_isVset ( io_enq_req_4_bits_isVset ),
    .io_enq_req_4_bits_firstUop ( io_enq_req_4_bits_firstUop ),
    .io_enq_req_4_bits_lastUop ( io_enq_req_4_bits_lastUop ),
    .io_enq_req_4_bits_numWB ( io_enq_req_4_bits_numWB ),
    .io_enq_req_4_bits_commitType ( io_enq_req_4_bits_commitType ),
    .io_enq_req_4_bits_pdest ( io_enq_req_4_bits_pdest ),
    .io_enq_req_4_bits_robIdx_flag ( io_enq_req_4_bits_robIdx_flag ),
    .io_enq_req_4_bits_robIdx_value ( io_enq_req_4_bits_robIdx_value ),
    .io_enq_req_4_bits_instrSize ( io_enq_req_4_bits_instrSize ),
    .io_enq_req_4_bits_dirtyFs ( io_enq_req_4_bits_dirtyFs ),
    .io_enq_req_4_bits_dirtyVs ( io_enq_req_4_bits_dirtyVs ),
    .io_enq_req_4_bits_traceBlockInPipe_itype ( io_enq_req_4_bits_traceBlockInPipe_itype ),
    .io_enq_req_4_bits_traceBlockInPipe_iretire ( io_enq_req_4_bits_traceBlockInPipe_iretire ),
    .io_enq_req_4_bits_traceBlockInPipe_ilastsize ( io_enq_req_4_bits_traceBlockInPipe_ilastsize ),
    .io_enq_req_4_bits_eliminatedMove ( io_enq_req_4_bits_eliminatedMove ),
    .io_enq_req_4_bits_snapshot ( io_enq_req_4_bits_snapshot ),
    .io_enq_req_4_bits_lqIdx_value ( io_enq_req_4_bits_lqIdx_value ),
    .io_enq_req_4_bits_sqIdx_value ( io_enq_req_4_bits_sqIdx_value ),
    .io_enq_req_4_bits_singleStep ( io_enq_req_4_bits_singleStep ),
    .io_enq_req_4_bits_debug_sim_trig ( io_enq_req_4_bits_debug_sim_trig ),
    .io_enq_req_5_valid   ( io_enq_req_5_valid   ),
    .io_enq_req_5_bits_instr ( io_enq_req_5_bits_instr ),
    .io_enq_req_5_bits_pc ( io_enq_req_5_bits_pc ),
    .io_enq_req_5_bits_exceptionVec_0 ( io_enq_req_5_bits_exceptionVec_0 ),
    .io_enq_req_5_bits_exceptionVec_1 ( io_enq_req_5_bits_exceptionVec_1 ),
    .io_enq_req_5_bits_exceptionVec_2 ( io_enq_req_5_bits_exceptionVec_2 ),
    .io_enq_req_5_bits_exceptionVec_3 ( io_enq_req_5_bits_exceptionVec_3 ),
    .io_enq_req_5_bits_exceptionVec_12 ( io_enq_req_5_bits_exceptionVec_12 ),
    .io_enq_req_5_bits_exceptionVec_20 ( io_enq_req_5_bits_exceptionVec_20 ),
    .io_enq_req_5_bits_exceptionVec_22 ( io_enq_req_5_bits_exceptionVec_22 ),
    .io_enq_req_5_bits_isFetchMalAddr ( io_enq_req_5_bits_isFetchMalAddr ),
    .io_enq_req_5_bits_hasException ( io_enq_req_5_bits_hasException ),
    .io_enq_req_5_bits_trigger ( io_enq_req_5_bits_trigger ),
    .io_enq_req_5_bits_preDecodeInfo_isRVC ( io_enq_req_5_bits_preDecodeInfo_isRVC ),
    .io_enq_req_5_bits_crossPageIPFFix ( io_enq_req_5_bits_crossPageIPFFix ),
    .io_enq_req_5_bits_ftqPtr_flag ( io_enq_req_5_bits_ftqPtr_flag ),
    .io_enq_req_5_bits_ftqPtr_value ( io_enq_req_5_bits_ftqPtr_value ),
    .io_enq_req_5_bits_ftqOffset ( io_enq_req_5_bits_ftqOffset ),
    .io_enq_req_5_bits_ldest ( io_enq_req_5_bits_ldest ),
    .io_enq_req_5_bits_fuType ( io_enq_req_5_bits_fuType ),
    .io_enq_req_5_bits_fuOpType ( io_enq_req_5_bits_fuOpType ),
    .io_enq_req_5_bits_rfWen ( io_enq_req_5_bits_rfWen ),
    .io_enq_req_5_bits_fpWen ( io_enq_req_5_bits_fpWen ),
    .io_enq_req_5_bits_vecWen ( io_enq_req_5_bits_vecWen ),
    .io_enq_req_5_bits_v0Wen ( io_enq_req_5_bits_v0Wen ),
    .io_enq_req_5_bits_vlWen ( io_enq_req_5_bits_vlWen ),
    .io_enq_req_5_bits_isXSTrap ( io_enq_req_5_bits_isXSTrap ),
    .io_enq_req_5_bits_waitForward ( io_enq_req_5_bits_waitForward ),
    .io_enq_req_5_bits_blockBackward ( io_enq_req_5_bits_blockBackward ),
    .io_enq_req_5_bits_flushPipe ( io_enq_req_5_bits_flushPipe ),
    .io_enq_req_5_bits_vpu_vill ( io_enq_req_5_bits_vpu_vill ),
    .io_enq_req_5_bits_vpu_vma ( io_enq_req_5_bits_vpu_vma ),
    .io_enq_req_5_bits_vpu_vta ( io_enq_req_5_bits_vpu_vta ),
    .io_enq_req_5_bits_vpu_vsew ( io_enq_req_5_bits_vpu_vsew ),
    .io_enq_req_5_bits_vpu_vlmul ( io_enq_req_5_bits_vpu_vlmul ),
    .io_enq_req_5_bits_vpu_specVill ( io_enq_req_5_bits_vpu_specVill ),
    .io_enq_req_5_bits_vpu_specVma ( io_enq_req_5_bits_vpu_specVma ),
    .io_enq_req_5_bits_vpu_specVta ( io_enq_req_5_bits_vpu_specVta ),
    .io_enq_req_5_bits_vpu_specVsew ( io_enq_req_5_bits_vpu_specVsew ),
    .io_enq_req_5_bits_vpu_specVlmul ( io_enq_req_5_bits_vpu_specVlmul ),
    .io_enq_req_5_bits_vlsInstr ( io_enq_req_5_bits_vlsInstr ),
    .io_enq_req_5_bits_wfflags ( io_enq_req_5_bits_wfflags ),
    .io_enq_req_5_bits_isMove ( io_enq_req_5_bits_isMove ),
    .io_enq_req_5_bits_isVset ( io_enq_req_5_bits_isVset ),
    .io_enq_req_5_bits_firstUop ( io_enq_req_5_bits_firstUop ),
    .io_enq_req_5_bits_lastUop ( io_enq_req_5_bits_lastUop ),
    .io_enq_req_5_bits_numWB ( io_enq_req_5_bits_numWB ),
    .io_enq_req_5_bits_commitType ( io_enq_req_5_bits_commitType ),
    .io_enq_req_5_bits_pdest ( io_enq_req_5_bits_pdest ),
    .io_enq_req_5_bits_robIdx_flag ( io_enq_req_5_bits_robIdx_flag ),
    .io_enq_req_5_bits_robIdx_value ( io_enq_req_5_bits_robIdx_value ),
    .io_enq_req_5_bits_instrSize ( io_enq_req_5_bits_instrSize ),
    .io_enq_req_5_bits_dirtyFs ( io_enq_req_5_bits_dirtyFs ),
    .io_enq_req_5_bits_dirtyVs ( io_enq_req_5_bits_dirtyVs ),
    .io_enq_req_5_bits_traceBlockInPipe_itype ( io_enq_req_5_bits_traceBlockInPipe_itype ),
    .io_enq_req_5_bits_traceBlockInPipe_iretire ( io_enq_req_5_bits_traceBlockInPipe_iretire ),
    .io_enq_req_5_bits_traceBlockInPipe_ilastsize ( io_enq_req_5_bits_traceBlockInPipe_ilastsize ),
    .io_enq_req_5_bits_eliminatedMove ( io_enq_req_5_bits_eliminatedMove ),
    .io_enq_req_5_bits_snapshot ( io_enq_req_5_bits_snapshot ),
    .io_enq_req_5_bits_lqIdx_value ( io_enq_req_5_bits_lqIdx_value ),
    .io_enq_req_5_bits_sqIdx_value ( io_enq_req_5_bits_sqIdx_value ),
    .io_enq_req_5_bits_singleStep ( io_enq_req_5_bits_singleStep ),
    .io_enq_req_5_bits_debug_sim_trig ( io_enq_req_5_bits_debug_sim_trig ),
    //WriteBack_in
    .io_writeback_24_valid ( io_writeback_24_valid ),
    .io_writeback_24_bits_data_0 ( io_writeback_24_bits_data_0 ),
    .io_writeback_24_bits_pdest ( io_writeback_24_bits_pdest ),
    .io_writeback_24_bits_robIdx_flag ( io_writeback_24_bits_robIdx_flag ),
    .io_writeback_24_bits_robIdx_value ( io_writeback_24_bits_robIdx_value ),
    .io_writeback_24_bits_vecWen ( io_writeback_24_bits_vecWen ),
    .io_writeback_24_bits_v0Wen ( io_writeback_24_bits_v0Wen ),
    .io_writeback_24_bits_vlWen ( io_writeback_24_bits_vlWen ),
    .io_writeback_24_bits_exceptionVec_0 ( io_writeback_24_bits_exceptionVec_0 ),
    .io_writeback_24_bits_exceptionVec_1 ( io_writeback_24_bits_exceptionVec_1 ),
    .io_writeback_24_bits_exceptionVec_2 ( io_writeback_24_bits_exceptionVec_2 ),
    .io_writeback_24_bits_exceptionVec_3 ( io_writeback_24_bits_exceptionVec_3 ),
    .io_writeback_24_bits_exceptionVec_4 ( io_writeback_24_bits_exceptionVec_4 ),
    .io_writeback_24_bits_exceptionVec_5 ( io_writeback_24_bits_exceptionVec_5 ),
    .io_writeback_24_bits_exceptionVec_6 ( io_writeback_24_bits_exceptionVec_6 ),
    .io_writeback_24_bits_exceptionVec_7 ( io_writeback_24_bits_exceptionVec_7 ),
    .io_writeback_24_bits_exceptionVec_8 ( io_writeback_24_bits_exceptionVec_8 ),
    .io_writeback_24_bits_exceptionVec_9 ( io_writeback_24_bits_exceptionVec_9 ),
    .io_writeback_24_bits_exceptionVec_10 ( io_writeback_24_bits_exceptionVec_10 ),
    .io_writeback_24_bits_exceptionVec_11 ( io_writeback_24_bits_exceptionVec_11 ),
    .io_writeback_24_bits_exceptionVec_12 ( io_writeback_24_bits_exceptionVec_12 ),
    .io_writeback_24_bits_exceptionVec_13 ( io_writeback_24_bits_exceptionVec_13 ),
    .io_writeback_24_bits_exceptionVec_14 ( io_writeback_24_bits_exceptionVec_14 ),
    .io_writeback_24_bits_exceptionVec_15 ( io_writeback_24_bits_exceptionVec_15 ),
    .io_writeback_24_bits_exceptionVec_16 ( io_writeback_24_bits_exceptionVec_16 ),
    .io_writeback_24_bits_exceptionVec_17 ( io_writeback_24_bits_exceptionVec_17 ),
    .io_writeback_24_bits_exceptionVec_18 ( io_writeback_24_bits_exceptionVec_18 ),
    .io_writeback_24_bits_exceptionVec_19 ( io_writeback_24_bits_exceptionVec_19 ),
    .io_writeback_24_bits_exceptionVec_20 ( io_writeback_24_bits_exceptionVec_20 ),
    .io_writeback_24_bits_exceptionVec_21 ( io_writeback_24_bits_exceptionVec_21 ),
    .io_writeback_24_bits_exceptionVec_22 ( io_writeback_24_bits_exceptionVec_22 ),
    .io_writeback_24_bits_exceptionVec_23 ( io_writeback_24_bits_exceptionVec_23 ),
    .io_writeback_24_bits_flushPipe ( io_writeback_24_bits_flushPipe ),
    .io_writeback_24_bits_replay ( io_writeback_24_bits_replay ),
    .io_writeback_24_bits_trigger ( io_writeback_24_bits_trigger ),
    .io_writeback_24_bits_vls_vpu_vill ( io_writeback_24_bits_vls_vpu_vill ),
    .io_writeback_24_bits_vls_vpu_vma ( io_writeback_24_bits_vls_vpu_vma ),
    .io_writeback_24_bits_vls_vpu_vta ( io_writeback_24_bits_vls_vpu_vta ),
    .io_writeback_24_bits_vls_vpu_vsew ( io_writeback_24_bits_vls_vpu_vsew ),
    .io_writeback_24_bits_vls_vpu_vlmul ( io_writeback_24_bits_vls_vpu_vlmul ),
    .io_writeback_24_bits_vls_vpu_specVill ( io_writeback_24_bits_vls_vpu_specVill ),
    .io_writeback_24_bits_vls_vpu_specVma ( io_writeback_24_bits_vls_vpu_specVma ),
    .io_writeback_24_bits_vls_vpu_specVta ( io_writeback_24_bits_vls_vpu_specVta ),
    .io_writeback_24_bits_vls_vpu_specVsew ( io_writeback_24_bits_vls_vpu_specVsew ),
    .io_writeback_24_bits_vls_vpu_specVlmul ( io_writeback_24_bits_vls_vpu_specVlmul ),
    .io_writeback_24_bits_vls_vpu_vm ( io_writeback_24_bits_vls_vpu_vm ),
    .io_writeback_24_bits_vls_vpu_vstart ( io_writeback_24_bits_vls_vpu_vstart ),
    .io_writeback_24_bits_vls_vpu_frm ( io_writeback_24_bits_vls_vpu_frm ),
    .io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst ( io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst ),
    .io_writeback_24_bits_vls_vpu_fpu_isFP32Instr ( io_writeback_24_bits_vls_vpu_fpu_isFP32Instr ),
    .io_writeback_24_bits_vls_vpu_fpu_isFP64Instr ( io_writeback_24_bits_vls_vpu_fpu_isFP64Instr ),
    .io_writeback_24_bits_vls_vpu_fpu_isReduction ( io_writeback_24_bits_vls_vpu_fpu_isReduction ),
    .io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2 ( io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2 ),
    .io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4 ( io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4 ),
    .io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8 ( io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8 ),
    .io_writeback_24_bits_vls_vpu_vxrm ( io_writeback_24_bits_vls_vpu_vxrm ),
    .io_writeback_24_bits_vls_vpu_vuopIdx ( io_writeback_24_bits_vls_vpu_vuopIdx ),
    .io_writeback_24_bits_vls_vpu_lastUop ( io_writeback_24_bits_vls_vpu_lastUop ),
    .io_writeback_24_bits_vls_vpu_vmask ( io_writeback_24_bits_vls_vpu_vmask ),
    .io_writeback_24_bits_vls_vpu_vl ( io_writeback_24_bits_vls_vpu_vl ),
    .io_writeback_24_bits_vls_vpu_nf ( io_writeback_24_bits_vls_vpu_nf ),
    .io_writeback_24_bits_vls_vpu_veew ( io_writeback_24_bits_vls_vpu_veew ),
    .io_writeback_24_bits_vls_vpu_isReverse ( io_writeback_24_bits_vls_vpu_isReverse ),
    .io_writeback_24_bits_vls_vpu_isExt ( io_writeback_24_bits_vls_vpu_isExt ),
    .io_writeback_24_bits_vls_vpu_isNarrow ( io_writeback_24_bits_vls_vpu_isNarrow ),
    .io_writeback_24_bits_vls_vpu_isDstMask ( io_writeback_24_bits_vls_vpu_isDstMask ),
    .io_writeback_24_bits_vls_vpu_isOpMask ( io_writeback_24_bits_vls_vpu_isOpMask ),
    .io_writeback_24_bits_vls_vpu_isMove ( io_writeback_24_bits_vls_vpu_isMove ),
    .io_writeback_24_bits_vls_vpu_isDependOldVd ( io_writeback_24_bits_vls_vpu_isDependOldVd ),
    .io_writeback_24_bits_vls_vpu_isWritePartVd ( io_writeback_24_bits_vls_vpu_isWritePartVd ),
    .io_writeback_24_bits_vls_vpu_isVleff ( io_writeback_24_bits_vls_vpu_isVleff ),
    .io_writeback_24_bits_vls_oldVdPsrc ( io_writeback_24_bits_vls_oldVdPsrc ),
    .io_writeback_24_bits_vls_vdIdx ( io_writeback_24_bits_vls_vdIdx ),
    .io_writeback_24_bits_vls_vdIdxInField ( io_writeback_24_bits_vls_vdIdxInField ),
    .io_writeback_24_bits_vls_isIndexed ( io_writeback_24_bits_vls_isIndexed ),
    .io_writeback_24_bits_vls_isMasked ( io_writeback_24_bits_vls_isMasked ),
    .io_writeback_24_bits_vls_isStrided ( io_writeback_24_bits_vls_isStrided ),
    .io_writeback_24_bits_vls_isWhole ( io_writeback_24_bits_vls_isWhole ),
    .io_writeback_24_bits_vls_isVecLoad ( io_writeback_24_bits_vls_isVecLoad ),
    .io_writeback_24_bits_vls_isVlm ( io_writeback_24_bits_vls_isVlm ),
    .io_writeback_24_bits_debug_isMMIO ( io_writeback_24_bits_debug_isMMIO ),
    .io_writeback_24_bits_debug_isNCIO ( io_writeback_24_bits_debug_isNCIO ),
    .io_writeback_24_bits_debug_isPerfCnt ( io_writeback_24_bits_debug_isPerfCnt ),
    .io_writeback_24_bits_debug_paddr ( io_writeback_24_bits_debug_paddr ),
    .io_writeback_24_bits_debug_vaddr ( io_writeback_24_bits_debug_vaddr ),
    .io_writeback_24_bits_debugInfo_eliminatedMove ( io_writeback_24_bits_debugInfo_eliminatedMove ),
    .io_writeback_24_bits_debugInfo_renameTime ( io_writeback_24_bits_debugInfo_renameTime ),
    .io_writeback_24_bits_debugInfo_dispatchTime ( io_writeback_24_bits_debugInfo_dispatchTime ),
    .io_writeback_24_bits_debugInfo_enqRsTime ( io_writeback_24_bits_debugInfo_enqRsTime ),
    .io_writeback_24_bits_debugInfo_selectTime ( io_writeback_24_bits_debugInfo_selectTime ),
    .io_writeback_24_bits_debugInfo_issueTime ( io_writeback_24_bits_debugInfo_issueTime ),
    .io_writeback_24_bits_debugInfo_writebackTime ( io_writeback_24_bits_debugInfo_writebackTime ),
    .io_writeback_24_bits_debugInfo_runahead_checkpoint_id ( io_writeback_24_bits_debugInfo_runahead_checkpoint_id ),
    .io_writeback_24_bits_debugInfo_tlbFirstReqTime ( io_writeback_24_bits_debugInfo_tlbFirstReqTime ),
    .io_writeback_24_bits_debugInfo_tlbRespTime ( io_writeback_24_bits_debugInfo_tlbRespTime ),
    .io_writeback_24_bits_debug_seqNum ( io_writeback_24_bits_debug_seqNum ),
    .io_writeback_23_valid ( io_writeback_23_valid ),
    .io_writeback_23_bits_data_0 ( io_writeback_23_bits_data_0 ),
    .io_writeback_23_bits_pdest ( io_writeback_23_bits_pdest ),
    .io_writeback_23_bits_robIdx_flag ( io_writeback_23_bits_robIdx_flag ),
    .io_writeback_23_bits_robIdx_value ( io_writeback_23_bits_robIdx_value ),
    .io_writeback_23_bits_vecWen ( io_writeback_23_bits_vecWen ),
    .io_writeback_23_bits_v0Wen ( io_writeback_23_bits_v0Wen ),
    .io_writeback_23_bits_vlWen ( io_writeback_23_bits_vlWen ),
    .io_writeback_23_bits_exceptionVec_0 ( io_writeback_23_bits_exceptionVec_0 ),
    .io_writeback_23_bits_exceptionVec_1 ( io_writeback_23_bits_exceptionVec_1 ),
    .io_writeback_23_bits_exceptionVec_2 ( io_writeback_23_bits_exceptionVec_2 ),
    .io_writeback_23_bits_exceptionVec_3 ( io_writeback_23_bits_exceptionVec_3 ),
    .io_writeback_23_bits_exceptionVec_4 ( io_writeback_23_bits_exceptionVec_4 ),
    .io_writeback_23_bits_exceptionVec_5 ( io_writeback_23_bits_exceptionVec_5 ),
    .io_writeback_23_bits_exceptionVec_6 ( io_writeback_23_bits_exceptionVec_6 ),
    .io_writeback_23_bits_exceptionVec_7 ( io_writeback_23_bits_exceptionVec_7 ),
    .io_writeback_23_bits_exceptionVec_8 ( io_writeback_23_bits_exceptionVec_8 ),
    .io_writeback_23_bits_exceptionVec_9 ( io_writeback_23_bits_exceptionVec_9 ),
    .io_writeback_23_bits_exceptionVec_10 ( io_writeback_23_bits_exceptionVec_10 ),
    .io_writeback_23_bits_exceptionVec_11 ( io_writeback_23_bits_exceptionVec_11 ),
    .io_writeback_23_bits_exceptionVec_12 ( io_writeback_23_bits_exceptionVec_12 ),
    .io_writeback_23_bits_exceptionVec_13 ( io_writeback_23_bits_exceptionVec_13 ),
    .io_writeback_23_bits_exceptionVec_14 ( io_writeback_23_bits_exceptionVec_14 ),
    .io_writeback_23_bits_exceptionVec_15 ( io_writeback_23_bits_exceptionVec_15 ),
    .io_writeback_23_bits_exceptionVec_16 ( io_writeback_23_bits_exceptionVec_16 ),
    .io_writeback_23_bits_exceptionVec_17 ( io_writeback_23_bits_exceptionVec_17 ),
    .io_writeback_23_bits_exceptionVec_18 ( io_writeback_23_bits_exceptionVec_18 ),
    .io_writeback_23_bits_exceptionVec_19 ( io_writeback_23_bits_exceptionVec_19 ),
    .io_writeback_23_bits_exceptionVec_20 ( io_writeback_23_bits_exceptionVec_20 ),
    .io_writeback_23_bits_exceptionVec_21 ( io_writeback_23_bits_exceptionVec_21 ),
    .io_writeback_23_bits_exceptionVec_22 ( io_writeback_23_bits_exceptionVec_22 ),
    .io_writeback_23_bits_exceptionVec_23 ( io_writeback_23_bits_exceptionVec_23 ),
    .io_writeback_23_bits_flushPipe ( io_writeback_23_bits_flushPipe ),
    .io_writeback_23_bits_replay ( io_writeback_23_bits_replay ),
    .io_writeback_23_bits_trigger ( io_writeback_23_bits_trigger ),
    .io_writeback_23_bits_vls_vpu_vill ( io_writeback_23_bits_vls_vpu_vill ),
    .io_writeback_23_bits_vls_vpu_vma ( io_writeback_23_bits_vls_vpu_vma ),
    .io_writeback_23_bits_vls_vpu_vta ( io_writeback_23_bits_vls_vpu_vta ),
    .io_writeback_23_bits_vls_vpu_vsew ( io_writeback_23_bits_vls_vpu_vsew ),
    .io_writeback_23_bits_vls_vpu_vlmul ( io_writeback_23_bits_vls_vpu_vlmul ),
    .io_writeback_23_bits_vls_vpu_specVill ( io_writeback_23_bits_vls_vpu_specVill ),
    .io_writeback_23_bits_vls_vpu_specVma ( io_writeback_23_bits_vls_vpu_specVma ),
    .io_writeback_23_bits_vls_vpu_specVta ( io_writeback_23_bits_vls_vpu_specVta ),
    .io_writeback_23_bits_vls_vpu_specVsew ( io_writeback_23_bits_vls_vpu_specVsew ),
    .io_writeback_23_bits_vls_vpu_specVlmul ( io_writeback_23_bits_vls_vpu_specVlmul ),
    .io_writeback_23_bits_vls_vpu_vm ( io_writeback_23_bits_vls_vpu_vm ),
    .io_writeback_23_bits_vls_vpu_vstart ( io_writeback_23_bits_vls_vpu_vstart ),
    .io_writeback_23_bits_vls_vpu_frm ( io_writeback_23_bits_vls_vpu_frm ),
    .io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst ( io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst ),
    .io_writeback_23_bits_vls_vpu_fpu_isFP32Instr ( io_writeback_23_bits_vls_vpu_fpu_isFP32Instr ),
    .io_writeback_23_bits_vls_vpu_fpu_isFP64Instr ( io_writeback_23_bits_vls_vpu_fpu_isFP64Instr ),
    .io_writeback_23_bits_vls_vpu_fpu_isReduction ( io_writeback_23_bits_vls_vpu_fpu_isReduction ),
    .io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2 ( io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2 ),
    .io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4 ( io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4 ),
    .io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8 ( io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8 ),
    .io_writeback_23_bits_vls_vpu_vxrm ( io_writeback_23_bits_vls_vpu_vxrm ),
    .io_writeback_23_bits_vls_vpu_vuopIdx ( io_writeback_23_bits_vls_vpu_vuopIdx ),
    .io_writeback_23_bits_vls_vpu_lastUop ( io_writeback_23_bits_vls_vpu_lastUop ),
    .io_writeback_23_bits_vls_vpu_vmask ( io_writeback_23_bits_vls_vpu_vmask ),
    .io_writeback_23_bits_vls_vpu_vl ( io_writeback_23_bits_vls_vpu_vl ),
    .io_writeback_23_bits_vls_vpu_nf ( io_writeback_23_bits_vls_vpu_nf ),
    .io_writeback_23_bits_vls_vpu_veew ( io_writeback_23_bits_vls_vpu_veew ),
    .io_writeback_23_bits_vls_vpu_isReverse ( io_writeback_23_bits_vls_vpu_isReverse ),
    .io_writeback_23_bits_vls_vpu_isExt ( io_writeback_23_bits_vls_vpu_isExt ),
    .io_writeback_23_bits_vls_vpu_isNarrow ( io_writeback_23_bits_vls_vpu_isNarrow ),
    .io_writeback_23_bits_vls_vpu_isDstMask ( io_writeback_23_bits_vls_vpu_isDstMask ),
    .io_writeback_23_bits_vls_vpu_isOpMask ( io_writeback_23_bits_vls_vpu_isOpMask ),
    .io_writeback_23_bits_vls_vpu_isMove ( io_writeback_23_bits_vls_vpu_isMove ),
    .io_writeback_23_bits_vls_vpu_isDependOldVd ( io_writeback_23_bits_vls_vpu_isDependOldVd ),
    .io_writeback_23_bits_vls_vpu_isWritePartVd ( io_writeback_23_bits_vls_vpu_isWritePartVd ),
    .io_writeback_23_bits_vls_vpu_isVleff ( io_writeback_23_bits_vls_vpu_isVleff ),
    .io_writeback_23_bits_vls_oldVdPsrc ( io_writeback_23_bits_vls_oldVdPsrc ),
    .io_writeback_23_bits_vls_vdIdx ( io_writeback_23_bits_vls_vdIdx ),
    .io_writeback_23_bits_vls_vdIdxInField ( io_writeback_23_bits_vls_vdIdxInField ),
    .io_writeback_23_bits_vls_isIndexed ( io_writeback_23_bits_vls_isIndexed ),
    .io_writeback_23_bits_vls_isMasked ( io_writeback_23_bits_vls_isMasked ),
    .io_writeback_23_bits_vls_isStrided ( io_writeback_23_bits_vls_isStrided ),
    .io_writeback_23_bits_vls_isWhole ( io_writeback_23_bits_vls_isWhole ),
    .io_writeback_23_bits_vls_isVecLoad ( io_writeback_23_bits_vls_isVecLoad ),
    .io_writeback_23_bits_vls_isVlm ( io_writeback_23_bits_vls_isVlm ),
    .io_writeback_23_bits_debug_isMMIO ( io_writeback_23_bits_debug_isMMIO ),
    .io_writeback_23_bits_debug_isNCIO ( io_writeback_23_bits_debug_isNCIO ),
    .io_writeback_23_bits_debug_isPerfCnt ( io_writeback_23_bits_debug_isPerfCnt ),
    .io_writeback_23_bits_debug_paddr ( io_writeback_23_bits_debug_paddr ),
    .io_writeback_23_bits_debug_vaddr ( io_writeback_23_bits_debug_vaddr ),
    .io_writeback_23_bits_debugInfo_eliminatedMove ( io_writeback_23_bits_debugInfo_eliminatedMove ),
    .io_writeback_23_bits_debugInfo_renameTime ( io_writeback_23_bits_debugInfo_renameTime ),
    .io_writeback_23_bits_debugInfo_dispatchTime ( io_writeback_23_bits_debugInfo_dispatchTime ),
    .io_writeback_23_bits_debugInfo_enqRsTime ( io_writeback_23_bits_debugInfo_enqRsTime ),
    .io_writeback_23_bits_debugInfo_selectTime ( io_writeback_23_bits_debugInfo_selectTime ),
    .io_writeback_23_bits_debugInfo_issueTime ( io_writeback_23_bits_debugInfo_issueTime ),
    .io_writeback_23_bits_debugInfo_writebackTime ( io_writeback_23_bits_debugInfo_writebackTime ),
    .io_writeback_23_bits_debugInfo_runahead_checkpoint_id ( io_writeback_23_bits_debugInfo_runahead_checkpoint_id ),
    .io_writeback_23_bits_debugInfo_tlbFirstReqTime ( io_writeback_23_bits_debugInfo_tlbFirstReqTime ),
    .io_writeback_23_bits_debugInfo_tlbRespTime ( io_writeback_23_bits_debugInfo_tlbRespTime ),
    .io_writeback_23_bits_debug_seqNum ( io_writeback_23_bits_debug_seqNum ),
    .io_writeback_22_valid ( io_writeback_22_valid ),
    .io_writeback_22_bits_data_0 ( io_writeback_22_bits_data_0 ),
    .io_writeback_22_bits_pdest ( io_writeback_22_bits_pdest ),
    .io_writeback_22_bits_robIdx_flag ( io_writeback_22_bits_robIdx_flag ),
    .io_writeback_22_bits_robIdx_value ( io_writeback_22_bits_robIdx_value ),
    .io_writeback_22_bits_intWen ( io_writeback_22_bits_intWen ),
    .io_writeback_22_bits_fpWen ( io_writeback_22_bits_fpWen ),
    .io_writeback_22_bits_exceptionVec_0 ( io_writeback_22_bits_exceptionVec_0 ),
    .io_writeback_22_bits_exceptionVec_1 ( io_writeback_22_bits_exceptionVec_1 ),
    .io_writeback_22_bits_exceptionVec_2 ( io_writeback_22_bits_exceptionVec_2 ),
    .io_writeback_22_bits_exceptionVec_3 ( io_writeback_22_bits_exceptionVec_3 ),
    .io_writeback_22_bits_exceptionVec_4 ( io_writeback_22_bits_exceptionVec_4 ),
    .io_writeback_22_bits_exceptionVec_5 ( io_writeback_22_bits_exceptionVec_5 ),
    .io_writeback_22_bits_exceptionVec_6 ( io_writeback_22_bits_exceptionVec_6 ),
    .io_writeback_22_bits_exceptionVec_7 ( io_writeback_22_bits_exceptionVec_7 ),
    .io_writeback_22_bits_exceptionVec_8 ( io_writeback_22_bits_exceptionVec_8 ),
    .io_writeback_22_bits_exceptionVec_9 ( io_writeback_22_bits_exceptionVec_9 ),
    .io_writeback_22_bits_exceptionVec_10 ( io_writeback_22_bits_exceptionVec_10 ),
    .io_writeback_22_bits_exceptionVec_11 ( io_writeback_22_bits_exceptionVec_11 ),
    .io_writeback_22_bits_exceptionVec_12 ( io_writeback_22_bits_exceptionVec_12 ),
    .io_writeback_22_bits_exceptionVec_13 ( io_writeback_22_bits_exceptionVec_13 ),
    .io_writeback_22_bits_exceptionVec_14 ( io_writeback_22_bits_exceptionVec_14 ),
    .io_writeback_22_bits_exceptionVec_15 ( io_writeback_22_bits_exceptionVec_15 ),
    .io_writeback_22_bits_exceptionVec_16 ( io_writeback_22_bits_exceptionVec_16 ),
    .io_writeback_22_bits_exceptionVec_17 ( io_writeback_22_bits_exceptionVec_17 ),
    .io_writeback_22_bits_exceptionVec_18 ( io_writeback_22_bits_exceptionVec_18 ),
    .io_writeback_22_bits_exceptionVec_19 ( io_writeback_22_bits_exceptionVec_19 ),
    .io_writeback_22_bits_exceptionVec_20 ( io_writeback_22_bits_exceptionVec_20 ),
    .io_writeback_22_bits_exceptionVec_21 ( io_writeback_22_bits_exceptionVec_21 ),
    .io_writeback_22_bits_exceptionVec_22 ( io_writeback_22_bits_exceptionVec_22 ),
    .io_writeback_22_bits_exceptionVec_23 ( io_writeback_22_bits_exceptionVec_23 ),
    .io_writeback_22_bits_flushPipe ( io_writeback_22_bits_flushPipe ),
    .io_writeback_22_bits_replay ( io_writeback_22_bits_replay ),
    .io_writeback_22_bits_lqIdx_flag ( io_writeback_22_bits_lqIdx_flag ),
    .io_writeback_22_bits_lqIdx_value ( io_writeback_22_bits_lqIdx_value ),
    .io_writeback_22_bits_trigger ( io_writeback_22_bits_trigger ),
    .io_writeback_22_bits_predecodeInfo_valid ( io_writeback_22_bits_predecodeInfo_valid ),
    .io_writeback_22_bits_predecodeInfo_isRVC ( io_writeback_22_bits_predecodeInfo_isRVC ),
    .io_writeback_22_bits_predecodeInfo_brType ( io_writeback_22_bits_predecodeInfo_brType ),
    .io_writeback_22_bits_predecodeInfo_isCall ( io_writeback_22_bits_predecodeInfo_isCall ),
    .io_writeback_22_bits_predecodeInfo_isRet ( io_writeback_22_bits_predecodeInfo_isRet ),
    .io_writeback_22_bits_debug_isMMIO ( io_writeback_22_bits_debug_isMMIO ),
    .io_writeback_22_bits_debug_isNCIO ( io_writeback_22_bits_debug_isNCIO ),
    .io_writeback_22_bits_debug_isPerfCnt ( io_writeback_22_bits_debug_isPerfCnt ),
    .io_writeback_22_bits_debug_paddr ( io_writeback_22_bits_debug_paddr ),
    .io_writeback_22_bits_debug_vaddr ( io_writeback_22_bits_debug_vaddr ),
    .io_writeback_22_bits_debugInfo_eliminatedMove ( io_writeback_22_bits_debugInfo_eliminatedMove ),
    .io_writeback_22_bits_debugInfo_renameTime ( io_writeback_22_bits_debugInfo_renameTime ),
    .io_writeback_22_bits_debugInfo_dispatchTime ( io_writeback_22_bits_debugInfo_dispatchTime ),
    .io_writeback_22_bits_debugInfo_enqRsTime ( io_writeback_22_bits_debugInfo_enqRsTime ),
    .io_writeback_22_bits_debugInfo_selectTime ( io_writeback_22_bits_debugInfo_selectTime ),
    .io_writeback_22_bits_debugInfo_issueTime ( io_writeback_22_bits_debugInfo_issueTime ),
    .io_writeback_22_bits_debugInfo_writebackTime ( io_writeback_22_bits_debugInfo_writebackTime ),
    .io_writeback_22_bits_debugInfo_runahead_checkpoint_id ( io_writeback_22_bits_debugInfo_runahead_checkpoint_id ),
    .io_writeback_22_bits_debugInfo_tlbFirstReqTime ( io_writeback_22_bits_debugInfo_tlbFirstReqTime ),
    .io_writeback_22_bits_debugInfo_tlbRespTime ( io_writeback_22_bits_debugInfo_tlbRespTime ),
    .io_writeback_22_bits_debug_seqNum ( io_writeback_22_bits_debug_seqNum ),
    .io_writeback_21_valid ( io_writeback_21_valid ),
    .io_writeback_21_bits_data_0 ( io_writeback_21_bits_data_0 ),
    .io_writeback_21_bits_pdest ( io_writeback_21_bits_pdest ),
    .io_writeback_21_bits_robIdx_flag ( io_writeback_21_bits_robIdx_flag ),
    .io_writeback_21_bits_robIdx_value ( io_writeback_21_bits_robIdx_value ),
    .io_writeback_21_bits_intWen ( io_writeback_21_bits_intWen ),
    .io_writeback_21_bits_fpWen ( io_writeback_21_bits_fpWen ),
    .io_writeback_21_bits_exceptionVec_0 ( io_writeback_21_bits_exceptionVec_0 ),
    .io_writeback_21_bits_exceptionVec_1 ( io_writeback_21_bits_exceptionVec_1 ),
    .io_writeback_21_bits_exceptionVec_2 ( io_writeback_21_bits_exceptionVec_2 ),
    .io_writeback_21_bits_exceptionVec_3 ( io_writeback_21_bits_exceptionVec_3 ),
    .io_writeback_21_bits_exceptionVec_4 ( io_writeback_21_bits_exceptionVec_4 ),
    .io_writeback_21_bits_exceptionVec_5 ( io_writeback_21_bits_exceptionVec_5 ),
    .io_writeback_21_bits_exceptionVec_6 ( io_writeback_21_bits_exceptionVec_6 ),
    .io_writeback_21_bits_exceptionVec_7 ( io_writeback_21_bits_exceptionVec_7 ),
    .io_writeback_21_bits_exceptionVec_8 ( io_writeback_21_bits_exceptionVec_8 ),
    .io_writeback_21_bits_exceptionVec_9 ( io_writeback_21_bits_exceptionVec_9 ),
    .io_writeback_21_bits_exceptionVec_10 ( io_writeback_21_bits_exceptionVec_10 ),
    .io_writeback_21_bits_exceptionVec_11 ( io_writeback_21_bits_exceptionVec_11 ),
    .io_writeback_21_bits_exceptionVec_12 ( io_writeback_21_bits_exceptionVec_12 ),
    .io_writeback_21_bits_exceptionVec_13 ( io_writeback_21_bits_exceptionVec_13 ),
    .io_writeback_21_bits_exceptionVec_14 ( io_writeback_21_bits_exceptionVec_14 ),
    .io_writeback_21_bits_exceptionVec_15 ( io_writeback_21_bits_exceptionVec_15 ),
    .io_writeback_21_bits_exceptionVec_16 ( io_writeback_21_bits_exceptionVec_16 ),
    .io_writeback_21_bits_exceptionVec_17 ( io_writeback_21_bits_exceptionVec_17 ),
    .io_writeback_21_bits_exceptionVec_18 ( io_writeback_21_bits_exceptionVec_18 ),
    .io_writeback_21_bits_exceptionVec_19 ( io_writeback_21_bits_exceptionVec_19 ),
    .io_writeback_21_bits_exceptionVec_20 ( io_writeback_21_bits_exceptionVec_20 ),
    .io_writeback_21_bits_exceptionVec_21 ( io_writeback_21_bits_exceptionVec_21 ),
    .io_writeback_21_bits_exceptionVec_22 ( io_writeback_21_bits_exceptionVec_22 ),
    .io_writeback_21_bits_exceptionVec_23 ( io_writeback_21_bits_exceptionVec_23 ),
    .io_writeback_21_bits_flushPipe ( io_writeback_21_bits_flushPipe ),
    .io_writeback_21_bits_replay ( io_writeback_21_bits_replay ),
    .io_writeback_21_bits_lqIdx_flag ( io_writeback_21_bits_lqIdx_flag ),
    .io_writeback_21_bits_lqIdx_value ( io_writeback_21_bits_lqIdx_value ),
    .io_writeback_21_bits_trigger ( io_writeback_21_bits_trigger ),
    .io_writeback_21_bits_predecodeInfo_valid ( io_writeback_21_bits_predecodeInfo_valid ),
    .io_writeback_21_bits_predecodeInfo_isRVC ( io_writeback_21_bits_predecodeInfo_isRVC ),
    .io_writeback_21_bits_predecodeInfo_brType ( io_writeback_21_bits_predecodeInfo_brType ),
    .io_writeback_21_bits_predecodeInfo_isCall ( io_writeback_21_bits_predecodeInfo_isCall ),
    .io_writeback_21_bits_predecodeInfo_isRet ( io_writeback_21_bits_predecodeInfo_isRet ),
    .io_writeback_21_bits_debug_isMMIO ( io_writeback_21_bits_debug_isMMIO ),
    .io_writeback_21_bits_debug_isNCIO ( io_writeback_21_bits_debug_isNCIO ),
    .io_writeback_21_bits_debug_isPerfCnt ( io_writeback_21_bits_debug_isPerfCnt ),
    .io_writeback_21_bits_debug_paddr ( io_writeback_21_bits_debug_paddr ),
    .io_writeback_21_bits_debug_vaddr ( io_writeback_21_bits_debug_vaddr ),
    .io_writeback_21_bits_debugInfo_eliminatedMove ( io_writeback_21_bits_debugInfo_eliminatedMove ),
    .io_writeback_21_bits_debugInfo_renameTime ( io_writeback_21_bits_debugInfo_renameTime ),
    .io_writeback_21_bits_debugInfo_dispatchTime ( io_writeback_21_bits_debugInfo_dispatchTime ),
    .io_writeback_21_bits_debugInfo_enqRsTime ( io_writeback_21_bits_debugInfo_enqRsTime ),
    .io_writeback_21_bits_debugInfo_selectTime ( io_writeback_21_bits_debugInfo_selectTime ),
    .io_writeback_21_bits_debugInfo_issueTime ( io_writeback_21_bits_debugInfo_issueTime ),
    .io_writeback_21_bits_debugInfo_writebackTime ( io_writeback_21_bits_debugInfo_writebackTime ),
    .io_writeback_21_bits_debugInfo_runahead_checkpoint_id ( io_writeback_21_bits_debugInfo_runahead_checkpoint_id ),
    .io_writeback_21_bits_debugInfo_tlbFirstReqTime ( io_writeback_21_bits_debugInfo_tlbFirstReqTime ),
    .io_writeback_21_bits_debugInfo_tlbRespTime ( io_writeback_21_bits_debugInfo_tlbRespTime ),
    .io_writeback_21_bits_debug_seqNum ( io_writeback_21_bits_debug_seqNum ),
    .io_writeback_20_valid ( io_writeback_20_valid ),
    .io_writeback_20_bits_data_0 ( io_writeback_20_bits_data_0 ),
    .io_writeback_20_bits_pdest ( io_writeback_20_bits_pdest ),
    .io_writeback_20_bits_robIdx_flag ( io_writeback_20_bits_robIdx_flag ),
    .io_writeback_20_bits_robIdx_value ( io_writeback_20_bits_robIdx_value ),
    .io_writeback_20_bits_intWen ( io_writeback_20_bits_intWen ),
    .io_writeback_20_bits_fpWen ( io_writeback_20_bits_fpWen ),
    .io_writeback_20_bits_exceptionVec_0 ( io_writeback_20_bits_exceptionVec_0 ),
    .io_writeback_20_bits_exceptionVec_1 ( io_writeback_20_bits_exceptionVec_1 ),
    .io_writeback_20_bits_exceptionVec_2 ( io_writeback_20_bits_exceptionVec_2 ),
    .io_writeback_20_bits_exceptionVec_3 ( io_writeback_20_bits_exceptionVec_3 ),
    .io_writeback_20_bits_exceptionVec_4 ( io_writeback_20_bits_exceptionVec_4 ),
    .io_writeback_20_bits_exceptionVec_5 ( io_writeback_20_bits_exceptionVec_5 ),
    .io_writeback_20_bits_exceptionVec_6 ( io_writeback_20_bits_exceptionVec_6 ),
    .io_writeback_20_bits_exceptionVec_7 ( io_writeback_20_bits_exceptionVec_7 ),
    .io_writeback_20_bits_exceptionVec_8 ( io_writeback_20_bits_exceptionVec_8 ),
    .io_writeback_20_bits_exceptionVec_9 ( io_writeback_20_bits_exceptionVec_9 ),
    .io_writeback_20_bits_exceptionVec_10 ( io_writeback_20_bits_exceptionVec_10 ),
    .io_writeback_20_bits_exceptionVec_11 ( io_writeback_20_bits_exceptionVec_11 ),
    .io_writeback_20_bits_exceptionVec_12 ( io_writeback_20_bits_exceptionVec_12 ),
    .io_writeback_20_bits_exceptionVec_13 ( io_writeback_20_bits_exceptionVec_13 ),
    .io_writeback_20_bits_exceptionVec_14 ( io_writeback_20_bits_exceptionVec_14 ),
    .io_writeback_20_bits_exceptionVec_15 ( io_writeback_20_bits_exceptionVec_15 ),
    .io_writeback_20_bits_exceptionVec_16 ( io_writeback_20_bits_exceptionVec_16 ),
    .io_writeback_20_bits_exceptionVec_17 ( io_writeback_20_bits_exceptionVec_17 ),
    .io_writeback_20_bits_exceptionVec_18 ( io_writeback_20_bits_exceptionVec_18 ),
    .io_writeback_20_bits_exceptionVec_19 ( io_writeback_20_bits_exceptionVec_19 ),
    .io_writeback_20_bits_exceptionVec_20 ( io_writeback_20_bits_exceptionVec_20 ),
    .io_writeback_20_bits_exceptionVec_21 ( io_writeback_20_bits_exceptionVec_21 ),
    .io_writeback_20_bits_exceptionVec_22 ( io_writeback_20_bits_exceptionVec_22 ),
    .io_writeback_20_bits_exceptionVec_23 ( io_writeback_20_bits_exceptionVec_23 ),
    .io_writeback_20_bits_flushPipe ( io_writeback_20_bits_flushPipe ),
    .io_writeback_20_bits_replay ( io_writeback_20_bits_replay ),
    .io_writeback_20_bits_lqIdx_flag ( io_writeback_20_bits_lqIdx_flag ),
    .io_writeback_20_bits_lqIdx_value ( io_writeback_20_bits_lqIdx_value ),
    .io_writeback_20_bits_trigger ( io_writeback_20_bits_trigger ),
    .io_writeback_20_bits_predecodeInfo_valid ( io_writeback_20_bits_predecodeInfo_valid ),
    .io_writeback_20_bits_predecodeInfo_isRVC ( io_writeback_20_bits_predecodeInfo_isRVC ),
    .io_writeback_20_bits_predecodeInfo_brType ( io_writeback_20_bits_predecodeInfo_brType ),
    .io_writeback_20_bits_predecodeInfo_isCall ( io_writeback_20_bits_predecodeInfo_isCall ),
    .io_writeback_20_bits_predecodeInfo_isRet ( io_writeback_20_bits_predecodeInfo_isRet ),
    .io_writeback_20_bits_debug_isMMIO ( io_writeback_20_bits_debug_isMMIO ),
    .io_writeback_20_bits_debug_isNCIO ( io_writeback_20_bits_debug_isNCIO ),
    .io_writeback_20_bits_debug_isPerfCnt ( io_writeback_20_bits_debug_isPerfCnt ),
    .io_writeback_20_bits_debug_paddr ( io_writeback_20_bits_debug_paddr ),
    .io_writeback_20_bits_debug_vaddr ( io_writeback_20_bits_debug_vaddr ),
    .io_writeback_20_bits_debugInfo_eliminatedMove ( io_writeback_20_bits_debugInfo_eliminatedMove ),
    .io_writeback_20_bits_debugInfo_renameTime ( io_writeback_20_bits_debugInfo_renameTime ),
    .io_writeback_20_bits_debugInfo_dispatchTime ( io_writeback_20_bits_debugInfo_dispatchTime ),
    .io_writeback_20_bits_debugInfo_enqRsTime ( io_writeback_20_bits_debugInfo_enqRsTime ),
    .io_writeback_20_bits_debugInfo_selectTime ( io_writeback_20_bits_debugInfo_selectTime ),
    .io_writeback_20_bits_debugInfo_issueTime ( io_writeback_20_bits_debugInfo_issueTime ),
    .io_writeback_20_bits_debugInfo_writebackTime ( io_writeback_20_bits_debugInfo_writebackTime ),
    .io_writeback_20_bits_debugInfo_runahead_checkpoint_id ( io_writeback_20_bits_debugInfo_runahead_checkpoint_id ),
    .io_writeback_20_bits_debugInfo_tlbFirstReqTime ( io_writeback_20_bits_debugInfo_tlbFirstReqTime ),
    .io_writeback_20_bits_debugInfo_tlbRespTime ( io_writeback_20_bits_debugInfo_tlbRespTime ),
    .io_writeback_20_bits_debug_seqNum ( io_writeback_20_bits_debug_seqNum ),
    .io_writeback_19_valid ( io_writeback_19_valid ),
    .io_writeback_19_bits_data_0 ( io_writeback_19_bits_data_0 ),
    .io_writeback_19_bits_pdest ( io_writeback_19_bits_pdest ),
    .io_writeback_19_bits_robIdx_flag ( io_writeback_19_bits_robIdx_flag ),
    .io_writeback_19_bits_robIdx_value ( io_writeback_19_bits_robIdx_value ),
    .io_writeback_19_bits_intWen ( io_writeback_19_bits_intWen ),
    .io_writeback_19_bits_exceptionVec_0 ( io_writeback_19_bits_exceptionVec_0 ),
    .io_writeback_19_bits_exceptionVec_1 ( io_writeback_19_bits_exceptionVec_1 ),
    .io_writeback_19_bits_exceptionVec_2 ( io_writeback_19_bits_exceptionVec_2 ),
    .io_writeback_19_bits_exceptionVec_3 ( io_writeback_19_bits_exceptionVec_3 ),
    .io_writeback_19_bits_exceptionVec_4 ( io_writeback_19_bits_exceptionVec_4 ),
    .io_writeback_19_bits_exceptionVec_5 ( io_writeback_19_bits_exceptionVec_5 ),
    .io_writeback_19_bits_exceptionVec_6 ( io_writeback_19_bits_exceptionVec_6 ),
    .io_writeback_19_bits_exceptionVec_7 ( io_writeback_19_bits_exceptionVec_7 ),
    .io_writeback_19_bits_exceptionVec_8 ( io_writeback_19_bits_exceptionVec_8 ),
    .io_writeback_19_bits_exceptionVec_9 ( io_writeback_19_bits_exceptionVec_9 ),
    .io_writeback_19_bits_exceptionVec_10 ( io_writeback_19_bits_exceptionVec_10 ),
    .io_writeback_19_bits_exceptionVec_11 ( io_writeback_19_bits_exceptionVec_11 ),
    .io_writeback_19_bits_exceptionVec_12 ( io_writeback_19_bits_exceptionVec_12 ),
    .io_writeback_19_bits_exceptionVec_13 ( io_writeback_19_bits_exceptionVec_13 ),
    .io_writeback_19_bits_exceptionVec_14 ( io_writeback_19_bits_exceptionVec_14 ),
    .io_writeback_19_bits_exceptionVec_15 ( io_writeback_19_bits_exceptionVec_15 ),
    .io_writeback_19_bits_exceptionVec_16 ( io_writeback_19_bits_exceptionVec_16 ),
    .io_writeback_19_bits_exceptionVec_17 ( io_writeback_19_bits_exceptionVec_17 ),
    .io_writeback_19_bits_exceptionVec_18 ( io_writeback_19_bits_exceptionVec_18 ),
    .io_writeback_19_bits_exceptionVec_19 ( io_writeback_19_bits_exceptionVec_19 ),
    .io_writeback_19_bits_exceptionVec_20 ( io_writeback_19_bits_exceptionVec_20 ),
    .io_writeback_19_bits_exceptionVec_21 ( io_writeback_19_bits_exceptionVec_21 ),
    .io_writeback_19_bits_exceptionVec_22 ( io_writeback_19_bits_exceptionVec_22 ),
    .io_writeback_19_bits_exceptionVec_23 ( io_writeback_19_bits_exceptionVec_23 ),
    .io_writeback_19_bits_flushPipe ( io_writeback_19_bits_flushPipe ),
    .io_writeback_19_bits_sqIdx_flag ( io_writeback_19_bits_sqIdx_flag ),
    .io_writeback_19_bits_sqIdx_value ( io_writeback_19_bits_sqIdx_value ),
    .io_writeback_19_bits_trigger ( io_writeback_19_bits_trigger ),
    .io_writeback_19_bits_debug_isMMIO ( io_writeback_19_bits_debug_isMMIO ),
    .io_writeback_19_bits_debug_isNCIO ( io_writeback_19_bits_debug_isNCIO ),
    .io_writeback_19_bits_debug_isPerfCnt ( io_writeback_19_bits_debug_isPerfCnt ),
    .io_writeback_19_bits_debug_paddr ( io_writeback_19_bits_debug_paddr ),
    .io_writeback_19_bits_debug_vaddr ( io_writeback_19_bits_debug_vaddr ),
    .io_writeback_19_bits_debugInfo_eliminatedMove ( io_writeback_19_bits_debugInfo_eliminatedMove ),
    .io_writeback_19_bits_debugInfo_renameTime ( io_writeback_19_bits_debugInfo_renameTime ),
    .io_writeback_19_bits_debugInfo_dispatchTime ( io_writeback_19_bits_debugInfo_dispatchTime ),
    .io_writeback_19_bits_debugInfo_enqRsTime ( io_writeback_19_bits_debugInfo_enqRsTime ),
    .io_writeback_19_bits_debugInfo_selectTime ( io_writeback_19_bits_debugInfo_selectTime ),
    .io_writeback_19_bits_debugInfo_issueTime ( io_writeback_19_bits_debugInfo_issueTime ),
    .io_writeback_19_bits_debugInfo_writebackTime ( io_writeback_19_bits_debugInfo_writebackTime ),
    .io_writeback_19_bits_debugInfo_runahead_checkpoint_id ( io_writeback_19_bits_debugInfo_runahead_checkpoint_id ),
    .io_writeback_19_bits_debugInfo_tlbFirstReqTime ( io_writeback_19_bits_debugInfo_tlbFirstReqTime ),
    .io_writeback_19_bits_debugInfo_tlbRespTime ( io_writeback_19_bits_debugInfo_tlbRespTime ),
    .io_writeback_19_bits_debug_seqNum ( io_writeback_19_bits_debug_seqNum ),
    .io_writeback_18_valid ( io_writeback_18_valid ),
    .io_writeback_18_bits_data_0 ( io_writeback_18_bits_data_0 ),
    .io_writeback_18_bits_pdest ( io_writeback_18_bits_pdest ),
    .io_writeback_18_bits_robIdx_flag ( io_writeback_18_bits_robIdx_flag ),
    .io_writeback_18_bits_robIdx_value ( io_writeback_18_bits_robIdx_value ),
    .io_writeback_18_bits_intWen ( io_writeback_18_bits_intWen ),
    .io_writeback_18_bits_exceptionVec_0 ( io_writeback_18_bits_exceptionVec_0 ),
    .io_writeback_18_bits_exceptionVec_1 ( io_writeback_18_bits_exceptionVec_1 ),
    .io_writeback_18_bits_exceptionVec_2 ( io_writeback_18_bits_exceptionVec_2 ),
    .io_writeback_18_bits_exceptionVec_3 ( io_writeback_18_bits_exceptionVec_3 ),
    .io_writeback_18_bits_exceptionVec_4 ( io_writeback_18_bits_exceptionVec_4 ),
    .io_writeback_18_bits_exceptionVec_5 ( io_writeback_18_bits_exceptionVec_5 ),
    .io_writeback_18_bits_exceptionVec_6 ( io_writeback_18_bits_exceptionVec_6 ),
    .io_writeback_18_bits_exceptionVec_7 ( io_writeback_18_bits_exceptionVec_7 ),
    .io_writeback_18_bits_exceptionVec_8 ( io_writeback_18_bits_exceptionVec_8 ),
    .io_writeback_18_bits_exceptionVec_9 ( io_writeback_18_bits_exceptionVec_9 ),
    .io_writeback_18_bits_exceptionVec_10 ( io_writeback_18_bits_exceptionVec_10 ),
    .io_writeback_18_bits_exceptionVec_11 ( io_writeback_18_bits_exceptionVec_11 ),
    .io_writeback_18_bits_exceptionVec_12 ( io_writeback_18_bits_exceptionVec_12 ),
    .io_writeback_18_bits_exceptionVec_13 ( io_writeback_18_bits_exceptionVec_13 ),
    .io_writeback_18_bits_exceptionVec_14 ( io_writeback_18_bits_exceptionVec_14 ),
    .io_writeback_18_bits_exceptionVec_15 ( io_writeback_18_bits_exceptionVec_15 ),
    .io_writeback_18_bits_exceptionVec_16 ( io_writeback_18_bits_exceptionVec_16 ),
    .io_writeback_18_bits_exceptionVec_17 ( io_writeback_18_bits_exceptionVec_17 ),
    .io_writeback_18_bits_exceptionVec_18 ( io_writeback_18_bits_exceptionVec_18 ),
    .io_writeback_18_bits_exceptionVec_19 ( io_writeback_18_bits_exceptionVec_19 ),
    .io_writeback_18_bits_exceptionVec_20 ( io_writeback_18_bits_exceptionVec_20 ),
    .io_writeback_18_bits_exceptionVec_21 ( io_writeback_18_bits_exceptionVec_21 ),
    .io_writeback_18_bits_exceptionVec_22 ( io_writeback_18_bits_exceptionVec_22 ),
    .io_writeback_18_bits_exceptionVec_23 ( io_writeback_18_bits_exceptionVec_23 ),
    .io_writeback_18_bits_flushPipe ( io_writeback_18_bits_flushPipe ),
    .io_writeback_18_bits_sqIdx_flag ( io_writeback_18_bits_sqIdx_flag ),
    .io_writeback_18_bits_sqIdx_value ( io_writeback_18_bits_sqIdx_value ),
    .io_writeback_18_bits_trigger ( io_writeback_18_bits_trigger ),
    .io_writeback_18_bits_debug_isMMIO ( io_writeback_18_bits_debug_isMMIO ),
    .io_writeback_18_bits_debug_isNCIO ( io_writeback_18_bits_debug_isNCIO ),
    .io_writeback_18_bits_debug_isPerfCnt ( io_writeback_18_bits_debug_isPerfCnt ),
    .io_writeback_18_bits_debug_paddr ( io_writeback_18_bits_debug_paddr ),
    .io_writeback_18_bits_debug_vaddr ( io_writeback_18_bits_debug_vaddr ),
    .io_writeback_18_bits_debugInfo_eliminatedMove ( io_writeback_18_bits_debugInfo_eliminatedMove ),
    .io_writeback_18_bits_debugInfo_renameTime ( io_writeback_18_bits_debugInfo_renameTime ),
    .io_writeback_18_bits_debugInfo_dispatchTime ( io_writeback_18_bits_debugInfo_dispatchTime ),
    .io_writeback_18_bits_debugInfo_enqRsTime ( io_writeback_18_bits_debugInfo_enqRsTime ),
    .io_writeback_18_bits_debugInfo_selectTime ( io_writeback_18_bits_debugInfo_selectTime ),
    .io_writeback_18_bits_debugInfo_issueTime ( io_writeback_18_bits_debugInfo_issueTime ),
    .io_writeback_18_bits_debugInfo_writebackTime ( io_writeback_18_bits_debugInfo_writebackTime ),
    .io_writeback_18_bits_debugInfo_runahead_checkpoint_id ( io_writeback_18_bits_debugInfo_runahead_checkpoint_id ),
    .io_writeback_18_bits_debugInfo_tlbFirstReqTime ( io_writeback_18_bits_debugInfo_tlbFirstReqTime ),
    .io_writeback_18_bits_debugInfo_tlbRespTime ( io_writeback_18_bits_debugInfo_tlbRespTime ),
    .io_writeback_18_bits_debug_seqNum ( io_writeback_18_bits_debug_seqNum ),
    .io_writeback_17_valid ( io_writeback_17_valid ),
    .io_writeback_17_bits_data_0 ( io_writeback_17_bits_data_0 ),
    .io_writeback_17_bits_data_1 ( io_writeback_17_bits_data_1 ),
    .io_writeback_17_bits_data_2 ( io_writeback_17_bits_data_2 ),
    .io_writeback_17_bits_pdest ( io_writeback_17_bits_pdest ),
    .io_writeback_17_bits_robIdx_flag ( io_writeback_17_bits_robIdx_flag ),
    .io_writeback_17_bits_robIdx_value ( io_writeback_17_bits_robIdx_value ),
    .io_writeback_17_bits_vecWen ( io_writeback_17_bits_vecWen ),
    .io_writeback_17_bits_v0Wen ( io_writeback_17_bits_v0Wen ),
    .io_writeback_17_bits_fflags ( io_writeback_17_bits_fflags ),
    .io_writeback_17_bits_wflags ( io_writeback_17_bits_wflags ),
    .io_writeback_17_bits_debugInfo_eliminatedMove ( io_writeback_17_bits_debugInfo_eliminatedMove ),
    .io_writeback_17_bits_debugInfo_renameTime ( io_writeback_17_bits_debugInfo_renameTime ),
    .io_writeback_17_bits_debugInfo_dispatchTime ( io_writeback_17_bits_debugInfo_dispatchTime ),
    .io_writeback_17_bits_debugInfo_enqRsTime ( io_writeback_17_bits_debugInfo_enqRsTime ),
    .io_writeback_17_bits_debugInfo_selectTime ( io_writeback_17_bits_debugInfo_selectTime ),
    .io_writeback_17_bits_debugInfo_issueTime ( io_writeback_17_bits_debugInfo_issueTime ),
    .io_writeback_17_bits_debugInfo_writebackTime ( io_writeback_17_bits_debugInfo_writebackTime ),
    .io_writeback_17_bits_debugInfo_runahead_checkpoint_id ( io_writeback_17_bits_debugInfo_runahead_checkpoint_id ),
    .io_writeback_17_bits_debugInfo_tlbFirstReqTime ( io_writeback_17_bits_debugInfo_tlbFirstReqTime ),
    .io_writeback_17_bits_debugInfo_tlbRespTime ( io_writeback_17_bits_debugInfo_tlbRespTime ),
    .io_writeback_17_bits_debug_seqNum ( io_writeback_17_bits_debug_seqNum ),
    .io_writeback_16_valid ( io_writeback_16_valid ),
    .io_writeback_16_bits_data_0 ( io_writeback_16_bits_data_0 ),
    .io_writeback_16_bits_data_1 ( io_writeback_16_bits_data_1 ),
    .io_writeback_16_bits_data_2 ( io_writeback_16_bits_data_2 ),
    .io_writeback_16_bits_data_3 ( io_writeback_16_bits_data_3 ),
    .io_writeback_16_bits_pdest ( io_writeback_16_bits_pdest ),
    .io_writeback_16_bits_robIdx_flag ( io_writeback_16_bits_robIdx_flag ),
    .io_writeback_16_bits_robIdx_value ( io_writeback_16_bits_robIdx_value ),
    .io_writeback_16_bits_fpWen ( io_writeback_16_bits_fpWen ),
    .io_writeback_16_bits_vecWen ( io_writeback_16_bits_vecWen ),
    .io_writeback_16_bits_v0Wen ( io_writeback_16_bits_v0Wen ),
    .io_writeback_16_bits_fflags ( io_writeback_16_bits_fflags ),
    .io_writeback_16_bits_wflags ( io_writeback_16_bits_wflags ),
    .io_writeback_16_bits_debugInfo_eliminatedMove ( io_writeback_16_bits_debugInfo_eliminatedMove ),
    .io_writeback_16_bits_debugInfo_renameTime ( io_writeback_16_bits_debugInfo_renameTime ),
    .io_writeback_16_bits_debugInfo_dispatchTime ( io_writeback_16_bits_debugInfo_dispatchTime ),
    .io_writeback_16_bits_debugInfo_enqRsTime ( io_writeback_16_bits_debugInfo_enqRsTime ),
    .io_writeback_16_bits_debugInfo_selectTime ( io_writeback_16_bits_debugInfo_selectTime ),
    .io_writeback_16_bits_debugInfo_issueTime ( io_writeback_16_bits_debugInfo_issueTime ),
    .io_writeback_16_bits_debugInfo_writebackTime ( io_writeback_16_bits_debugInfo_writebackTime ),
    .io_writeback_16_bits_debugInfo_runahead_checkpoint_id ( io_writeback_16_bits_debugInfo_runahead_checkpoint_id ),
    .io_writeback_16_bits_debugInfo_tlbFirstReqTime ( io_writeback_16_bits_debugInfo_tlbFirstReqTime ),
    .io_writeback_16_bits_debugInfo_tlbRespTime ( io_writeback_16_bits_debugInfo_tlbRespTime ),
    .io_writeback_16_bits_debug_seqNum ( io_writeback_16_bits_debug_seqNum ),
    .io_writeback_15_valid ( io_writeback_15_valid ),
    .io_writeback_15_bits_data_0 ( io_writeback_15_bits_data_0 ),
    .io_writeback_15_bits_data_1 ( io_writeback_15_bits_data_1 ),
    .io_writeback_15_bits_data_2 ( io_writeback_15_bits_data_2 ),
    .io_writeback_15_bits_pdest ( io_writeback_15_bits_pdest ),
    .io_writeback_15_bits_robIdx_flag ( io_writeback_15_bits_robIdx_flag ),
    .io_writeback_15_bits_robIdx_value ( io_writeback_15_bits_robIdx_value ),
    .io_writeback_15_bits_vecWen ( io_writeback_15_bits_vecWen ),
    .io_writeback_15_bits_v0Wen ( io_writeback_15_bits_v0Wen ),
    .io_writeback_15_bits_fflags ( io_writeback_15_bits_fflags ),
    .io_writeback_15_bits_wflags ( io_writeback_15_bits_wflags ),
    .io_writeback_15_bits_vxsat ( io_writeback_15_bits_vxsat ),
    .io_writeback_15_bits_debugInfo_eliminatedMove ( io_writeback_15_bits_debugInfo_eliminatedMove ),
    .io_writeback_15_bits_debugInfo_renameTime ( io_writeback_15_bits_debugInfo_renameTime ),
    .io_writeback_15_bits_debugInfo_dispatchTime ( io_writeback_15_bits_debugInfo_dispatchTime ),
    .io_writeback_15_bits_debugInfo_enqRsTime ( io_writeback_15_bits_debugInfo_enqRsTime ),
    .io_writeback_15_bits_debugInfo_selectTime ( io_writeback_15_bits_debugInfo_selectTime ),
    .io_writeback_15_bits_debugInfo_issueTime ( io_writeback_15_bits_debugInfo_issueTime ),
    .io_writeback_15_bits_debugInfo_writebackTime ( io_writeback_15_bits_debugInfo_writebackTime ),
    .io_writeback_15_bits_debugInfo_runahead_checkpoint_id ( io_writeback_15_bits_debugInfo_runahead_checkpoint_id ),
    .io_writeback_15_bits_debugInfo_tlbFirstReqTime ( io_writeback_15_bits_debugInfo_tlbFirstReqTime ),
    .io_writeback_15_bits_debugInfo_tlbRespTime ( io_writeback_15_bits_debugInfo_tlbRespTime ),
    .io_writeback_15_bits_debug_seqNum ( io_writeback_15_bits_debug_seqNum ),
    .io_writeback_14_valid ( io_writeback_14_valid ),
    .io_writeback_14_bits_data_0 ( io_writeback_14_bits_data_0 ),
    .io_writeback_14_bits_data_1 ( io_writeback_14_bits_data_1 ),
    .io_writeback_14_bits_data_2 ( io_writeback_14_bits_data_2 ),
    .io_writeback_14_bits_data_3 ( io_writeback_14_bits_data_3 ),
    .io_writeback_14_bits_data_4 ( io_writeback_14_bits_data_4 ),
    .io_writeback_14_bits_data_5 ( io_writeback_14_bits_data_5 ),
    .io_writeback_14_bits_pdest ( io_writeback_14_bits_pdest ),
    .io_writeback_14_bits_robIdx_flag ( io_writeback_14_bits_robIdx_flag ),
    .io_writeback_14_bits_robIdx_value ( io_writeback_14_bits_robIdx_value ),
    .io_writeback_14_bits_intWen ( io_writeback_14_bits_intWen ),
    .io_writeback_14_bits_fpWen ( io_writeback_14_bits_fpWen ),
    .io_writeback_14_bits_vecWen ( io_writeback_14_bits_vecWen ),
    .io_writeback_14_bits_v0Wen ( io_writeback_14_bits_v0Wen ),
    .io_writeback_14_bits_vlWen ( io_writeback_14_bits_vlWen ),
    .io_writeback_14_bits_fflags ( io_writeback_14_bits_fflags ),
    .io_writeback_14_bits_wflags ( io_writeback_14_bits_wflags ),
    .io_writeback_14_bits_exceptionVec_2 ( io_writeback_14_bits_exceptionVec_2 ),
    .io_writeback_14_bits_debugInfo_eliminatedMove ( io_writeback_14_bits_debugInfo_eliminatedMove ),
    .io_writeback_14_bits_debugInfo_renameTime ( io_writeback_14_bits_debugInfo_renameTime ),
    .io_writeback_14_bits_debugInfo_dispatchTime ( io_writeback_14_bits_debugInfo_dispatchTime ),
    .io_writeback_14_bits_debugInfo_enqRsTime ( io_writeback_14_bits_debugInfo_enqRsTime ),
    .io_writeback_14_bits_debugInfo_selectTime ( io_writeback_14_bits_debugInfo_selectTime ),
    .io_writeback_14_bits_debugInfo_issueTime ( io_writeback_14_bits_debugInfo_issueTime ),
    .io_writeback_14_bits_debugInfo_writebackTime ( io_writeback_14_bits_debugInfo_writebackTime ),
    .io_writeback_14_bits_debugInfo_runahead_checkpoint_id ( io_writeback_14_bits_debugInfo_runahead_checkpoint_id ),
    .io_writeback_14_bits_debugInfo_tlbFirstReqTime ( io_writeback_14_bits_debugInfo_tlbFirstReqTime ),
    .io_writeback_14_bits_debugInfo_tlbRespTime ( io_writeback_14_bits_debugInfo_tlbRespTime ),
    .io_writeback_14_bits_debug_seqNum ( io_writeback_14_bits_debug_seqNum ),
    .io_writeback_13_valid ( io_writeback_13_valid ),
    .io_writeback_13_bits_data_0 ( io_writeback_13_bits_data_0 ),
    .io_writeback_13_bits_data_1 ( io_writeback_13_bits_data_1 ),
    .io_writeback_13_bits_data_2 ( io_writeback_13_bits_data_2 ),
    .io_writeback_13_bits_pdest ( io_writeback_13_bits_pdest ),
    .io_writeback_13_bits_robIdx_flag ( io_writeback_13_bits_robIdx_flag ),
    .io_writeback_13_bits_robIdx_value ( io_writeback_13_bits_robIdx_value ),
    .io_writeback_13_bits_vecWen ( io_writeback_13_bits_vecWen ),
    .io_writeback_13_bits_v0Wen ( io_writeback_13_bits_v0Wen ),
    .io_writeback_13_bits_fflags ( io_writeback_13_bits_fflags ),
    .io_writeback_13_bits_wflags ( io_writeback_13_bits_wflags ),
    .io_writeback_13_bits_vxsat ( io_writeback_13_bits_vxsat ),
    .io_writeback_13_bits_exceptionVec_2 ( io_writeback_13_bits_exceptionVec_2 ),
    .io_writeback_13_bits_debugInfo_eliminatedMove ( io_writeback_13_bits_debugInfo_eliminatedMove ),
    .io_writeback_13_bits_debugInfo_renameTime ( io_writeback_13_bits_debugInfo_renameTime ),
    .io_writeback_13_bits_debugInfo_dispatchTime ( io_writeback_13_bits_debugInfo_dispatchTime ),
    .io_writeback_13_bits_debugInfo_enqRsTime ( io_writeback_13_bits_debugInfo_enqRsTime ),
    .io_writeback_13_bits_debugInfo_selectTime ( io_writeback_13_bits_debugInfo_selectTime ),
    .io_writeback_13_bits_debugInfo_issueTime ( io_writeback_13_bits_debugInfo_issueTime ),
    .io_writeback_13_bits_debugInfo_writebackTime ( io_writeback_13_bits_debugInfo_writebackTime ),
    .io_writeback_13_bits_debugInfo_runahead_checkpoint_id ( io_writeback_13_bits_debugInfo_runahead_checkpoint_id ),
    .io_writeback_13_bits_debugInfo_tlbFirstReqTime ( io_writeback_13_bits_debugInfo_tlbFirstReqTime ),
    .io_writeback_13_bits_debugInfo_tlbRespTime ( io_writeback_13_bits_debugInfo_tlbRespTime ),
    .io_writeback_13_bits_debug_seqNum ( io_writeback_13_bits_debug_seqNum ),
    .io_writeback_7_valid ( io_writeback_7_valid ),
    .io_writeback_7_bits_data_0 ( io_writeback_7_bits_data_0 ),
    .io_writeback_7_bits_data_1 ( io_writeback_7_bits_data_1 ),
    .io_writeback_7_bits_pdest ( io_writeback_7_bits_pdest ),
    .io_writeback_7_bits_robIdx_flag ( io_writeback_7_bits_robIdx_flag ),
    .io_writeback_7_bits_robIdx_value ( io_writeback_7_bits_robIdx_value ),
    .io_writeback_7_bits_intWen ( io_writeback_7_bits_intWen ),
    .io_writeback_7_bits_redirect_valid ( io_writeback_7_bits_redirect_valid ),
    .io_writeback_7_bits_redirect_bits_isRVC ( io_writeback_7_bits_redirect_bits_isRVC ),
    .io_writeback_7_bits_redirect_bits_robIdx_flag ( io_writeback_7_bits_redirect_bits_robIdx_flag ),
    .io_writeback_7_bits_redirect_bits_robIdx_value ( io_writeback_7_bits_redirect_bits_robIdx_value ),
    .io_writeback_7_bits_redirect_bits_ftqIdx_flag ( io_writeback_7_bits_redirect_bits_ftqIdx_flag ),
    .io_writeback_7_bits_redirect_bits_ftqIdx_value ( io_writeback_7_bits_redirect_bits_ftqIdx_value ),
    .io_writeback_7_bits_redirect_bits_ftqOffset ( io_writeback_7_bits_redirect_bits_ftqOffset ),
    .io_writeback_7_bits_redirect_bits_level ( io_writeback_7_bits_redirect_bits_level ),
    .io_writeback_7_bits_redirect_bits_interrupt ( io_writeback_7_bits_redirect_bits_interrupt ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_pc ( io_writeback_7_bits_redirect_bits_cfiUpdate_pc ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid ( io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC ( io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType ( io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall ( io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet ( io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_ssp ( io_writeback_7_bits_redirect_bits_cfiUpdate_ssp ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_sctr ( io_writeback_7_bits_redirect_bits_cfiUpdate_sctr ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag ( io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value ( io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag ( io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value ( io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag ( io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value ( io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr ( io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist ( io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist ( io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist ( io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist ( io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist ( io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist ( io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist ( io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist ( io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist ( io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist ( io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist ( io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist ( io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist ( io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist ( io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist ( io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist ( io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist ( io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist ( io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0 ( io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0 ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1 ( io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1 ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2 ( io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2 ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3 ( io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3 ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0 ( io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0 ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1 ( io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1 ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2 ( io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2 ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3 ( io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3 ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0 ( io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0 ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1 ( io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1 ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2 ( io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2 ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3 ( io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3 ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0 ( io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0 ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1 ( io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1 ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2 ( io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2 ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3 ( io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3 ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0 ( io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0 ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1 ( io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1 ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2 ( io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2 ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3 ( io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3 ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0 ( io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0 ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1 ( io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1 ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2 ( io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2 ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3 ( io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3 ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH ( io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_ghr ( io_writeback_7_bits_redirect_bits_cfiUpdate_ghr ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag ( io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value ( io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0 ( io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0 ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1 ( io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1 ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit ( io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit ( io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit ( io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken ( io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_target ( io_writeback_7_bits_redirect_bits_cfiUpdate_target ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_taken ( io_writeback_7_bits_redirect_bits_cfiUpdate_taken ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred ( io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_shift ( io_writeback_7_bits_redirect_bits_cfiUpdate_shift ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist ( io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF ( io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF ( io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF ),
    .io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF ( io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF ),
    .io_writeback_7_bits_redirect_bits_fullTarget ( io_writeback_7_bits_redirect_bits_fullTarget ),
    .io_writeback_7_bits_redirect_bits_stFtqIdx_flag ( io_writeback_7_bits_redirect_bits_stFtqIdx_flag ),
    .io_writeback_7_bits_redirect_bits_stFtqIdx_value ( io_writeback_7_bits_redirect_bits_stFtqIdx_value ),
    .io_writeback_7_bits_redirect_bits_stFtqOffset ( io_writeback_7_bits_redirect_bits_stFtqOffset ),
    .io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id ( io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id ),
    .io_writeback_7_bits_redirect_bits_debugIsCtrl ( io_writeback_7_bits_redirect_bits_debugIsCtrl ),
    .io_writeback_7_bits_redirect_bits_debugIsMemVio ( io_writeback_7_bits_redirect_bits_debugIsMemVio ),
    .io_writeback_7_bits_exceptionVec_2 ( io_writeback_7_bits_exceptionVec_2 ),
    .io_writeback_7_bits_exceptionVec_3 ( io_writeback_7_bits_exceptionVec_3 ),
    .io_writeback_7_bits_exceptionVec_8 ( io_writeback_7_bits_exceptionVec_8 ),
    .io_writeback_7_bits_exceptionVec_9 ( io_writeback_7_bits_exceptionVec_9 ),
    .io_writeback_7_bits_exceptionVec_10 ( io_writeback_7_bits_exceptionVec_10 ),
    .io_writeback_7_bits_exceptionVec_11 ( io_writeback_7_bits_exceptionVec_11 ),
    .io_writeback_7_bits_exceptionVec_22 ( io_writeback_7_bits_exceptionVec_22 ),
    .io_writeback_7_bits_flushPipe ( io_writeback_7_bits_flushPipe ),
    .io_writeback_7_bits_predecodeInfo_valid ( io_writeback_7_bits_predecodeInfo_valid ),
    .io_writeback_7_bits_predecodeInfo_isRVC ( io_writeback_7_bits_predecodeInfo_isRVC ),
    .io_writeback_7_bits_predecodeInfo_brType ( io_writeback_7_bits_predecodeInfo_brType ),
    .io_writeback_7_bits_predecodeInfo_isCall ( io_writeback_7_bits_predecodeInfo_isCall ),
    .io_writeback_7_bits_predecodeInfo_isRet ( io_writeback_7_bits_predecodeInfo_isRet ),
    .io_writeback_7_bits_debug_isPerfCnt ( io_writeback_7_bits_debug_isPerfCnt ),
    .io_writeback_7_bits_debugInfo_eliminatedMove ( io_writeback_7_bits_debugInfo_eliminatedMove ),
    .io_writeback_7_bits_debugInfo_renameTime ( io_writeback_7_bits_debugInfo_renameTime ),
    .io_writeback_7_bits_debugInfo_dispatchTime ( io_writeback_7_bits_debugInfo_dispatchTime ),
    .io_writeback_7_bits_debugInfo_enqRsTime ( io_writeback_7_bits_debugInfo_enqRsTime ),
    .io_writeback_7_bits_debugInfo_selectTime ( io_writeback_7_bits_debugInfo_selectTime ),
    .io_writeback_7_bits_debugInfo_issueTime ( io_writeback_7_bits_debugInfo_issueTime ),
    .io_writeback_7_bits_debugInfo_writebackTime ( io_writeback_7_bits_debugInfo_writebackTime ),
    .io_writeback_7_bits_debugInfo_runahead_checkpoint_id ( io_writeback_7_bits_debugInfo_runahead_checkpoint_id ),
    .io_writeback_7_bits_debugInfo_tlbFirstReqTime ( io_writeback_7_bits_debugInfo_tlbFirstReqTime ),
    .io_writeback_7_bits_debugInfo_tlbRespTime ( io_writeback_7_bits_debugInfo_tlbRespTime ),
    .io_writeback_7_bits_debug_seqNum ( io_writeback_7_bits_debug_seqNum ),
    .io_writeback_5_valid ( io_writeback_5_valid ),
    .io_writeback_5_bits_redirect_valid ( io_writeback_5_bits_redirect_valid ),
    .io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred ( io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred ),
    .io_writeback_3_valid ( io_writeback_3_valid ),
    .io_writeback_3_bits_redirect_valid ( io_writeback_3_bits_redirect_valid ),
    .io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred ( io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred ),
    .io_writeback_1_valid ( io_writeback_1_valid ),
    .io_writeback_1_bits_redirect_valid ( io_writeback_1_bits_redirect_valid ),
    .io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred ( io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred ),
    .io_exuWriteback_26_valid ( io_exuWriteback_26_valid ),
    .io_exuWriteback_26_bits_robIdx_value ( io_exuWriteback_26_bits_robIdx_value ),
    .io_exuWriteback_25_valid ( io_exuWriteback_25_valid ),
    .io_exuWriteback_25_bits_robIdx_value ( io_exuWriteback_25_bits_robIdx_value ),
    .io_exuWriteback_24_valid ( io_exuWriteback_24_valid ),
    .io_exuWriteback_24_bits_data_0 ( io_exuWriteback_24_bits_data_0 ),
    .io_exuWriteback_24_bits_pdest ( io_exuWriteback_24_bits_pdest ),
    .io_exuWriteback_24_bits_robIdx_value ( io_exuWriteback_24_bits_robIdx_value ),
    .io_exuWriteback_24_bits_vecWen ( io_exuWriteback_24_bits_vecWen ),
    .io_exuWriteback_24_bits_v0Wen ( io_exuWriteback_24_bits_v0Wen ),
    .io_exuWriteback_24_bits_vls_vdIdx ( io_exuWriteback_24_bits_vls_vdIdx ),
    .io_exuWriteback_24_bits_debug_isMMIO ( io_exuWriteback_24_bits_debug_isMMIO ),
    .io_exuWriteback_24_bits_debug_isNCIO ( io_exuWriteback_24_bits_debug_isNCIO ),
    .io_exuWriteback_24_bits_debug_isPerfCnt ( io_exuWriteback_24_bits_debug_isPerfCnt ),
    .io_exuWriteback_24_bits_debug_paddr ( io_exuWriteback_24_bits_debug_paddr ),
    .io_exuWriteback_23_valid ( io_exuWriteback_23_valid ),
    .io_exuWriteback_23_bits_data_0 ( io_exuWriteback_23_bits_data_0 ),
    .io_exuWriteback_23_bits_pdest ( io_exuWriteback_23_bits_pdest ),
    .io_exuWriteback_23_bits_robIdx_value ( io_exuWriteback_23_bits_robIdx_value ),
    .io_exuWriteback_23_bits_vecWen ( io_exuWriteback_23_bits_vecWen ),
    .io_exuWriteback_23_bits_v0Wen ( io_exuWriteback_23_bits_v0Wen ),
    .io_exuWriteback_23_bits_vls_vdIdx ( io_exuWriteback_23_bits_vls_vdIdx ),
    .io_exuWriteback_23_bits_debug_isMMIO ( io_exuWriteback_23_bits_debug_isMMIO ),
    .io_exuWriteback_23_bits_debug_isNCIO ( io_exuWriteback_23_bits_debug_isNCIO ),
    .io_exuWriteback_23_bits_debug_isPerfCnt ( io_exuWriteback_23_bits_debug_isPerfCnt ),
    .io_exuWriteback_23_bits_debug_paddr ( io_exuWriteback_23_bits_debug_paddr ),
    .io_exuWriteback_22_valid ( io_exuWriteback_22_valid ),
    .io_exuWriteback_22_bits_data_0 ( io_exuWriteback_22_bits_data_0 ),
    .io_exuWriteback_22_bits_robIdx_value ( io_exuWriteback_22_bits_robIdx_value ),
    .io_exuWriteback_22_bits_lqIdx_value ( io_exuWriteback_22_bits_lqIdx_value ),
    .io_exuWriteback_22_bits_debug_isMMIO ( io_exuWriteback_22_bits_debug_isMMIO ),
    .io_exuWriteback_22_bits_debug_isNCIO ( io_exuWriteback_22_bits_debug_isNCIO ),
    .io_exuWriteback_22_bits_debug_isPerfCnt ( io_exuWriteback_22_bits_debug_isPerfCnt ),
    .io_exuWriteback_22_bits_debug_paddr ( io_exuWriteback_22_bits_debug_paddr ),
    .io_exuWriteback_21_valid ( io_exuWriteback_21_valid ),
    .io_exuWriteback_21_bits_data_0 ( io_exuWriteback_21_bits_data_0 ),
    .io_exuWriteback_21_bits_robIdx_value ( io_exuWriteback_21_bits_robIdx_value ),
    .io_exuWriteback_21_bits_lqIdx_value ( io_exuWriteback_21_bits_lqIdx_value ),
    .io_exuWriteback_21_bits_debug_isMMIO ( io_exuWriteback_21_bits_debug_isMMIO ),
    .io_exuWriteback_21_bits_debug_isNCIO ( io_exuWriteback_21_bits_debug_isNCIO ),
    .io_exuWriteback_21_bits_debug_isPerfCnt ( io_exuWriteback_21_bits_debug_isPerfCnt ),
    .io_exuWriteback_21_bits_debug_paddr ( io_exuWriteback_21_bits_debug_paddr ),
    .io_exuWriteback_20_valid ( io_exuWriteback_20_valid ),
    .io_exuWriteback_20_bits_data_0 ( io_exuWriteback_20_bits_data_0 ),
    .io_exuWriteback_20_bits_robIdx_value ( io_exuWriteback_20_bits_robIdx_value ),
    .io_exuWriteback_20_bits_lqIdx_value ( io_exuWriteback_20_bits_lqIdx_value ),
    .io_exuWriteback_20_bits_debug_isMMIO ( io_exuWriteback_20_bits_debug_isMMIO ),
    .io_exuWriteback_20_bits_debug_isNCIO ( io_exuWriteback_20_bits_debug_isNCIO ),
    .io_exuWriteback_20_bits_debug_isPerfCnt ( io_exuWriteback_20_bits_debug_isPerfCnt ),
    .io_exuWriteback_20_bits_debug_paddr ( io_exuWriteback_20_bits_debug_paddr ),
    .io_exuWriteback_19_valid ( io_exuWriteback_19_valid ),
    .io_exuWriteback_19_bits_data_0 ( io_exuWriteback_19_bits_data_0 ),
    .io_exuWriteback_19_bits_robIdx_value ( io_exuWriteback_19_bits_robIdx_value ),
    .io_exuWriteback_19_bits_sqIdx_value ( io_exuWriteback_19_bits_sqIdx_value ),
    .io_exuWriteback_19_bits_debug_isMMIO ( io_exuWriteback_19_bits_debug_isMMIO ),
    .io_exuWriteback_19_bits_debug_isNCIO ( io_exuWriteback_19_bits_debug_isNCIO ),
    .io_exuWriteback_19_bits_debug_isPerfCnt ( io_exuWriteback_19_bits_debug_isPerfCnt ),
    .io_exuWriteback_19_bits_debug_paddr ( io_exuWriteback_19_bits_debug_paddr ),
    .io_exuWriteback_18_valid ( io_exuWriteback_18_valid ),
    .io_exuWriteback_18_bits_data_0 ( io_exuWriteback_18_bits_data_0 ),
    .io_exuWriteback_18_bits_robIdx_value ( io_exuWriteback_18_bits_robIdx_value ),
    .io_exuWriteback_18_bits_sqIdx_value ( io_exuWriteback_18_bits_sqIdx_value ),
    .io_exuWriteback_18_bits_debug_isMMIO ( io_exuWriteback_18_bits_debug_isMMIO ),
    .io_exuWriteback_18_bits_debug_isNCIO ( io_exuWriteback_18_bits_debug_isNCIO ),
    .io_exuWriteback_18_bits_debug_isPerfCnt ( io_exuWriteback_18_bits_debug_isPerfCnt ),
    .io_exuWriteback_18_bits_debug_paddr ( io_exuWriteback_18_bits_debug_paddr ),
    .io_exuWriteback_17_valid ( io_exuWriteback_17_valid ),
    .io_exuWriteback_17_bits_data_0 ( io_exuWriteback_17_bits_data_0 ),
    .io_exuWriteback_17_bits_robIdx_value ( io_exuWriteback_17_bits_robIdx_value ),
    .io_exuWriteback_17_bits_fflags ( io_exuWriteback_17_bits_fflags ),
    .io_exuWriteback_17_bits_wflags ( io_exuWriteback_17_bits_wflags ),
    .io_exuWriteback_16_valid ( io_exuWriteback_16_valid ),
    .io_exuWriteback_16_bits_data_0 ( io_exuWriteback_16_bits_data_0 ),
    .io_exuWriteback_16_bits_robIdx_value ( io_exuWriteback_16_bits_robIdx_value ),
    .io_exuWriteback_16_bits_fflags ( io_exuWriteback_16_bits_fflags ),
    .io_exuWriteback_16_bits_wflags ( io_exuWriteback_16_bits_wflags ),
    .io_exuWriteback_15_valid ( io_exuWriteback_15_valid ),
    .io_exuWriteback_15_bits_data_0 ( io_exuWriteback_15_bits_data_0 ),
    .io_exuWriteback_15_bits_robIdx_value ( io_exuWriteback_15_bits_robIdx_value ),
    .io_exuWriteback_15_bits_fflags ( io_exuWriteback_15_bits_fflags ),
    .io_exuWriteback_15_bits_wflags ( io_exuWriteback_15_bits_wflags ),
    .io_exuWriteback_15_bits_vxsat ( io_exuWriteback_15_bits_vxsat ),
    .io_exuWriteback_14_valid ( io_exuWriteback_14_valid ),
    .io_exuWriteback_14_bits_data_0 ( io_exuWriteback_14_bits_data_0 ),
    .io_exuWriteback_14_bits_robIdx_value ( io_exuWriteback_14_bits_robIdx_value ),
    .io_exuWriteback_14_bits_fflags ( io_exuWriteback_14_bits_fflags ),
    .io_exuWriteback_14_bits_wflags ( io_exuWriteback_14_bits_wflags ),
    .io_exuWriteback_13_valid ( io_exuWriteback_13_valid ),
    .io_exuWriteback_13_bits_data_0 ( io_exuWriteback_13_bits_data_0 ),
    .io_exuWriteback_13_bits_robIdx_value ( io_exuWriteback_13_bits_robIdx_value ),
    .io_exuWriteback_13_bits_fflags ( io_exuWriteback_13_bits_fflags ),
    .io_exuWriteback_13_bits_wflags ( io_exuWriteback_13_bits_wflags ),
    .io_exuWriteback_13_bits_vxsat ( io_exuWriteback_13_bits_vxsat ),
    .io_exuWriteback_12_valid ( io_exuWriteback_12_valid ),
    .io_exuWriteback_12_bits_data_0 ( io_exuWriteback_12_bits_data_0 ),
    .io_exuWriteback_12_bits_robIdx_value ( io_exuWriteback_12_bits_robIdx_value ),
    .io_exuWriteback_12_bits_fflags ( io_exuWriteback_12_bits_fflags ),
    .io_exuWriteback_12_bits_wflags ( io_exuWriteback_12_bits_wflags ),
    .io_exuWriteback_11_valid ( io_exuWriteback_11_valid ),
    .io_exuWriteback_11_bits_data_0 ( io_exuWriteback_11_bits_data_0 ),
    .io_exuWriteback_11_bits_robIdx_value ( io_exuWriteback_11_bits_robIdx_value ),
    .io_exuWriteback_11_bits_fflags ( io_exuWriteback_11_bits_fflags ),
    .io_exuWriteback_11_bits_wflags ( io_exuWriteback_11_bits_wflags ),
    .io_exuWriteback_10_valid ( io_exuWriteback_10_valid ),
    .io_exuWriteback_10_bits_data_0 ( io_exuWriteback_10_bits_data_0 ),
    .io_exuWriteback_10_bits_robIdx_value ( io_exuWriteback_10_bits_robIdx_value ),
    .io_exuWriteback_10_bits_fflags ( io_exuWriteback_10_bits_fflags ),
    .io_exuWriteback_10_bits_wflags ( io_exuWriteback_10_bits_wflags ),
    .io_exuWriteback_9_valid ( io_exuWriteback_9_valid ),
    .io_exuWriteback_9_bits_data_0 ( io_exuWriteback_9_bits_data_0 ),
    .io_exuWriteback_9_bits_robIdx_value ( io_exuWriteback_9_bits_robIdx_value ),
    .io_exuWriteback_9_bits_fflags ( io_exuWriteback_9_bits_fflags ),
    .io_exuWriteback_9_bits_wflags ( io_exuWriteback_9_bits_wflags ),
    .io_exuWriteback_8_valid ( io_exuWriteback_8_valid ),
    .io_exuWriteback_8_bits_data_0 ( io_exuWriteback_8_bits_data_0 ),
    .io_exuWriteback_8_bits_robIdx_value ( io_exuWriteback_8_bits_robIdx_value ),
    .io_exuWriteback_8_bits_fflags ( io_exuWriteback_8_bits_fflags ),
    .io_exuWriteback_8_bits_wflags ( io_exuWriteback_8_bits_wflags ),
    .io_exuWriteback_7_valid ( io_exuWriteback_7_valid ),
    .io_exuWriteback_7_bits_data_0 ( io_exuWriteback_7_bits_data_0 ),
    .io_exuWriteback_7_bits_robIdx_value ( io_exuWriteback_7_bits_robIdx_value ),
    .io_exuWriteback_7_bits_debug_isPerfCnt ( io_exuWriteback_7_bits_debug_isPerfCnt ),
    .io_exuWriteback_6_valid ( io_exuWriteback_6_valid ),
    .io_exuWriteback_6_bits_data_0 ( io_exuWriteback_6_bits_data_0 ),
    .io_exuWriteback_6_bits_robIdx_value ( io_exuWriteback_6_bits_robIdx_value ),
    .io_exuWriteback_5_valid ( io_exuWriteback_5_valid ),
    .io_exuWriteback_5_bits_data_0 ( io_exuWriteback_5_bits_data_0 ),
    .io_exuWriteback_5_bits_robIdx_value ( io_exuWriteback_5_bits_robIdx_value ),
    .io_exuWriteback_5_bits_redirect_valid ( io_exuWriteback_5_bits_redirect_valid ),
    .io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken ( io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken ),
    .io_exuWriteback_5_bits_fflags ( io_exuWriteback_5_bits_fflags ),
    .io_exuWriteback_5_bits_wflags ( io_exuWriteback_5_bits_wflags ),
    .io_exuWriteback_4_valid ( io_exuWriteback_4_valid ),
    .io_exuWriteback_4_bits_data_0 ( io_exuWriteback_4_bits_data_0 ),
    .io_exuWriteback_4_bits_robIdx_value ( io_exuWriteback_4_bits_robIdx_value ),
    .io_exuWriteback_3_valid ( io_exuWriteback_3_valid ),
    .io_exuWriteback_3_bits_data_0 ( io_exuWriteback_3_bits_data_0 ),
    .io_exuWriteback_3_bits_robIdx_value ( io_exuWriteback_3_bits_robIdx_value ),
    .io_exuWriteback_3_bits_redirect_valid ( io_exuWriteback_3_bits_redirect_valid ),
    .io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken ( io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken ),
    .io_exuWriteback_2_valid ( io_exuWriteback_2_valid ),
    .io_exuWriteback_2_bits_data_0 ( io_exuWriteback_2_bits_data_0 ),
    .io_exuWriteback_2_bits_robIdx_value ( io_exuWriteback_2_bits_robIdx_value ),
    .io_exuWriteback_1_valid ( io_exuWriteback_1_valid ),
    .io_exuWriteback_1_bits_data_0 ( io_exuWriteback_1_bits_data_0 ),
    .io_exuWriteback_1_bits_robIdx_value ( io_exuWriteback_1_bits_robIdx_value ),
    .io_exuWriteback_1_bits_redirect_valid ( io_exuWriteback_1_bits_redirect_valid ),
    .io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken ( io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken ),
    .io_exuWriteback_0_valid ( io_exuWriteback_0_valid ),
    .io_exuWriteback_0_bits_data_0 ( io_exuWriteback_0_bits_data_0 ),
    .io_exuWriteback_0_bits_robIdx_value ( io_exuWriteback_0_bits_robIdx_value ),
    .io_writebackNums_0_bits ( io_writebackNums_0_bits ),
    .io_writebackNums_1_bits ( io_writebackNums_1_bits ),
    .io_writebackNums_2_bits ( io_writebackNums_2_bits ),
    .io_writebackNums_3_bits ( io_writebackNums_3_bits ),
    .io_writebackNums_4_bits ( io_writebackNums_4_bits ),
    .io_writebackNums_5_bits ( io_writebackNums_5_bits ),
    .io_writebackNums_6_bits ( io_writebackNums_6_bits ),
    .io_writebackNums_7_bits ( io_writebackNums_7_bits ),
    .io_writebackNums_8_bits ( io_writebackNums_8_bits ),
    .io_writebackNums_9_bits ( io_writebackNums_9_bits ),
    .io_writebackNums_10_bits ( io_writebackNums_10_bits ),
    .io_writebackNums_11_bits ( io_writebackNums_11_bits ),
    .io_writebackNums_12_bits ( io_writebackNums_12_bits ),
    .io_writebackNums_13_bits ( io_writebackNums_13_bits ),
    .io_writebackNums_14_bits ( io_writebackNums_14_bits ),
    .io_writebackNums_15_bits ( io_writebackNums_15_bits ),
    .io_writebackNums_16_bits ( io_writebackNums_16_bits ),
    .io_writebackNums_17_bits ( io_writebackNums_17_bits ),
    .io_writebackNums_18_bits ( io_writebackNums_18_bits ),
    .io_writebackNums_19_bits ( io_writebackNums_19_bits ),
    .io_writebackNums_20_bits ( io_writebackNums_20_bits ),
    .io_writebackNums_21_bits ( io_writebackNums_21_bits ),
    .io_writebackNums_22_bits ( io_writebackNums_22_bits ),
    .io_writebackNums_23_bits ( io_writebackNums_23_bits ),
    .io_writebackNums_24_bits ( io_writebackNums_24_bits ),
    .io_writebackNeedFlush_0 ( io_writebackNeedFlush_0 ),
    .io_writebackNeedFlush_1 ( io_writebackNeedFlush_1 ),
    .io_writebackNeedFlush_2 ( io_writebackNeedFlush_2 ),
    .io_writebackNeedFlush_6 ( io_writebackNeedFlush_6 ),
    .io_writebackNeedFlush_7 ( io_writebackNeedFlush_7 ),
    .io_writebackNeedFlush_8 ( io_writebackNeedFlush_8 ),
    .io_writebackNeedFlush_9 ( io_writebackNeedFlush_9 ),
    .io_writebackNeedFlush_10 ( io_writebackNeedFlush_10 ),
    .io_writebackNeedFlush_11 ( io_writebackNeedFlush_11 ),
    .io_writebackNeedFlush_12 ( io_writebackNeedFlush_12 ),
    //Redirect_in
    .io_redirect_valid    ( io_redirect_valid    ),
    .io_redirect_bits_robIdx_flag ( io_redirect_bits_robIdx_flag ),
    .io_redirect_bits_robIdx_value ( io_redirect_bits_robIdx_value ),
    .io_redirect_bits_level ( io_redirect_bits_level ),
    //CSR_in
    .io_csr_intrBitSet    ( io_csr_intrBitSet    ),
    .io_csr_wfiEvent      ( io_csr_wfiEvent      ),
    .io_csr_criticalErrorState ( io_csr_criticalErrorState ),
    .io_snpt_snptDeq      ( io_snpt_snptDeq      ),
    .io_snpt_useSnpt      ( io_snpt_useSnpt      ),
    .io_snpt_snptSelect   ( io_snpt_snptSelect   ),
    .io_snpt_flushVec_0   ( io_snpt_flushVec_0   ),
    .io_snpt_flushVec_1   ( io_snpt_flushVec_1   ),
    .io_snpt_flushVec_2   ( io_snpt_flushVec_2   ),
    .io_snpt_flushVec_3   ( io_snpt_flushVec_3   ),
    .io_wfi_safeFromMem   ( io_wfi_safeFromMem   ),
    .io_wfi_safeFromFrontend ( io_wfi_safeFromFrontend ),
    .io_wfi_enable        ( io_wfi_enable        ),
    .io_fromVecExcpMod_busy ( io_fromVecExcpMod_busy ),
    .io_readGPAMemData_gpaddr ( io_readGPAMemData_gpaddr ),
    .io_readGPAMemData_isForVSnonLeafPTE ( io_readGPAMemData_isForVSnonLeafPTE ),
    .io_vstartIsZero      ( io_vstartIsZero      ),
    .io_debugEnqLsq_canAccept ( io_debugEnqLsq_canAccept ),
    .io_debugEnqLsq_needAlloc_0 ( io_debugEnqLsq_needAlloc_0 ),
    .io_debugEnqLsq_needAlloc_1 ( io_debugEnqLsq_needAlloc_1 ),
    .io_debugEnqLsq_needAlloc_2 ( io_debugEnqLsq_needAlloc_2 ),
    .io_debugEnqLsq_needAlloc_3 ( io_debugEnqLsq_needAlloc_3 ),
    .io_debugEnqLsq_needAlloc_4 ( io_debugEnqLsq_needAlloc_4 ),
    .io_debugEnqLsq_needAlloc_5 ( io_debugEnqLsq_needAlloc_5 ),
    .io_debugEnqLsq_req_0_valid ( io_debugEnqLsq_req_0_valid ),
    .io_debugEnqLsq_req_0_bits_robIdx_value ( io_debugEnqLsq_req_0_bits_robIdx_value ),
    .io_debugEnqLsq_req_0_bits_lqIdx_value ( io_debugEnqLsq_req_0_bits_lqIdx_value ),
    .io_debugEnqLsq_req_1_valid ( io_debugEnqLsq_req_1_valid ),
    .io_debugEnqLsq_req_1_bits_robIdx_value ( io_debugEnqLsq_req_1_bits_robIdx_value ),
    .io_debugEnqLsq_req_1_bits_lqIdx_value ( io_debugEnqLsq_req_1_bits_lqIdx_value ),
    .io_debugEnqLsq_req_2_valid ( io_debugEnqLsq_req_2_valid ),
    .io_debugEnqLsq_req_2_bits_robIdx_value ( io_debugEnqLsq_req_2_bits_robIdx_value ),
    .io_debugEnqLsq_req_2_bits_lqIdx_value ( io_debugEnqLsq_req_2_bits_lqIdx_value ),
    .io_debugEnqLsq_req_3_valid ( io_debugEnqLsq_req_3_valid ),
    .io_debugEnqLsq_req_3_bits_robIdx_value ( io_debugEnqLsq_req_3_bits_robIdx_value ),
    .io_debugEnqLsq_req_3_bits_lqIdx_value ( io_debugEnqLsq_req_3_bits_lqIdx_value ),
    .io_debugEnqLsq_req_4_valid ( io_debugEnqLsq_req_4_valid ),
    .io_debugEnqLsq_req_4_bits_robIdx_value ( io_debugEnqLsq_req_4_bits_robIdx_value ),
    .io_debugEnqLsq_req_4_bits_lqIdx_value ( io_debugEnqLsq_req_4_bits_lqIdx_value ),
    .io_debugEnqLsq_req_5_valid ( io_debugEnqLsq_req_5_valid ),
    .io_debugEnqLsq_req_5_bits_robIdx_value ( io_debugEnqLsq_req_5_bits_robIdx_value ),
    .io_debugEnqLsq_req_5_bits_lqIdx_value ( io_debugEnqLsq_req_5_bits_lqIdx_value ),
    .io_debugInstrAddrTransType_bare ( io_debugInstrAddrTransType_bare ),
    .io_debugInstrAddrTransType_sv39 ( io_debugInstrAddrTransType_sv39 ),
    .io_debugInstrAddrTransType_sv39x4 ( io_debugInstrAddrTransType_sv39x4 ),
    .io_debugInstrAddrTransType_sv48 ( io_debugInstrAddrTransType_sv48 ),
    .io_debugInstrAddrTransType_sv48x4 ( io_debugInstrAddrTransType_sv48x4 ),
    .io_storeDebugInfo_0_robidx_value ( io_storeDebugInfo_0_robidx_value ),
    .io_storeDebugInfo_1_robidx_value ( io_storeDebugInfo_1_robidx_value ),
    //Mem_in
    .io_lsq_mmio_0        ( io_lsq_mmio_0        ),
    .io_lsq_mmio_1        ( io_lsq_mmio_1        ),
    .io_lsq_mmio_2        ( io_lsq_mmio_2        ),
    .io_lsq_uop_0_robIdx_value ( io_lsq_uop_0_robIdx_value ),
    .io_lsq_uop_1_robIdx_value ( io_lsq_uop_1_robIdx_value ),
    .io_lsq_uop_2_robIdx_value ( io_lsq_uop_2_robIdx_value ),
    //Rob_output
    .io_enq_canAccept     ( io_enq_canAccept     ),
    .io_enq_canAcceptForDispatch ( io_enq_canAcceptForDispatch ),
    .io_enq_isEmpty       ( io_enq_isEmpty       ),
    .io_flushOut_valid    ( io_flushOut_valid    ),
    .io_flushOut_bits_isRVC ( io_flushOut_bits_isRVC ),
    .io_flushOut_bits_robIdx_flag ( io_flushOut_bits_robIdx_flag ),
    .io_flushOut_bits_robIdx_value ( io_flushOut_bits_robIdx_value ),
    .io_flushOut_bits_ftqIdx_flag ( io_flushOut_bits_ftqIdx_flag ),
    .io_flushOut_bits_ftqIdx_value ( io_flushOut_bits_ftqIdx_value ),
    .io_flushOut_bits_ftqOffset ( io_flushOut_bits_ftqOffset ),
    .io_flushOut_bits_level ( io_flushOut_bits_level ),
    .io_exception_valid   ( io_exception_valid   ),
    .io_exception_bits_instr ( io_exception_bits_instr ),
    .io_exception_bits_commitType ( io_exception_bits_commitType ),
    .io_exception_bits_exceptionVec_0 ( io_exception_bits_exceptionVec_0 ),
    .io_exception_bits_exceptionVec_1 ( io_exception_bits_exceptionVec_1 ),
    .io_exception_bits_exceptionVec_2 ( io_exception_bits_exceptionVec_2 ),
    .io_exception_bits_exceptionVec_3 ( io_exception_bits_exceptionVec_3 ),
    .io_exception_bits_exceptionVec_4 ( io_exception_bits_exceptionVec_4 ),
    .io_exception_bits_exceptionVec_5 ( io_exception_bits_exceptionVec_5 ),
    .io_exception_bits_exceptionVec_6 ( io_exception_bits_exceptionVec_6 ),
    .io_exception_bits_exceptionVec_7 ( io_exception_bits_exceptionVec_7 ),
    .io_exception_bits_exceptionVec_8 ( io_exception_bits_exceptionVec_8 ),
    .io_exception_bits_exceptionVec_9 ( io_exception_bits_exceptionVec_9 ),
    .io_exception_bits_exceptionVec_10 ( io_exception_bits_exceptionVec_10 ),
    .io_exception_bits_exceptionVec_11 ( io_exception_bits_exceptionVec_11 ),
    .io_exception_bits_exceptionVec_12 ( io_exception_bits_exceptionVec_12 ),
    .io_exception_bits_exceptionVec_13 ( io_exception_bits_exceptionVec_13 ),
    .io_exception_bits_exceptionVec_14 ( io_exception_bits_exceptionVec_14 ),
    .io_exception_bits_exceptionVec_15 ( io_exception_bits_exceptionVec_15 ),
    .io_exception_bits_exceptionVec_16 ( io_exception_bits_exceptionVec_16 ),
    .io_exception_bits_exceptionVec_17 ( io_exception_bits_exceptionVec_17 ),
    .io_exception_bits_exceptionVec_18 ( io_exception_bits_exceptionVec_18 ),
    .io_exception_bits_exceptionVec_19 ( io_exception_bits_exceptionVec_19 ),
    .io_exception_bits_exceptionVec_20 ( io_exception_bits_exceptionVec_20 ),
    .io_exception_bits_exceptionVec_21 ( io_exception_bits_exceptionVec_21 ),
    .io_exception_bits_exceptionVec_22 ( io_exception_bits_exceptionVec_22 ),
    .io_exception_bits_exceptionVec_23 ( io_exception_bits_exceptionVec_23 ),
    .io_exception_bits_isPcBkpt ( io_exception_bits_isPcBkpt ),
    .io_exception_bits_isFetchMalAddr ( io_exception_bits_isFetchMalAddr ),
    .io_exception_bits_gpaddr ( io_exception_bits_gpaddr ),
    .io_exception_bits_singleStep ( io_exception_bits_singleStep ),
    .io_exception_bits_crossPageIPFFix ( io_exception_bits_crossPageIPFFix ),
    .io_exception_bits_isInterrupt ( io_exception_bits_isInterrupt ),
    .io_exception_bits_isHls ( io_exception_bits_isHls ),
    .io_exception_bits_trigger ( io_exception_bits_trigger ),
    .io_exception_bits_isForVSnonLeafPTE ( io_exception_bits_isForVSnonLeafPTE ),
    .io_commits_isCommit  ( io_commits_isCommit  ),
    .io_commits_commitValid_0 ( io_commits_commitValid_0 ),
    .io_commits_commitValid_1 ( io_commits_commitValid_1 ),
    .io_commits_commitValid_2 ( io_commits_commitValid_2 ),
    .io_commits_commitValid_3 ( io_commits_commitValid_3 ),
    .io_commits_commitValid_4 ( io_commits_commitValid_4 ),
    .io_commits_commitValid_5 ( io_commits_commitValid_5 ),
    .io_commits_commitValid_6 ( io_commits_commitValid_6 ),
    .io_commits_commitValid_7 ( io_commits_commitValid_7 ),
    .io_commits_isWalk    ( io_commits_isWalk    ),
    .io_commits_walkValid_0 ( io_commits_walkValid_0 ),
    .io_commits_walkValid_1 ( io_commits_walkValid_1 ),
    .io_commits_walkValid_2 ( io_commits_walkValid_2 ),
    .io_commits_walkValid_3 ( io_commits_walkValid_3 ),
    .io_commits_walkValid_4 ( io_commits_walkValid_4 ),
    .io_commits_walkValid_5 ( io_commits_walkValid_5 ),
    .io_commits_walkValid_6 ( io_commits_walkValid_6 ),
    .io_commits_walkValid_7 ( io_commits_walkValid_7 ),
    .io_commits_info_0_walk_v ( io_commits_info_0_walk_v ),
    .io_commits_info_0_commit_v ( io_commits_info_0_commit_v ),
    .io_commits_info_0_commit_w ( io_commits_info_0_commit_w ),
    .io_commits_info_0_realDestSize ( io_commits_info_0_realDestSize ),
    .io_commits_info_0_interrupt_safe ( io_commits_info_0_interrupt_safe ),
    .io_commits_info_0_wflags ( io_commits_info_0_wflags ),
    .io_commits_info_0_fflags ( io_commits_info_0_fflags ),
    .io_commits_info_0_vxsat ( io_commits_info_0_vxsat ),
    .io_commits_info_0_isRVC ( io_commits_info_0_isRVC ),
    .io_commits_info_0_isVset ( io_commits_info_0_isVset ),
    .io_commits_info_0_isHls ( io_commits_info_0_isHls ),
    .io_commits_info_0_isVls ( io_commits_info_0_isVls ),
    .io_commits_info_0_vls ( io_commits_info_0_vls ),
    .io_commits_info_0_mmio ( io_commits_info_0_mmio ),
    .io_commits_info_0_commitType ( io_commits_info_0_commitType ),
    .io_commits_info_0_ftqIdx_flag ( io_commits_info_0_ftqIdx_flag ),
    .io_commits_info_0_ftqIdx_value ( io_commits_info_0_ftqIdx_value ),
    .io_commits_info_0_ftqOffset ( io_commits_info_0_ftqOffset ),
    .io_commits_info_0_instrSize ( io_commits_info_0_instrSize ),
    .io_commits_info_0_fpWen ( io_commits_info_0_fpWen ),
    .io_commits_info_0_rfWen ( io_commits_info_0_rfWen ),
    .io_commits_info_0_needFlush ( io_commits_info_0_needFlush ),
    .io_commits_info_0_traceBlockInPipe_itype ( io_commits_info_0_traceBlockInPipe_itype ),
    .io_commits_info_0_traceBlockInPipe_iretire ( io_commits_info_0_traceBlockInPipe_iretire ),
    .io_commits_info_0_traceBlockInPipe_ilastsize ( io_commits_info_0_traceBlockInPipe_ilastsize ),
    .io_commits_info_0_debug_pc ( io_commits_info_0_debug_pc ),
    .io_commits_info_0_debug_instr ( io_commits_info_0_debug_instr ),
    .io_commits_info_0_debug_ldest ( io_commits_info_0_debug_ldest ),
    .io_commits_info_0_debug_pdest ( io_commits_info_0_debug_pdest ),
    .io_commits_info_0_debug_otherPdest_0 ( io_commits_info_0_debug_otherPdest_0 ),
    .io_commits_info_0_debug_otherPdest_1 ( io_commits_info_0_debug_otherPdest_1 ),
    .io_commits_info_0_debug_otherPdest_2 ( io_commits_info_0_debug_otherPdest_2 ),
    .io_commits_info_0_debug_otherPdest_3 ( io_commits_info_0_debug_otherPdest_3 ),
    .io_commits_info_0_debug_otherPdest_4 ( io_commits_info_0_debug_otherPdest_4 ),
    .io_commits_info_0_debug_otherPdest_5 ( io_commits_info_0_debug_otherPdest_5 ),
    .io_commits_info_0_debug_otherPdest_6 ( io_commits_info_0_debug_otherPdest_6 ),
    .io_commits_info_0_debug_fuType ( io_commits_info_0_debug_fuType ),
    .io_commits_info_0_dirtyFs ( io_commits_info_0_dirtyFs ),
    .io_commits_info_0_dirtyVs ( io_commits_info_0_dirtyVs ),
    .io_commits_info_1_walk_v ( io_commits_info_1_walk_v ),
    .io_commits_info_1_commit_v ( io_commits_info_1_commit_v ),
    .io_commits_info_1_commit_w ( io_commits_info_1_commit_w ),
    .io_commits_info_1_realDestSize ( io_commits_info_1_realDestSize ),
    .io_commits_info_1_interrupt_safe ( io_commits_info_1_interrupt_safe ),
    .io_commits_info_1_wflags ( io_commits_info_1_wflags ),
    .io_commits_info_1_fflags ( io_commits_info_1_fflags ),
    .io_commits_info_1_vxsat ( io_commits_info_1_vxsat ),
    .io_commits_info_1_isRVC ( io_commits_info_1_isRVC ),
    .io_commits_info_1_isVset ( io_commits_info_1_isVset ),
    .io_commits_info_1_isHls ( io_commits_info_1_isHls ),
    .io_commits_info_1_isVls ( io_commits_info_1_isVls ),
    .io_commits_info_1_vls ( io_commits_info_1_vls ),
    .io_commits_info_1_mmio ( io_commits_info_1_mmio ),
    .io_commits_info_1_commitType ( io_commits_info_1_commitType ),
    .io_commits_info_1_ftqIdx_flag ( io_commits_info_1_ftqIdx_flag ),
    .io_commits_info_1_ftqIdx_value ( io_commits_info_1_ftqIdx_value ),
    .io_commits_info_1_ftqOffset ( io_commits_info_1_ftqOffset ),
    .io_commits_info_1_instrSize ( io_commits_info_1_instrSize ),
    .io_commits_info_1_fpWen ( io_commits_info_1_fpWen ),
    .io_commits_info_1_rfWen ( io_commits_info_1_rfWen ),
    .io_commits_info_1_needFlush ( io_commits_info_1_needFlush ),
    .io_commits_info_1_traceBlockInPipe_itype ( io_commits_info_1_traceBlockInPipe_itype ),
    .io_commits_info_1_traceBlockInPipe_iretire ( io_commits_info_1_traceBlockInPipe_iretire ),
    .io_commits_info_1_traceBlockInPipe_ilastsize ( io_commits_info_1_traceBlockInPipe_ilastsize ),
    .io_commits_info_1_debug_pc ( io_commits_info_1_debug_pc ),
    .io_commits_info_1_debug_instr ( io_commits_info_1_debug_instr ),
    .io_commits_info_1_debug_ldest ( io_commits_info_1_debug_ldest ),
    .io_commits_info_1_debug_pdest ( io_commits_info_1_debug_pdest ),
    .io_commits_info_1_debug_otherPdest_0 ( io_commits_info_1_debug_otherPdest_0 ),
    .io_commits_info_1_debug_otherPdest_1 ( io_commits_info_1_debug_otherPdest_1 ),
    .io_commits_info_1_debug_otherPdest_2 ( io_commits_info_1_debug_otherPdest_2 ),
    .io_commits_info_1_debug_otherPdest_3 ( io_commits_info_1_debug_otherPdest_3 ),
    .io_commits_info_1_debug_otherPdest_4 ( io_commits_info_1_debug_otherPdest_4 ),
    .io_commits_info_1_debug_otherPdest_5 ( io_commits_info_1_debug_otherPdest_5 ),
    .io_commits_info_1_debug_otherPdest_6 ( io_commits_info_1_debug_otherPdest_6 ),
    .io_commits_info_1_debug_fuType ( io_commits_info_1_debug_fuType ),
    .io_commits_info_1_dirtyFs ( io_commits_info_1_dirtyFs ),
    .io_commits_info_1_dirtyVs ( io_commits_info_1_dirtyVs ),
    .io_commits_info_2_walk_v ( io_commits_info_2_walk_v ),
    .io_commits_info_2_commit_v ( io_commits_info_2_commit_v ),
    .io_commits_info_2_commit_w ( io_commits_info_2_commit_w ),
    .io_commits_info_2_realDestSize ( io_commits_info_2_realDestSize ),
    .io_commits_info_2_interrupt_safe ( io_commits_info_2_interrupt_safe ),
    .io_commits_info_2_wflags ( io_commits_info_2_wflags ),
    .io_commits_info_2_fflags ( io_commits_info_2_fflags ),
    .io_commits_info_2_vxsat ( io_commits_info_2_vxsat ),
    .io_commits_info_2_isRVC ( io_commits_info_2_isRVC ),
    .io_commits_info_2_isVset ( io_commits_info_2_isVset ),
    .io_commits_info_2_isHls ( io_commits_info_2_isHls ),
    .io_commits_info_2_isVls ( io_commits_info_2_isVls ),
    .io_commits_info_2_vls ( io_commits_info_2_vls ),
    .io_commits_info_2_mmio ( io_commits_info_2_mmio ),
    .io_commits_info_2_commitType ( io_commits_info_2_commitType ),
    .io_commits_info_2_ftqIdx_flag ( io_commits_info_2_ftqIdx_flag ),
    .io_commits_info_2_ftqIdx_value ( io_commits_info_2_ftqIdx_value ),
    .io_commits_info_2_ftqOffset ( io_commits_info_2_ftqOffset ),
    .io_commits_info_2_instrSize ( io_commits_info_2_instrSize ),
    .io_commits_info_2_fpWen ( io_commits_info_2_fpWen ),
    .io_commits_info_2_rfWen ( io_commits_info_2_rfWen ),
    .io_commits_info_2_needFlush ( io_commits_info_2_needFlush ),
    .io_commits_info_2_traceBlockInPipe_itype ( io_commits_info_2_traceBlockInPipe_itype ),
    .io_commits_info_2_traceBlockInPipe_iretire ( io_commits_info_2_traceBlockInPipe_iretire ),
    .io_commits_info_2_traceBlockInPipe_ilastsize ( io_commits_info_2_traceBlockInPipe_ilastsize ),
    .io_commits_info_2_debug_pc ( io_commits_info_2_debug_pc ),
    .io_commits_info_2_debug_instr ( io_commits_info_2_debug_instr ),
    .io_commits_info_2_debug_ldest ( io_commits_info_2_debug_ldest ),
    .io_commits_info_2_debug_pdest ( io_commits_info_2_debug_pdest ),
    .io_commits_info_2_debug_otherPdest_0 ( io_commits_info_2_debug_otherPdest_0 ),
    .io_commits_info_2_debug_otherPdest_1 ( io_commits_info_2_debug_otherPdest_1 ),
    .io_commits_info_2_debug_otherPdest_2 ( io_commits_info_2_debug_otherPdest_2 ),
    .io_commits_info_2_debug_otherPdest_3 ( io_commits_info_2_debug_otherPdest_3 ),
    .io_commits_info_2_debug_otherPdest_4 ( io_commits_info_2_debug_otherPdest_4 ),
    .io_commits_info_2_debug_otherPdest_5 ( io_commits_info_2_debug_otherPdest_5 ),
    .io_commits_info_2_debug_otherPdest_6 ( io_commits_info_2_debug_otherPdest_6 ),
    .io_commits_info_2_debug_fuType ( io_commits_info_2_debug_fuType ),
    .io_commits_info_2_dirtyFs ( io_commits_info_2_dirtyFs ),
    .io_commits_info_2_dirtyVs ( io_commits_info_2_dirtyVs ),
    .io_commits_info_3_walk_v ( io_commits_info_3_walk_v ),
    .io_commits_info_3_commit_v ( io_commits_info_3_commit_v ),
    .io_commits_info_3_commit_w ( io_commits_info_3_commit_w ),
    .io_commits_info_3_realDestSize ( io_commits_info_3_realDestSize ),
    .io_commits_info_3_interrupt_safe ( io_commits_info_3_interrupt_safe ),
    .io_commits_info_3_wflags ( io_commits_info_3_wflags ),
    .io_commits_info_3_fflags ( io_commits_info_3_fflags ),
    .io_commits_info_3_vxsat ( io_commits_info_3_vxsat ),
    .io_commits_info_3_isRVC ( io_commits_info_3_isRVC ),
    .io_commits_info_3_isVset ( io_commits_info_3_isVset ),
    .io_commits_info_3_isHls ( io_commits_info_3_isHls ),
    .io_commits_info_3_isVls ( io_commits_info_3_isVls ),
    .io_commits_info_3_vls ( io_commits_info_3_vls ),
    .io_commits_info_3_mmio ( io_commits_info_3_mmio ),
    .io_commits_info_3_commitType ( io_commits_info_3_commitType ),
    .io_commits_info_3_ftqIdx_flag ( io_commits_info_3_ftqIdx_flag ),
    .io_commits_info_3_ftqIdx_value ( io_commits_info_3_ftqIdx_value ),
    .io_commits_info_3_ftqOffset ( io_commits_info_3_ftqOffset ),
    .io_commits_info_3_instrSize ( io_commits_info_3_instrSize ),
    .io_commits_info_3_fpWen ( io_commits_info_3_fpWen ),
    .io_commits_info_3_rfWen ( io_commits_info_3_rfWen ),
    .io_commits_info_3_needFlush ( io_commits_info_3_needFlush ),
    .io_commits_info_3_traceBlockInPipe_itype ( io_commits_info_3_traceBlockInPipe_itype ),
    .io_commits_info_3_traceBlockInPipe_iretire ( io_commits_info_3_traceBlockInPipe_iretire ),
    .io_commits_info_3_traceBlockInPipe_ilastsize ( io_commits_info_3_traceBlockInPipe_ilastsize ),
    .io_commits_info_3_debug_pc ( io_commits_info_3_debug_pc ),
    .io_commits_info_3_debug_instr ( io_commits_info_3_debug_instr ),
    .io_commits_info_3_debug_ldest ( io_commits_info_3_debug_ldest ),
    .io_commits_info_3_debug_pdest ( io_commits_info_3_debug_pdest ),
    .io_commits_info_3_debug_otherPdest_0 ( io_commits_info_3_debug_otherPdest_0 ),
    .io_commits_info_3_debug_otherPdest_1 ( io_commits_info_3_debug_otherPdest_1 ),
    .io_commits_info_3_debug_otherPdest_2 ( io_commits_info_3_debug_otherPdest_2 ),
    .io_commits_info_3_debug_otherPdest_3 ( io_commits_info_3_debug_otherPdest_3 ),
    .io_commits_info_3_debug_otherPdest_4 ( io_commits_info_3_debug_otherPdest_4 ),
    .io_commits_info_3_debug_otherPdest_5 ( io_commits_info_3_debug_otherPdest_5 ),
    .io_commits_info_3_debug_otherPdest_6 ( io_commits_info_3_debug_otherPdest_6 ),
    .io_commits_info_3_debug_fuType ( io_commits_info_3_debug_fuType ),
    .io_commits_info_3_dirtyFs ( io_commits_info_3_dirtyFs ),
    .io_commits_info_3_dirtyVs ( io_commits_info_3_dirtyVs ),
    .io_commits_info_4_walk_v ( io_commits_info_4_walk_v ),
    .io_commits_info_4_commit_v ( io_commits_info_4_commit_v ),
    .io_commits_info_4_commit_w ( io_commits_info_4_commit_w ),
    .io_commits_info_4_realDestSize ( io_commits_info_4_realDestSize ),
    .io_commits_info_4_interrupt_safe ( io_commits_info_4_interrupt_safe ),
    .io_commits_info_4_wflags ( io_commits_info_4_wflags ),
    .io_commits_info_4_fflags ( io_commits_info_4_fflags ),
    .io_commits_info_4_vxsat ( io_commits_info_4_vxsat ),
    .io_commits_info_4_isRVC ( io_commits_info_4_isRVC ),
    .io_commits_info_4_isVset ( io_commits_info_4_isVset ),
    .io_commits_info_4_isHls ( io_commits_info_4_isHls ),
    .io_commits_info_4_isVls ( io_commits_info_4_isVls ),
    .io_commits_info_4_vls ( io_commits_info_4_vls ),
    .io_commits_info_4_mmio ( io_commits_info_4_mmio ),
    .io_commits_info_4_commitType ( io_commits_info_4_commitType ),
    .io_commits_info_4_ftqIdx_flag ( io_commits_info_4_ftqIdx_flag ),
    .io_commits_info_4_ftqIdx_value ( io_commits_info_4_ftqIdx_value ),
    .io_commits_info_4_ftqOffset ( io_commits_info_4_ftqOffset ),
    .io_commits_info_4_instrSize ( io_commits_info_4_instrSize ),
    .io_commits_info_4_fpWen ( io_commits_info_4_fpWen ),
    .io_commits_info_4_rfWen ( io_commits_info_4_rfWen ),
    .io_commits_info_4_needFlush ( io_commits_info_4_needFlush ),
    .io_commits_info_4_traceBlockInPipe_itype ( io_commits_info_4_traceBlockInPipe_itype ),
    .io_commits_info_4_traceBlockInPipe_iretire ( io_commits_info_4_traceBlockInPipe_iretire ),
    .io_commits_info_4_traceBlockInPipe_ilastsize ( io_commits_info_4_traceBlockInPipe_ilastsize ),
    .io_commits_info_4_debug_pc ( io_commits_info_4_debug_pc ),
    .io_commits_info_4_debug_instr ( io_commits_info_4_debug_instr ),
    .io_commits_info_4_debug_ldest ( io_commits_info_4_debug_ldest ),
    .io_commits_info_4_debug_pdest ( io_commits_info_4_debug_pdest ),
    .io_commits_info_4_debug_otherPdest_0 ( io_commits_info_4_debug_otherPdest_0 ),
    .io_commits_info_4_debug_otherPdest_1 ( io_commits_info_4_debug_otherPdest_1 ),
    .io_commits_info_4_debug_otherPdest_2 ( io_commits_info_4_debug_otherPdest_2 ),
    .io_commits_info_4_debug_otherPdest_3 ( io_commits_info_4_debug_otherPdest_3 ),
    .io_commits_info_4_debug_otherPdest_4 ( io_commits_info_4_debug_otherPdest_4 ),
    .io_commits_info_4_debug_otherPdest_5 ( io_commits_info_4_debug_otherPdest_5 ),
    .io_commits_info_4_debug_otherPdest_6 ( io_commits_info_4_debug_otherPdest_6 ),
    .io_commits_info_4_debug_fuType ( io_commits_info_4_debug_fuType ),
    .io_commits_info_4_dirtyFs ( io_commits_info_4_dirtyFs ),
    .io_commits_info_4_dirtyVs ( io_commits_info_4_dirtyVs ),
    .io_commits_info_5_walk_v ( io_commits_info_5_walk_v ),
    .io_commits_info_5_commit_v ( io_commits_info_5_commit_v ),
    .io_commits_info_5_commit_w ( io_commits_info_5_commit_w ),
    .io_commits_info_5_realDestSize ( io_commits_info_5_realDestSize ),
    .io_commits_info_5_interrupt_safe ( io_commits_info_5_interrupt_safe ),
    .io_commits_info_5_wflags ( io_commits_info_5_wflags ),
    .io_commits_info_5_fflags ( io_commits_info_5_fflags ),
    .io_commits_info_5_vxsat ( io_commits_info_5_vxsat ),
    .io_commits_info_5_isRVC ( io_commits_info_5_isRVC ),
    .io_commits_info_5_isVset ( io_commits_info_5_isVset ),
    .io_commits_info_5_isHls ( io_commits_info_5_isHls ),
    .io_commits_info_5_isVls ( io_commits_info_5_isVls ),
    .io_commits_info_5_vls ( io_commits_info_5_vls ),
    .io_commits_info_5_mmio ( io_commits_info_5_mmio ),
    .io_commits_info_5_commitType ( io_commits_info_5_commitType ),
    .io_commits_info_5_ftqIdx_flag ( io_commits_info_5_ftqIdx_flag ),
    .io_commits_info_5_ftqIdx_value ( io_commits_info_5_ftqIdx_value ),
    .io_commits_info_5_ftqOffset ( io_commits_info_5_ftqOffset ),
    .io_commits_info_5_instrSize ( io_commits_info_5_instrSize ),
    .io_commits_info_5_fpWen ( io_commits_info_5_fpWen ),
    .io_commits_info_5_rfWen ( io_commits_info_5_rfWen ),
    .io_commits_info_5_needFlush ( io_commits_info_5_needFlush ),
    .io_commits_info_5_traceBlockInPipe_itype ( io_commits_info_5_traceBlockInPipe_itype ),
    .io_commits_info_5_traceBlockInPipe_iretire ( io_commits_info_5_traceBlockInPipe_iretire ),
    .io_commits_info_5_traceBlockInPipe_ilastsize ( io_commits_info_5_traceBlockInPipe_ilastsize ),
    .io_commits_info_5_debug_pc ( io_commits_info_5_debug_pc ),
    .io_commits_info_5_debug_instr ( io_commits_info_5_debug_instr ),
    .io_commits_info_5_debug_ldest ( io_commits_info_5_debug_ldest ),
    .io_commits_info_5_debug_pdest ( io_commits_info_5_debug_pdest ),
    .io_commits_info_5_debug_otherPdest_0 ( io_commits_info_5_debug_otherPdest_0 ),
    .io_commits_info_5_debug_otherPdest_1 ( io_commits_info_5_debug_otherPdest_1 ),
    .io_commits_info_5_debug_otherPdest_2 ( io_commits_info_5_debug_otherPdest_2 ),
    .io_commits_info_5_debug_otherPdest_3 ( io_commits_info_5_debug_otherPdest_3 ),
    .io_commits_info_5_debug_otherPdest_4 ( io_commits_info_5_debug_otherPdest_4 ),
    .io_commits_info_5_debug_otherPdest_5 ( io_commits_info_5_debug_otherPdest_5 ),
    .io_commits_info_5_debug_otherPdest_6 ( io_commits_info_5_debug_otherPdest_6 ),
    .io_commits_info_5_debug_fuType ( io_commits_info_5_debug_fuType ),
    .io_commits_info_5_dirtyFs ( io_commits_info_5_dirtyFs ),
    .io_commits_info_5_dirtyVs ( io_commits_info_5_dirtyVs ),
    .io_commits_info_6_walk_v ( io_commits_info_6_walk_v ),
    .io_commits_info_6_commit_v ( io_commits_info_6_commit_v ),
    .io_commits_info_6_commit_w ( io_commits_info_6_commit_w ),
    .io_commits_info_6_realDestSize ( io_commits_info_6_realDestSize ),
    .io_commits_info_6_interrupt_safe ( io_commits_info_6_interrupt_safe ),
    .io_commits_info_6_wflags ( io_commits_info_6_wflags ),
    .io_commits_info_6_fflags ( io_commits_info_6_fflags ),
    .io_commits_info_6_vxsat ( io_commits_info_6_vxsat ),
    .io_commits_info_6_isRVC ( io_commits_info_6_isRVC ),
    .io_commits_info_6_isVset ( io_commits_info_6_isVset ),
    .io_commits_info_6_isHls ( io_commits_info_6_isHls ),
    .io_commits_info_6_isVls ( io_commits_info_6_isVls ),
    .io_commits_info_6_vls ( io_commits_info_6_vls ),
    .io_commits_info_6_mmio ( io_commits_info_6_mmio ),
    .io_commits_info_6_commitType ( io_commits_info_6_commitType ),
    .io_commits_info_6_ftqIdx_flag ( io_commits_info_6_ftqIdx_flag ),
    .io_commits_info_6_ftqIdx_value ( io_commits_info_6_ftqIdx_value ),
    .io_commits_info_6_ftqOffset ( io_commits_info_6_ftqOffset ),
    .io_commits_info_6_instrSize ( io_commits_info_6_instrSize ),
    .io_commits_info_6_fpWen ( io_commits_info_6_fpWen ),
    .io_commits_info_6_rfWen ( io_commits_info_6_rfWen ),
    .io_commits_info_6_needFlush ( io_commits_info_6_needFlush ),
    .io_commits_info_6_traceBlockInPipe_itype ( io_commits_info_6_traceBlockInPipe_itype ),
    .io_commits_info_6_traceBlockInPipe_iretire ( io_commits_info_6_traceBlockInPipe_iretire ),
    .io_commits_info_6_traceBlockInPipe_ilastsize ( io_commits_info_6_traceBlockInPipe_ilastsize ),
    .io_commits_info_6_debug_pc ( io_commits_info_6_debug_pc ),
    .io_commits_info_6_debug_instr ( io_commits_info_6_debug_instr ),
    .io_commits_info_6_debug_ldest ( io_commits_info_6_debug_ldest ),
    .io_commits_info_6_debug_pdest ( io_commits_info_6_debug_pdest ),
    .io_commits_info_6_debug_otherPdest_0 ( io_commits_info_6_debug_otherPdest_0 ),
    .io_commits_info_6_debug_otherPdest_1 ( io_commits_info_6_debug_otherPdest_1 ),
    .io_commits_info_6_debug_otherPdest_2 ( io_commits_info_6_debug_otherPdest_2 ),
    .io_commits_info_6_debug_otherPdest_3 ( io_commits_info_6_debug_otherPdest_3 ),
    .io_commits_info_6_debug_otherPdest_4 ( io_commits_info_6_debug_otherPdest_4 ),
    .io_commits_info_6_debug_otherPdest_5 ( io_commits_info_6_debug_otherPdest_5 ),
    .io_commits_info_6_debug_otherPdest_6 ( io_commits_info_6_debug_otherPdest_6 ),
    .io_commits_info_6_debug_fuType ( io_commits_info_6_debug_fuType ),
    .io_commits_info_6_dirtyFs ( io_commits_info_6_dirtyFs ),
    .io_commits_info_6_dirtyVs ( io_commits_info_6_dirtyVs ),
    .io_commits_info_7_walk_v ( io_commits_info_7_walk_v ),
    .io_commits_info_7_commit_v ( io_commits_info_7_commit_v ),
    .io_commits_info_7_commit_w ( io_commits_info_7_commit_w ),
    .io_commits_info_7_realDestSize ( io_commits_info_7_realDestSize ),
    .io_commits_info_7_interrupt_safe ( io_commits_info_7_interrupt_safe ),
    .io_commits_info_7_wflags ( io_commits_info_7_wflags ),
    .io_commits_info_7_fflags ( io_commits_info_7_fflags ),
    .io_commits_info_7_vxsat ( io_commits_info_7_vxsat ),
    .io_commits_info_7_isRVC ( io_commits_info_7_isRVC ),
    .io_commits_info_7_isVset ( io_commits_info_7_isVset ),
    .io_commits_info_7_isHls ( io_commits_info_7_isHls ),
    .io_commits_info_7_isVls ( io_commits_info_7_isVls ),
    .io_commits_info_7_vls ( io_commits_info_7_vls ),
    .io_commits_info_7_mmio ( io_commits_info_7_mmio ),
    .io_commits_info_7_commitType ( io_commits_info_7_commitType ),
    .io_commits_info_7_ftqIdx_flag ( io_commits_info_7_ftqIdx_flag ),
    .io_commits_info_7_ftqIdx_value ( io_commits_info_7_ftqIdx_value ),
    .io_commits_info_7_ftqOffset ( io_commits_info_7_ftqOffset ),
    .io_commits_info_7_instrSize ( io_commits_info_7_instrSize ),
    .io_commits_info_7_fpWen ( io_commits_info_7_fpWen ),
    .io_commits_info_7_rfWen ( io_commits_info_7_rfWen ),
    .io_commits_info_7_needFlush ( io_commits_info_7_needFlush ),
    .io_commits_info_7_traceBlockInPipe_itype ( io_commits_info_7_traceBlockInPipe_itype ),
    .io_commits_info_7_traceBlockInPipe_iretire ( io_commits_info_7_traceBlockInPipe_iretire ),
    .io_commits_info_7_traceBlockInPipe_ilastsize ( io_commits_info_7_traceBlockInPipe_ilastsize ),
    .io_commits_info_7_debug_pc ( io_commits_info_7_debug_pc ),
    .io_commits_info_7_debug_instr ( io_commits_info_7_debug_instr ),
    .io_commits_info_7_debug_ldest ( io_commits_info_7_debug_ldest ),
    .io_commits_info_7_debug_pdest ( io_commits_info_7_debug_pdest ),
    .io_commits_info_7_debug_otherPdest_0 ( io_commits_info_7_debug_otherPdest_0 ),
    .io_commits_info_7_debug_otherPdest_1 ( io_commits_info_7_debug_otherPdest_1 ),
    .io_commits_info_7_debug_otherPdest_2 ( io_commits_info_7_debug_otherPdest_2 ),
    .io_commits_info_7_debug_otherPdest_3 ( io_commits_info_7_debug_otherPdest_3 ),
    .io_commits_info_7_debug_otherPdest_4 ( io_commits_info_7_debug_otherPdest_4 ),
    .io_commits_info_7_debug_otherPdest_5 ( io_commits_info_7_debug_otherPdest_5 ),
    .io_commits_info_7_debug_otherPdest_6 ( io_commits_info_7_debug_otherPdest_6 ),
    .io_commits_info_7_debug_fuType ( io_commits_info_7_debug_fuType ),
    .io_commits_info_7_dirtyFs ( io_commits_info_7_dirtyFs ),
    .io_commits_info_7_dirtyVs ( io_commits_info_7_dirtyVs ),
    .io_commits_robIdx_0_flag ( io_commits_robIdx_0_flag ),
    .io_commits_robIdx_0_value ( io_commits_robIdx_0_value ),
    .io_commits_robIdx_1_flag ( io_commits_robIdx_1_flag ),
    .io_commits_robIdx_1_value ( io_commits_robIdx_1_value ),
    .io_commits_robIdx_2_flag ( io_commits_robIdx_2_flag ),
    .io_commits_robIdx_2_value ( io_commits_robIdx_2_value ),
    .io_commits_robIdx_3_flag ( io_commits_robIdx_3_flag ),
    .io_commits_robIdx_3_value ( io_commits_robIdx_3_value ),
    .io_commits_robIdx_4_flag ( io_commits_robIdx_4_flag ),
    .io_commits_robIdx_4_value ( io_commits_robIdx_4_value ),
    .io_commits_robIdx_5_flag ( io_commits_robIdx_5_flag ),
    .io_commits_robIdx_5_value ( io_commits_robIdx_5_value ),
    .io_commits_robIdx_6_flag ( io_commits_robIdx_6_flag ),
    .io_commits_robIdx_6_value ( io_commits_robIdx_6_value ),
    .io_commits_robIdx_7_flag ( io_commits_robIdx_7_flag ),
    .io_commits_robIdx_7_value ( io_commits_robIdx_7_value ),
    .io_trace_blockCommit ( io_trace_blockCommit ),
    .io_trace_traceCommitInfo_blocks_0_valid ( io_trace_traceCommitInfo_blocks_0_valid ),
    .io_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value ( io_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value ),
    .io_trace_traceCommitInfo_blocks_0_bits_ftqOffset ( io_trace_traceCommitInfo_blocks_0_bits_ftqOffset ),
    .io_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype ( io_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype ),
    .io_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire ( io_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire ),
    .io_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize ( io_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize ),
    .io_trace_traceCommitInfo_blocks_1_valid ( io_trace_traceCommitInfo_blocks_1_valid ),
    .io_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value ( io_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value ),
    .io_trace_traceCommitInfo_blocks_1_bits_ftqOffset ( io_trace_traceCommitInfo_blocks_1_bits_ftqOffset ),
    .io_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype ( io_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype ),
    .io_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire ( io_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire ),
    .io_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize ( io_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize ),
    .io_trace_traceCommitInfo_blocks_2_valid ( io_trace_traceCommitInfo_blocks_2_valid ),
    .io_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value ( io_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value ),
    .io_trace_traceCommitInfo_blocks_2_bits_ftqOffset ( io_trace_traceCommitInfo_blocks_2_bits_ftqOffset ),
    .io_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype ( io_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype ),
    .io_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire ( io_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire ),
    .io_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize ( io_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize ),
    .io_trace_traceCommitInfo_blocks_3_valid ( io_trace_traceCommitInfo_blocks_3_valid ),
    .io_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value ( io_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value ),
    .io_trace_traceCommitInfo_blocks_3_bits_ftqOffset ( io_trace_traceCommitInfo_blocks_3_bits_ftqOffset ),
    .io_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype ( io_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype ),
    .io_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire ( io_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire ),
    .io_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize ( io_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize ),
    .io_trace_traceCommitInfo_blocks_4_valid ( io_trace_traceCommitInfo_blocks_4_valid ),
    .io_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value ( io_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value ),
    .io_trace_traceCommitInfo_blocks_4_bits_ftqOffset ( io_trace_traceCommitInfo_blocks_4_bits_ftqOffset ),
    .io_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype ( io_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype ),
    .io_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire ( io_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire ),
    .io_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize ( io_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize ),
    .io_trace_traceCommitInfo_blocks_5_valid ( io_trace_traceCommitInfo_blocks_5_valid ),
    .io_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value ( io_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value ),
    .io_trace_traceCommitInfo_blocks_5_bits_ftqOffset ( io_trace_traceCommitInfo_blocks_5_bits_ftqOffset ),
    .io_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype ( io_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype ),
    .io_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire ( io_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire ),
    .io_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize ( io_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize ),
    .io_trace_traceCommitInfo_blocks_6_valid ( io_trace_traceCommitInfo_blocks_6_valid ),
    .io_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value ( io_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value ),
    .io_trace_traceCommitInfo_blocks_6_bits_ftqOffset ( io_trace_traceCommitInfo_blocks_6_bits_ftqOffset ),
    .io_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype ( io_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype ),
    .io_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire ( io_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire ),
    .io_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize ( io_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize ),
    .io_trace_traceCommitInfo_blocks_7_valid ( io_trace_traceCommitInfo_blocks_7_valid ),
    .io_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value ( io_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value ),
    .io_trace_traceCommitInfo_blocks_7_bits_ftqOffset ( io_trace_traceCommitInfo_blocks_7_bits_ftqOffset ),
    .io_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype ( io_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype ),
    .io_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire ( io_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire ),
    .io_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize ( io_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize ),
    .io_rabCommits_isCommit ( io_rabCommits_isCommit ),
    .io_rabCommits_commitValid_0 ( io_rabCommits_commitValid_0 ),
    .io_rabCommits_commitValid_1 ( io_rabCommits_commitValid_1 ),
    .io_rabCommits_commitValid_2 ( io_rabCommits_commitValid_2 ),
    .io_rabCommits_commitValid_3 ( io_rabCommits_commitValid_3 ),
    .io_rabCommits_commitValid_4 ( io_rabCommits_commitValid_4 ),
    .io_rabCommits_commitValid_5 ( io_rabCommits_commitValid_5 ),
    .io_rabCommits_isWalk ( io_rabCommits_isWalk ),
    .io_rabCommits_walkValid_0 ( io_rabCommits_walkValid_0 ),
    .io_rabCommits_walkValid_1 ( io_rabCommits_walkValid_1 ),
    .io_rabCommits_walkValid_2 ( io_rabCommits_walkValid_2 ),
    .io_rabCommits_walkValid_3 ( io_rabCommits_walkValid_3 ),
    .io_rabCommits_walkValid_4 ( io_rabCommits_walkValid_4 ),
    .io_rabCommits_walkValid_5 ( io_rabCommits_walkValid_5 ),
    .io_rabCommits_info_0_ldest ( io_rabCommits_info_0_ldest ),
    .io_rabCommits_info_0_pdest ( io_rabCommits_info_0_pdest ),
    .io_rabCommits_info_0_rfWen ( io_rabCommits_info_0_rfWen ),
    .io_rabCommits_info_0_fpWen ( io_rabCommits_info_0_fpWen ),
    .io_rabCommits_info_0_vecWen ( io_rabCommits_info_0_vecWen ),
    .io_rabCommits_info_0_v0Wen ( io_rabCommits_info_0_v0Wen ),
    .io_rabCommits_info_0_vlWen ( io_rabCommits_info_0_vlWen ),
    .io_rabCommits_info_0_isMove ( io_rabCommits_info_0_isMove ),
    .io_rabCommits_info_1_ldest ( io_rabCommits_info_1_ldest ),
    .io_rabCommits_info_1_pdest ( io_rabCommits_info_1_pdest ),
    .io_rabCommits_info_1_rfWen ( io_rabCommits_info_1_rfWen ),
    .io_rabCommits_info_1_fpWen ( io_rabCommits_info_1_fpWen ),
    .io_rabCommits_info_1_vecWen ( io_rabCommits_info_1_vecWen ),
    .io_rabCommits_info_1_v0Wen ( io_rabCommits_info_1_v0Wen ),
    .io_rabCommits_info_1_vlWen ( io_rabCommits_info_1_vlWen ),
    .io_rabCommits_info_1_isMove ( io_rabCommits_info_1_isMove ),
    .io_rabCommits_info_2_ldest ( io_rabCommits_info_2_ldest ),
    .io_rabCommits_info_2_pdest ( io_rabCommits_info_2_pdest ),
    .io_rabCommits_info_2_rfWen ( io_rabCommits_info_2_rfWen ),
    .io_rabCommits_info_2_fpWen ( io_rabCommits_info_2_fpWen ),
    .io_rabCommits_info_2_vecWen ( io_rabCommits_info_2_vecWen ),
    .io_rabCommits_info_2_v0Wen ( io_rabCommits_info_2_v0Wen ),
    .io_rabCommits_info_2_vlWen ( io_rabCommits_info_2_vlWen ),
    .io_rabCommits_info_2_isMove ( io_rabCommits_info_2_isMove ),
    .io_rabCommits_info_3_ldest ( io_rabCommits_info_3_ldest ),
    .io_rabCommits_info_3_pdest ( io_rabCommits_info_3_pdest ),
    .io_rabCommits_info_3_rfWen ( io_rabCommits_info_3_rfWen ),
    .io_rabCommits_info_3_fpWen ( io_rabCommits_info_3_fpWen ),
    .io_rabCommits_info_3_vecWen ( io_rabCommits_info_3_vecWen ),
    .io_rabCommits_info_3_v0Wen ( io_rabCommits_info_3_v0Wen ),
    .io_rabCommits_info_3_vlWen ( io_rabCommits_info_3_vlWen ),
    .io_rabCommits_info_3_isMove ( io_rabCommits_info_3_isMove ),
    .io_rabCommits_info_4_ldest ( io_rabCommits_info_4_ldest ),
    .io_rabCommits_info_4_pdest ( io_rabCommits_info_4_pdest ),
    .io_rabCommits_info_4_rfWen ( io_rabCommits_info_4_rfWen ),
    .io_rabCommits_info_4_fpWen ( io_rabCommits_info_4_fpWen ),
    .io_rabCommits_info_4_vecWen ( io_rabCommits_info_4_vecWen ),
    .io_rabCommits_info_4_v0Wen ( io_rabCommits_info_4_v0Wen ),
    .io_rabCommits_info_4_vlWen ( io_rabCommits_info_4_vlWen ),
    .io_rabCommits_info_4_isMove ( io_rabCommits_info_4_isMove ),
    .io_rabCommits_info_5_ldest ( io_rabCommits_info_5_ldest ),
    .io_rabCommits_info_5_pdest ( io_rabCommits_info_5_pdest ),
    .io_rabCommits_info_5_rfWen ( io_rabCommits_info_5_rfWen ),
    .io_rabCommits_info_5_fpWen ( io_rabCommits_info_5_fpWen ),
    .io_rabCommits_info_5_vecWen ( io_rabCommits_info_5_vecWen ),
    .io_rabCommits_info_5_v0Wen ( io_rabCommits_info_5_v0Wen ),
    .io_rabCommits_info_5_vlWen ( io_rabCommits_info_5_vlWen ),
    .io_rabCommits_info_5_isMove ( io_rabCommits_info_5_isMove ),
    .io_diffCommits_commitValid_0 ( io_diffCommits_commitValid_0 ),
    .io_diffCommits_commitValid_1 ( io_diffCommits_commitValid_1 ),
    .io_diffCommits_commitValid_2 ( io_diffCommits_commitValid_2 ),
    .io_diffCommits_commitValid_3 ( io_diffCommits_commitValid_3 ),
    .io_diffCommits_commitValid_4 ( io_diffCommits_commitValid_4 ),
    .io_diffCommits_commitValid_5 ( io_diffCommits_commitValid_5 ),
    .io_diffCommits_commitValid_6 ( io_diffCommits_commitValid_6 ),
    .io_diffCommits_commitValid_7 ( io_diffCommits_commitValid_7 ),
    .io_diffCommits_commitValid_8 ( io_diffCommits_commitValid_8 ),
    .io_diffCommits_commitValid_9 ( io_diffCommits_commitValid_9 ),
    .io_diffCommits_commitValid_10 ( io_diffCommits_commitValid_10 ),
    .io_diffCommits_commitValid_11 ( io_diffCommits_commitValid_11 ),
    .io_diffCommits_commitValid_12 ( io_diffCommits_commitValid_12 ),
    .io_diffCommits_commitValid_13 ( io_diffCommits_commitValid_13 ),
    .io_diffCommits_commitValid_14 ( io_diffCommits_commitValid_14 ),
    .io_diffCommits_commitValid_15 ( io_diffCommits_commitValid_15 ),
    .io_diffCommits_commitValid_16 ( io_diffCommits_commitValid_16 ),
    .io_diffCommits_commitValid_17 ( io_diffCommits_commitValid_17 ),
    .io_diffCommits_commitValid_18 ( io_diffCommits_commitValid_18 ),
    .io_diffCommits_commitValid_19 ( io_diffCommits_commitValid_19 ),
    .io_diffCommits_commitValid_20 ( io_diffCommits_commitValid_20 ),
    .io_diffCommits_commitValid_21 ( io_diffCommits_commitValid_21 ),
    .io_diffCommits_commitValid_22 ( io_diffCommits_commitValid_22 ),
    .io_diffCommits_commitValid_23 ( io_diffCommits_commitValid_23 ),
    .io_diffCommits_commitValid_24 ( io_diffCommits_commitValid_24 ),
    .io_diffCommits_commitValid_25 ( io_diffCommits_commitValid_25 ),
    .io_diffCommits_commitValid_26 ( io_diffCommits_commitValid_26 ),
    .io_diffCommits_commitValid_27 ( io_diffCommits_commitValid_27 ),
    .io_diffCommits_commitValid_28 ( io_diffCommits_commitValid_28 ),
    .io_diffCommits_commitValid_29 ( io_diffCommits_commitValid_29 ),
    .io_diffCommits_commitValid_30 ( io_diffCommits_commitValid_30 ),
    .io_diffCommits_commitValid_31 ( io_diffCommits_commitValid_31 ),
    .io_diffCommits_commitValid_32 ( io_diffCommits_commitValid_32 ),
    .io_diffCommits_commitValid_33 ( io_diffCommits_commitValid_33 ),
    .io_diffCommits_commitValid_34 ( io_diffCommits_commitValid_34 ),
    .io_diffCommits_commitValid_35 ( io_diffCommits_commitValid_35 ),
    .io_diffCommits_commitValid_36 ( io_diffCommits_commitValid_36 ),
    .io_diffCommits_commitValid_37 ( io_diffCommits_commitValid_37 ),
    .io_diffCommits_commitValid_38 ( io_diffCommits_commitValid_38 ),
    .io_diffCommits_commitValid_39 ( io_diffCommits_commitValid_39 ),
    .io_diffCommits_commitValid_40 ( io_diffCommits_commitValid_40 ),
    .io_diffCommits_commitValid_41 ( io_diffCommits_commitValid_41 ),
    .io_diffCommits_commitValid_42 ( io_diffCommits_commitValid_42 ),
    .io_diffCommits_commitValid_43 ( io_diffCommits_commitValid_43 ),
    .io_diffCommits_commitValid_44 ( io_diffCommits_commitValid_44 ),
    .io_diffCommits_commitValid_45 ( io_diffCommits_commitValid_45 ),
    .io_diffCommits_commitValid_46 ( io_diffCommits_commitValid_46 ),
    .io_diffCommits_commitValid_47 ( io_diffCommits_commitValid_47 ),
    .io_diffCommits_commitValid_48 ( io_diffCommits_commitValid_48 ),
    .io_diffCommits_commitValid_49 ( io_diffCommits_commitValid_49 ),
    .io_diffCommits_commitValid_50 ( io_diffCommits_commitValid_50 ),
    .io_diffCommits_commitValid_51 ( io_diffCommits_commitValid_51 ),
    .io_diffCommits_commitValid_52 ( io_diffCommits_commitValid_52 ),
    .io_diffCommits_commitValid_53 ( io_diffCommits_commitValid_53 ),
    .io_diffCommits_commitValid_54 ( io_diffCommits_commitValid_54 ),
    .io_diffCommits_commitValid_55 ( io_diffCommits_commitValid_55 ),
    .io_diffCommits_commitValid_56 ( io_diffCommits_commitValid_56 ),
    .io_diffCommits_commitValid_57 ( io_diffCommits_commitValid_57 ),
    .io_diffCommits_commitValid_58 ( io_diffCommits_commitValid_58 ),
    .io_diffCommits_commitValid_59 ( io_diffCommits_commitValid_59 ),
    .io_diffCommits_commitValid_60 ( io_diffCommits_commitValid_60 ),
    .io_diffCommits_commitValid_61 ( io_diffCommits_commitValid_61 ),
    .io_diffCommits_commitValid_62 ( io_diffCommits_commitValid_62 ),
    .io_diffCommits_commitValid_63 ( io_diffCommits_commitValid_63 ),
    .io_diffCommits_commitValid_64 ( io_diffCommits_commitValid_64 ),
    .io_diffCommits_commitValid_65 ( io_diffCommits_commitValid_65 ),
    .io_diffCommits_commitValid_66 ( io_diffCommits_commitValid_66 ),
    .io_diffCommits_commitValid_67 ( io_diffCommits_commitValid_67 ),
    .io_diffCommits_commitValid_68 ( io_diffCommits_commitValid_68 ),
    .io_diffCommits_commitValid_69 ( io_diffCommits_commitValid_69 ),
    .io_diffCommits_commitValid_70 ( io_diffCommits_commitValid_70 ),
    .io_diffCommits_commitValid_71 ( io_diffCommits_commitValid_71 ),
    .io_diffCommits_commitValid_72 ( io_diffCommits_commitValid_72 ),
    .io_diffCommits_commitValid_73 ( io_diffCommits_commitValid_73 ),
    .io_diffCommits_commitValid_74 ( io_diffCommits_commitValid_74 ),
    .io_diffCommits_commitValid_75 ( io_diffCommits_commitValid_75 ),
    .io_diffCommits_commitValid_76 ( io_diffCommits_commitValid_76 ),
    .io_diffCommits_commitValid_77 ( io_diffCommits_commitValid_77 ),
    .io_diffCommits_commitValid_78 ( io_diffCommits_commitValid_78 ),
    .io_diffCommits_commitValid_79 ( io_diffCommits_commitValid_79 ),
    .io_diffCommits_commitValid_80 ( io_diffCommits_commitValid_80 ),
    .io_diffCommits_commitValid_81 ( io_diffCommits_commitValid_81 ),
    .io_diffCommits_commitValid_82 ( io_diffCommits_commitValid_82 ),
    .io_diffCommits_commitValid_83 ( io_diffCommits_commitValid_83 ),
    .io_diffCommits_commitValid_84 ( io_diffCommits_commitValid_84 ),
    .io_diffCommits_commitValid_85 ( io_diffCommits_commitValid_85 ),
    .io_diffCommits_commitValid_86 ( io_diffCommits_commitValid_86 ),
    .io_diffCommits_commitValid_87 ( io_diffCommits_commitValid_87 ),
    .io_diffCommits_commitValid_88 ( io_diffCommits_commitValid_88 ),
    .io_diffCommits_commitValid_89 ( io_diffCommits_commitValid_89 ),
    .io_diffCommits_commitValid_90 ( io_diffCommits_commitValid_90 ),
    .io_diffCommits_commitValid_91 ( io_diffCommits_commitValid_91 ),
    .io_diffCommits_commitValid_92 ( io_diffCommits_commitValid_92 ),
    .io_diffCommits_commitValid_93 ( io_diffCommits_commitValid_93 ),
    .io_diffCommits_commitValid_94 ( io_diffCommits_commitValid_94 ),
    .io_diffCommits_commitValid_95 ( io_diffCommits_commitValid_95 ),
    .io_diffCommits_commitValid_96 ( io_diffCommits_commitValid_96 ),
    .io_diffCommits_commitValid_97 ( io_diffCommits_commitValid_97 ),
    .io_diffCommits_commitValid_98 ( io_diffCommits_commitValid_98 ),
    .io_diffCommits_commitValid_99 ( io_diffCommits_commitValid_99 ),
    .io_diffCommits_commitValid_100 ( io_diffCommits_commitValid_100 ),
    .io_diffCommits_commitValid_101 ( io_diffCommits_commitValid_101 ),
    .io_diffCommits_commitValid_102 ( io_diffCommits_commitValid_102 ),
    .io_diffCommits_commitValid_103 ( io_diffCommits_commitValid_103 ),
    .io_diffCommits_commitValid_104 ( io_diffCommits_commitValid_104 ),
    .io_diffCommits_commitValid_105 ( io_diffCommits_commitValid_105 ),
    .io_diffCommits_commitValid_106 ( io_diffCommits_commitValid_106 ),
    .io_diffCommits_commitValid_107 ( io_diffCommits_commitValid_107 ),
    .io_diffCommits_commitValid_108 ( io_diffCommits_commitValid_108 ),
    .io_diffCommits_commitValid_109 ( io_diffCommits_commitValid_109 ),
    .io_diffCommits_commitValid_110 ( io_diffCommits_commitValid_110 ),
    .io_diffCommits_commitValid_111 ( io_diffCommits_commitValid_111 ),
    .io_diffCommits_commitValid_112 ( io_diffCommits_commitValid_112 ),
    .io_diffCommits_commitValid_113 ( io_diffCommits_commitValid_113 ),
    .io_diffCommits_commitValid_114 ( io_diffCommits_commitValid_114 ),
    .io_diffCommits_commitValid_115 ( io_diffCommits_commitValid_115 ),
    .io_diffCommits_commitValid_116 ( io_diffCommits_commitValid_116 ),
    .io_diffCommits_commitValid_117 ( io_diffCommits_commitValid_117 ),
    .io_diffCommits_commitValid_118 ( io_diffCommits_commitValid_118 ),
    .io_diffCommits_commitValid_119 ( io_diffCommits_commitValid_119 ),
    .io_diffCommits_commitValid_120 ( io_diffCommits_commitValid_120 ),
    .io_diffCommits_commitValid_121 ( io_diffCommits_commitValid_121 ),
    .io_diffCommits_commitValid_122 ( io_diffCommits_commitValid_122 ),
    .io_diffCommits_commitValid_123 ( io_diffCommits_commitValid_123 ),
    .io_diffCommits_commitValid_124 ( io_diffCommits_commitValid_124 ),
    .io_diffCommits_commitValid_125 ( io_diffCommits_commitValid_125 ),
    .io_diffCommits_commitValid_126 ( io_diffCommits_commitValid_126 ),
    .io_diffCommits_commitValid_127 ( io_diffCommits_commitValid_127 ),
    .io_diffCommits_commitValid_128 ( io_diffCommits_commitValid_128 ),
    .io_diffCommits_commitValid_129 ( io_diffCommits_commitValid_129 ),
    .io_diffCommits_commitValid_130 ( io_diffCommits_commitValid_130 ),
    .io_diffCommits_commitValid_131 ( io_diffCommits_commitValid_131 ),
    .io_diffCommits_commitValid_132 ( io_diffCommits_commitValid_132 ),
    .io_diffCommits_commitValid_133 ( io_diffCommits_commitValid_133 ),
    .io_diffCommits_commitValid_134 ( io_diffCommits_commitValid_134 ),
    .io_diffCommits_commitValid_135 ( io_diffCommits_commitValid_135 ),
    .io_diffCommits_commitValid_136 ( io_diffCommits_commitValid_136 ),
    .io_diffCommits_commitValid_137 ( io_diffCommits_commitValid_137 ),
    .io_diffCommits_commitValid_138 ( io_diffCommits_commitValid_138 ),
    .io_diffCommits_commitValid_139 ( io_diffCommits_commitValid_139 ),
    .io_diffCommits_commitValid_140 ( io_diffCommits_commitValid_140 ),
    .io_diffCommits_commitValid_141 ( io_diffCommits_commitValid_141 ),
    .io_diffCommits_commitValid_142 ( io_diffCommits_commitValid_142 ),
    .io_diffCommits_commitValid_143 ( io_diffCommits_commitValid_143 ),
    .io_diffCommits_commitValid_144 ( io_diffCommits_commitValid_144 ),
    .io_diffCommits_commitValid_145 ( io_diffCommits_commitValid_145 ),
    .io_diffCommits_commitValid_146 ( io_diffCommits_commitValid_146 ),
    .io_diffCommits_commitValid_147 ( io_diffCommits_commitValid_147 ),
    .io_diffCommits_commitValid_148 ( io_diffCommits_commitValid_148 ),
    .io_diffCommits_commitValid_149 ( io_diffCommits_commitValid_149 ),
    .io_diffCommits_commitValid_150 ( io_diffCommits_commitValid_150 ),
    .io_diffCommits_commitValid_151 ( io_diffCommits_commitValid_151 ),
    .io_diffCommits_commitValid_152 ( io_diffCommits_commitValid_152 ),
    .io_diffCommits_commitValid_153 ( io_diffCommits_commitValid_153 ),
    .io_diffCommits_commitValid_154 ( io_diffCommits_commitValid_154 ),
    .io_diffCommits_commitValid_155 ( io_diffCommits_commitValid_155 ),
    .io_diffCommits_commitValid_156 ( io_diffCommits_commitValid_156 ),
    .io_diffCommits_commitValid_157 ( io_diffCommits_commitValid_157 ),
    .io_diffCommits_commitValid_158 ( io_diffCommits_commitValid_158 ),
    .io_diffCommits_commitValid_159 ( io_diffCommits_commitValid_159 ),
    .io_diffCommits_commitValid_160 ( io_diffCommits_commitValid_160 ),
    .io_diffCommits_commitValid_161 ( io_diffCommits_commitValid_161 ),
    .io_diffCommits_commitValid_162 ( io_diffCommits_commitValid_162 ),
    .io_diffCommits_commitValid_163 ( io_diffCommits_commitValid_163 ),
    .io_diffCommits_commitValid_164 ( io_diffCommits_commitValid_164 ),
    .io_diffCommits_commitValid_165 ( io_diffCommits_commitValid_165 ),
    .io_diffCommits_commitValid_166 ( io_diffCommits_commitValid_166 ),
    .io_diffCommits_commitValid_167 ( io_diffCommits_commitValid_167 ),
    .io_diffCommits_commitValid_168 ( io_diffCommits_commitValid_168 ),
    .io_diffCommits_commitValid_169 ( io_diffCommits_commitValid_169 ),
    .io_diffCommits_commitValid_170 ( io_diffCommits_commitValid_170 ),
    .io_diffCommits_commitValid_171 ( io_diffCommits_commitValid_171 ),
    .io_diffCommits_commitValid_172 ( io_diffCommits_commitValid_172 ),
    .io_diffCommits_commitValid_173 ( io_diffCommits_commitValid_173 ),
    .io_diffCommits_commitValid_174 ( io_diffCommits_commitValid_174 ),
    .io_diffCommits_commitValid_175 ( io_diffCommits_commitValid_175 ),
    .io_diffCommits_commitValid_176 ( io_diffCommits_commitValid_176 ),
    .io_diffCommits_commitValid_177 ( io_diffCommits_commitValid_177 ),
    .io_diffCommits_commitValid_178 ( io_diffCommits_commitValid_178 ),
    .io_diffCommits_commitValid_179 ( io_diffCommits_commitValid_179 ),
    .io_diffCommits_commitValid_180 ( io_diffCommits_commitValid_180 ),
    .io_diffCommits_commitValid_181 ( io_diffCommits_commitValid_181 ),
    .io_diffCommits_commitValid_182 ( io_diffCommits_commitValid_182 ),
    .io_diffCommits_commitValid_183 ( io_diffCommits_commitValid_183 ),
    .io_diffCommits_commitValid_184 ( io_diffCommits_commitValid_184 ),
    .io_diffCommits_commitValid_185 ( io_diffCommits_commitValid_185 ),
    .io_diffCommits_commitValid_186 ( io_diffCommits_commitValid_186 ),
    .io_diffCommits_commitValid_187 ( io_diffCommits_commitValid_187 ),
    .io_diffCommits_commitValid_188 ( io_diffCommits_commitValid_188 ),
    .io_diffCommits_commitValid_189 ( io_diffCommits_commitValid_189 ),
    .io_diffCommits_commitValid_190 ( io_diffCommits_commitValid_190 ),
    .io_diffCommits_commitValid_191 ( io_diffCommits_commitValid_191 ),
    .io_diffCommits_commitValid_192 ( io_diffCommits_commitValid_192 ),
    .io_diffCommits_commitValid_193 ( io_diffCommits_commitValid_193 ),
    .io_diffCommits_commitValid_194 ( io_diffCommits_commitValid_194 ),
    .io_diffCommits_commitValid_195 ( io_diffCommits_commitValid_195 ),
    .io_diffCommits_commitValid_196 ( io_diffCommits_commitValid_196 ),
    .io_diffCommits_commitValid_197 ( io_diffCommits_commitValid_197 ),
    .io_diffCommits_commitValid_198 ( io_diffCommits_commitValid_198 ),
    .io_diffCommits_commitValid_199 ( io_diffCommits_commitValid_199 ),
    .io_diffCommits_commitValid_200 ( io_diffCommits_commitValid_200 ),
    .io_diffCommits_commitValid_201 ( io_diffCommits_commitValid_201 ),
    .io_diffCommits_commitValid_202 ( io_diffCommits_commitValid_202 ),
    .io_diffCommits_commitValid_203 ( io_diffCommits_commitValid_203 ),
    .io_diffCommits_commitValid_204 ( io_diffCommits_commitValid_204 ),
    .io_diffCommits_commitValid_205 ( io_diffCommits_commitValid_205 ),
    .io_diffCommits_commitValid_206 ( io_diffCommits_commitValid_206 ),
    .io_diffCommits_commitValid_207 ( io_diffCommits_commitValid_207 ),
    .io_diffCommits_commitValid_208 ( io_diffCommits_commitValid_208 ),
    .io_diffCommits_commitValid_209 ( io_diffCommits_commitValid_209 ),
    .io_diffCommits_commitValid_210 ( io_diffCommits_commitValid_210 ),
    .io_diffCommits_commitValid_211 ( io_diffCommits_commitValid_211 ),
    .io_diffCommits_commitValid_212 ( io_diffCommits_commitValid_212 ),
    .io_diffCommits_commitValid_213 ( io_diffCommits_commitValid_213 ),
    .io_diffCommits_commitValid_214 ( io_diffCommits_commitValid_214 ),
    .io_diffCommits_commitValid_215 ( io_diffCommits_commitValid_215 ),
    .io_diffCommits_commitValid_216 ( io_diffCommits_commitValid_216 ),
    .io_diffCommits_commitValid_217 ( io_diffCommits_commitValid_217 ),
    .io_diffCommits_commitValid_218 ( io_diffCommits_commitValid_218 ),
    .io_diffCommits_commitValid_219 ( io_diffCommits_commitValid_219 ),
    .io_diffCommits_commitValid_220 ( io_diffCommits_commitValid_220 ),
    .io_diffCommits_commitValid_221 ( io_diffCommits_commitValid_221 ),
    .io_diffCommits_commitValid_222 ( io_diffCommits_commitValid_222 ),
    .io_diffCommits_commitValid_223 ( io_diffCommits_commitValid_223 ),
    .io_diffCommits_commitValid_224 ( io_diffCommits_commitValid_224 ),
    .io_diffCommits_commitValid_225 ( io_diffCommits_commitValid_225 ),
    .io_diffCommits_commitValid_226 ( io_diffCommits_commitValid_226 ),
    .io_diffCommits_commitValid_227 ( io_diffCommits_commitValid_227 ),
    .io_diffCommits_commitValid_228 ( io_diffCommits_commitValid_228 ),
    .io_diffCommits_commitValid_229 ( io_diffCommits_commitValid_229 ),
    .io_diffCommits_commitValid_230 ( io_diffCommits_commitValid_230 ),
    .io_diffCommits_commitValid_231 ( io_diffCommits_commitValid_231 ),
    .io_diffCommits_commitValid_232 ( io_diffCommits_commitValid_232 ),
    .io_diffCommits_commitValid_233 ( io_diffCommits_commitValid_233 ),
    .io_diffCommits_commitValid_234 ( io_diffCommits_commitValid_234 ),
    .io_diffCommits_commitValid_235 ( io_diffCommits_commitValid_235 ),
    .io_diffCommits_commitValid_236 ( io_diffCommits_commitValid_236 ),
    .io_diffCommits_commitValid_237 ( io_diffCommits_commitValid_237 ),
    .io_diffCommits_commitValid_238 ( io_diffCommits_commitValid_238 ),
    .io_diffCommits_commitValid_239 ( io_diffCommits_commitValid_239 ),
    .io_diffCommits_commitValid_240 ( io_diffCommits_commitValid_240 ),
    .io_diffCommits_commitValid_241 ( io_diffCommits_commitValid_241 ),
    .io_diffCommits_commitValid_242 ( io_diffCommits_commitValid_242 ),
    .io_diffCommits_commitValid_243 ( io_diffCommits_commitValid_243 ),
    .io_diffCommits_commitValid_244 ( io_diffCommits_commitValid_244 ),
    .io_diffCommits_commitValid_245 ( io_diffCommits_commitValid_245 ),
    .io_diffCommits_commitValid_246 ( io_diffCommits_commitValid_246 ),
    .io_diffCommits_commitValid_247 ( io_diffCommits_commitValid_247 ),
    .io_diffCommits_commitValid_248 ( io_diffCommits_commitValid_248 ),
    .io_diffCommits_commitValid_249 ( io_diffCommits_commitValid_249 ),
    .io_diffCommits_commitValid_250 ( io_diffCommits_commitValid_250 ),
    .io_diffCommits_commitValid_251 ( io_diffCommits_commitValid_251 ),
    .io_diffCommits_commitValid_252 ( io_diffCommits_commitValid_252 ),
    .io_diffCommits_commitValid_253 ( io_diffCommits_commitValid_253 ),
    .io_diffCommits_commitValid_254 ( io_diffCommits_commitValid_254 ),
    .io_diffCommits_info_0_ldest ( io_diffCommits_info_0_ldest ),
    .io_diffCommits_info_0_pdest ( io_diffCommits_info_0_pdest ),
    .io_diffCommits_info_0_rfWen ( io_diffCommits_info_0_rfWen ),
    .io_diffCommits_info_0_fpWen ( io_diffCommits_info_0_fpWen ),
    .io_diffCommits_info_0_vecWen ( io_diffCommits_info_0_vecWen ),
    .io_diffCommits_info_0_v0Wen ( io_diffCommits_info_0_v0Wen ),
    .io_diffCommits_info_0_vlWen ( io_diffCommits_info_0_vlWen ),
    .io_diffCommits_info_1_ldest ( io_diffCommits_info_1_ldest ),
    .io_diffCommits_info_1_pdest ( io_diffCommits_info_1_pdest ),
    .io_diffCommits_info_1_rfWen ( io_diffCommits_info_1_rfWen ),
    .io_diffCommits_info_1_fpWen ( io_diffCommits_info_1_fpWen ),
    .io_diffCommits_info_1_vecWen ( io_diffCommits_info_1_vecWen ),
    .io_diffCommits_info_1_v0Wen ( io_diffCommits_info_1_v0Wen ),
    .io_diffCommits_info_1_vlWen ( io_diffCommits_info_1_vlWen ),
    .io_diffCommits_info_2_ldest ( io_diffCommits_info_2_ldest ),
    .io_diffCommits_info_2_pdest ( io_diffCommits_info_2_pdest ),
    .io_diffCommits_info_2_rfWen ( io_diffCommits_info_2_rfWen ),
    .io_diffCommits_info_2_fpWen ( io_diffCommits_info_2_fpWen ),
    .io_diffCommits_info_2_vecWen ( io_diffCommits_info_2_vecWen ),
    .io_diffCommits_info_2_v0Wen ( io_diffCommits_info_2_v0Wen ),
    .io_diffCommits_info_2_vlWen ( io_diffCommits_info_2_vlWen ),
    .io_diffCommits_info_3_ldest ( io_diffCommits_info_3_ldest ),
    .io_diffCommits_info_3_pdest ( io_diffCommits_info_3_pdest ),
    .io_diffCommits_info_3_rfWen ( io_diffCommits_info_3_rfWen ),
    .io_diffCommits_info_3_fpWen ( io_diffCommits_info_3_fpWen ),
    .io_diffCommits_info_3_vecWen ( io_diffCommits_info_3_vecWen ),
    .io_diffCommits_info_3_v0Wen ( io_diffCommits_info_3_v0Wen ),
    .io_diffCommits_info_3_vlWen ( io_diffCommits_info_3_vlWen ),
    .io_diffCommits_info_4_ldest ( io_diffCommits_info_4_ldest ),
    .io_diffCommits_info_4_pdest ( io_diffCommits_info_4_pdest ),
    .io_diffCommits_info_4_rfWen ( io_diffCommits_info_4_rfWen ),
    .io_diffCommits_info_4_fpWen ( io_diffCommits_info_4_fpWen ),
    .io_diffCommits_info_4_vecWen ( io_diffCommits_info_4_vecWen ),
    .io_diffCommits_info_4_v0Wen ( io_diffCommits_info_4_v0Wen ),
    .io_diffCommits_info_4_vlWen ( io_diffCommits_info_4_vlWen ),
    .io_diffCommits_info_5_ldest ( io_diffCommits_info_5_ldest ),
    .io_diffCommits_info_5_pdest ( io_diffCommits_info_5_pdest ),
    .io_diffCommits_info_5_rfWen ( io_diffCommits_info_5_rfWen ),
    .io_diffCommits_info_5_fpWen ( io_diffCommits_info_5_fpWen ),
    .io_diffCommits_info_5_vecWen ( io_diffCommits_info_5_vecWen ),
    .io_diffCommits_info_5_v0Wen ( io_diffCommits_info_5_v0Wen ),
    .io_diffCommits_info_5_vlWen ( io_diffCommits_info_5_vlWen ),
    .io_diffCommits_info_6_ldest ( io_diffCommits_info_6_ldest ),
    .io_diffCommits_info_6_pdest ( io_diffCommits_info_6_pdest ),
    .io_diffCommits_info_6_rfWen ( io_diffCommits_info_6_rfWen ),
    .io_diffCommits_info_6_fpWen ( io_diffCommits_info_6_fpWen ),
    .io_diffCommits_info_6_vecWen ( io_diffCommits_info_6_vecWen ),
    .io_diffCommits_info_6_v0Wen ( io_diffCommits_info_6_v0Wen ),
    .io_diffCommits_info_6_vlWen ( io_diffCommits_info_6_vlWen ),
    .io_diffCommits_info_7_ldest ( io_diffCommits_info_7_ldest ),
    .io_diffCommits_info_7_pdest ( io_diffCommits_info_7_pdest ),
    .io_diffCommits_info_7_rfWen ( io_diffCommits_info_7_rfWen ),
    .io_diffCommits_info_7_fpWen ( io_diffCommits_info_7_fpWen ),
    .io_diffCommits_info_7_vecWen ( io_diffCommits_info_7_vecWen ),
    .io_diffCommits_info_7_v0Wen ( io_diffCommits_info_7_v0Wen ),
    .io_diffCommits_info_7_vlWen ( io_diffCommits_info_7_vlWen ),
    .io_diffCommits_info_8_ldest ( io_diffCommits_info_8_ldest ),
    .io_diffCommits_info_8_pdest ( io_diffCommits_info_8_pdest ),
    .io_diffCommits_info_8_rfWen ( io_diffCommits_info_8_rfWen ),
    .io_diffCommits_info_8_fpWen ( io_diffCommits_info_8_fpWen ),
    .io_diffCommits_info_8_vecWen ( io_diffCommits_info_8_vecWen ),
    .io_diffCommits_info_8_v0Wen ( io_diffCommits_info_8_v0Wen ),
    .io_diffCommits_info_8_vlWen ( io_diffCommits_info_8_vlWen ),
    .io_diffCommits_info_9_ldest ( io_diffCommits_info_9_ldest ),
    .io_diffCommits_info_9_pdest ( io_diffCommits_info_9_pdest ),
    .io_diffCommits_info_9_rfWen ( io_diffCommits_info_9_rfWen ),
    .io_diffCommits_info_9_fpWen ( io_diffCommits_info_9_fpWen ),
    .io_diffCommits_info_9_vecWen ( io_diffCommits_info_9_vecWen ),
    .io_diffCommits_info_9_v0Wen ( io_diffCommits_info_9_v0Wen ),
    .io_diffCommits_info_9_vlWen ( io_diffCommits_info_9_vlWen ),
    .io_diffCommits_info_10_ldest ( io_diffCommits_info_10_ldest ),
    .io_diffCommits_info_10_pdest ( io_diffCommits_info_10_pdest ),
    .io_diffCommits_info_10_rfWen ( io_diffCommits_info_10_rfWen ),
    .io_diffCommits_info_10_fpWen ( io_diffCommits_info_10_fpWen ),
    .io_diffCommits_info_10_vecWen ( io_diffCommits_info_10_vecWen ),
    .io_diffCommits_info_10_v0Wen ( io_diffCommits_info_10_v0Wen ),
    .io_diffCommits_info_10_vlWen ( io_diffCommits_info_10_vlWen ),
    .io_diffCommits_info_11_ldest ( io_diffCommits_info_11_ldest ),
    .io_diffCommits_info_11_pdest ( io_diffCommits_info_11_pdest ),
    .io_diffCommits_info_11_rfWen ( io_diffCommits_info_11_rfWen ),
    .io_diffCommits_info_11_fpWen ( io_diffCommits_info_11_fpWen ),
    .io_diffCommits_info_11_vecWen ( io_diffCommits_info_11_vecWen ),
    .io_diffCommits_info_11_v0Wen ( io_diffCommits_info_11_v0Wen ),
    .io_diffCommits_info_11_vlWen ( io_diffCommits_info_11_vlWen ),
    .io_diffCommits_info_12_ldest ( io_diffCommits_info_12_ldest ),
    .io_diffCommits_info_12_pdest ( io_diffCommits_info_12_pdest ),
    .io_diffCommits_info_12_rfWen ( io_diffCommits_info_12_rfWen ),
    .io_diffCommits_info_12_fpWen ( io_diffCommits_info_12_fpWen ),
    .io_diffCommits_info_12_vecWen ( io_diffCommits_info_12_vecWen ),
    .io_diffCommits_info_12_v0Wen ( io_diffCommits_info_12_v0Wen ),
    .io_diffCommits_info_12_vlWen ( io_diffCommits_info_12_vlWen ),
    .io_diffCommits_info_13_ldest ( io_diffCommits_info_13_ldest ),
    .io_diffCommits_info_13_pdest ( io_diffCommits_info_13_pdest ),
    .io_diffCommits_info_13_rfWen ( io_diffCommits_info_13_rfWen ),
    .io_diffCommits_info_13_fpWen ( io_diffCommits_info_13_fpWen ),
    .io_diffCommits_info_13_vecWen ( io_diffCommits_info_13_vecWen ),
    .io_diffCommits_info_13_v0Wen ( io_diffCommits_info_13_v0Wen ),
    .io_diffCommits_info_13_vlWen ( io_diffCommits_info_13_vlWen ),
    .io_diffCommits_info_14_ldest ( io_diffCommits_info_14_ldest ),
    .io_diffCommits_info_14_pdest ( io_diffCommits_info_14_pdest ),
    .io_diffCommits_info_14_rfWen ( io_diffCommits_info_14_rfWen ),
    .io_diffCommits_info_14_fpWen ( io_diffCommits_info_14_fpWen ),
    .io_diffCommits_info_14_vecWen ( io_diffCommits_info_14_vecWen ),
    .io_diffCommits_info_14_v0Wen ( io_diffCommits_info_14_v0Wen ),
    .io_diffCommits_info_14_vlWen ( io_diffCommits_info_14_vlWen ),
    .io_diffCommits_info_15_ldest ( io_diffCommits_info_15_ldest ),
    .io_diffCommits_info_15_pdest ( io_diffCommits_info_15_pdest ),
    .io_diffCommits_info_15_rfWen ( io_diffCommits_info_15_rfWen ),
    .io_diffCommits_info_15_fpWen ( io_diffCommits_info_15_fpWen ),
    .io_diffCommits_info_15_vecWen ( io_diffCommits_info_15_vecWen ),
    .io_diffCommits_info_15_v0Wen ( io_diffCommits_info_15_v0Wen ),
    .io_diffCommits_info_15_vlWen ( io_diffCommits_info_15_vlWen ),
    .io_diffCommits_info_16_ldest ( io_diffCommits_info_16_ldest ),
    .io_diffCommits_info_16_pdest ( io_diffCommits_info_16_pdest ),
    .io_diffCommits_info_16_rfWen ( io_diffCommits_info_16_rfWen ),
    .io_diffCommits_info_16_fpWen ( io_diffCommits_info_16_fpWen ),
    .io_diffCommits_info_16_vecWen ( io_diffCommits_info_16_vecWen ),
    .io_diffCommits_info_16_v0Wen ( io_diffCommits_info_16_v0Wen ),
    .io_diffCommits_info_16_vlWen ( io_diffCommits_info_16_vlWen ),
    .io_diffCommits_info_17_ldest ( io_diffCommits_info_17_ldest ),
    .io_diffCommits_info_17_pdest ( io_diffCommits_info_17_pdest ),
    .io_diffCommits_info_17_rfWen ( io_diffCommits_info_17_rfWen ),
    .io_diffCommits_info_17_fpWen ( io_diffCommits_info_17_fpWen ),
    .io_diffCommits_info_17_vecWen ( io_diffCommits_info_17_vecWen ),
    .io_diffCommits_info_17_v0Wen ( io_diffCommits_info_17_v0Wen ),
    .io_diffCommits_info_17_vlWen ( io_diffCommits_info_17_vlWen ),
    .io_diffCommits_info_18_ldest ( io_diffCommits_info_18_ldest ),
    .io_diffCommits_info_18_pdest ( io_diffCommits_info_18_pdest ),
    .io_diffCommits_info_18_rfWen ( io_diffCommits_info_18_rfWen ),
    .io_diffCommits_info_18_fpWen ( io_diffCommits_info_18_fpWen ),
    .io_diffCommits_info_18_vecWen ( io_diffCommits_info_18_vecWen ),
    .io_diffCommits_info_18_v0Wen ( io_diffCommits_info_18_v0Wen ),
    .io_diffCommits_info_18_vlWen ( io_diffCommits_info_18_vlWen ),
    .io_diffCommits_info_19_ldest ( io_diffCommits_info_19_ldest ),
    .io_diffCommits_info_19_pdest ( io_diffCommits_info_19_pdest ),
    .io_diffCommits_info_19_rfWen ( io_diffCommits_info_19_rfWen ),
    .io_diffCommits_info_19_fpWen ( io_diffCommits_info_19_fpWen ),
    .io_diffCommits_info_19_vecWen ( io_diffCommits_info_19_vecWen ),
    .io_diffCommits_info_19_v0Wen ( io_diffCommits_info_19_v0Wen ),
    .io_diffCommits_info_19_vlWen ( io_diffCommits_info_19_vlWen ),
    .io_diffCommits_info_20_ldest ( io_diffCommits_info_20_ldest ),
    .io_diffCommits_info_20_pdest ( io_diffCommits_info_20_pdest ),
    .io_diffCommits_info_20_rfWen ( io_diffCommits_info_20_rfWen ),
    .io_diffCommits_info_20_fpWen ( io_diffCommits_info_20_fpWen ),
    .io_diffCommits_info_20_vecWen ( io_diffCommits_info_20_vecWen ),
    .io_diffCommits_info_20_v0Wen ( io_diffCommits_info_20_v0Wen ),
    .io_diffCommits_info_20_vlWen ( io_diffCommits_info_20_vlWen ),
    .io_diffCommits_info_21_ldest ( io_diffCommits_info_21_ldest ),
    .io_diffCommits_info_21_pdest ( io_diffCommits_info_21_pdest ),
    .io_diffCommits_info_21_rfWen ( io_diffCommits_info_21_rfWen ),
    .io_diffCommits_info_21_fpWen ( io_diffCommits_info_21_fpWen ),
    .io_diffCommits_info_21_vecWen ( io_diffCommits_info_21_vecWen ),
    .io_diffCommits_info_21_v0Wen ( io_diffCommits_info_21_v0Wen ),
    .io_diffCommits_info_21_vlWen ( io_diffCommits_info_21_vlWen ),
    .io_diffCommits_info_22_ldest ( io_diffCommits_info_22_ldest ),
    .io_diffCommits_info_22_pdest ( io_diffCommits_info_22_pdest ),
    .io_diffCommits_info_22_rfWen ( io_diffCommits_info_22_rfWen ),
    .io_diffCommits_info_22_fpWen ( io_diffCommits_info_22_fpWen ),
    .io_diffCommits_info_22_vecWen ( io_diffCommits_info_22_vecWen ),
    .io_diffCommits_info_22_v0Wen ( io_diffCommits_info_22_v0Wen ),
    .io_diffCommits_info_22_vlWen ( io_diffCommits_info_22_vlWen ),
    .io_diffCommits_info_23_ldest ( io_diffCommits_info_23_ldest ),
    .io_diffCommits_info_23_pdest ( io_diffCommits_info_23_pdest ),
    .io_diffCommits_info_23_rfWen ( io_diffCommits_info_23_rfWen ),
    .io_diffCommits_info_23_fpWen ( io_diffCommits_info_23_fpWen ),
    .io_diffCommits_info_23_vecWen ( io_diffCommits_info_23_vecWen ),
    .io_diffCommits_info_23_v0Wen ( io_diffCommits_info_23_v0Wen ),
    .io_diffCommits_info_23_vlWen ( io_diffCommits_info_23_vlWen ),
    .io_diffCommits_info_24_ldest ( io_diffCommits_info_24_ldest ),
    .io_diffCommits_info_24_pdest ( io_diffCommits_info_24_pdest ),
    .io_diffCommits_info_24_rfWen ( io_diffCommits_info_24_rfWen ),
    .io_diffCommits_info_24_fpWen ( io_diffCommits_info_24_fpWen ),
    .io_diffCommits_info_24_vecWen ( io_diffCommits_info_24_vecWen ),
    .io_diffCommits_info_24_v0Wen ( io_diffCommits_info_24_v0Wen ),
    .io_diffCommits_info_24_vlWen ( io_diffCommits_info_24_vlWen ),
    .io_diffCommits_info_25_ldest ( io_diffCommits_info_25_ldest ),
    .io_diffCommits_info_25_pdest ( io_diffCommits_info_25_pdest ),
    .io_diffCommits_info_25_rfWen ( io_diffCommits_info_25_rfWen ),
    .io_diffCommits_info_25_fpWen ( io_diffCommits_info_25_fpWen ),
    .io_diffCommits_info_25_vecWen ( io_diffCommits_info_25_vecWen ),
    .io_diffCommits_info_25_v0Wen ( io_diffCommits_info_25_v0Wen ),
    .io_diffCommits_info_25_vlWen ( io_diffCommits_info_25_vlWen ),
    .io_diffCommits_info_26_ldest ( io_diffCommits_info_26_ldest ),
    .io_diffCommits_info_26_pdest ( io_diffCommits_info_26_pdest ),
    .io_diffCommits_info_26_rfWen ( io_diffCommits_info_26_rfWen ),
    .io_diffCommits_info_26_fpWen ( io_diffCommits_info_26_fpWen ),
    .io_diffCommits_info_26_vecWen ( io_diffCommits_info_26_vecWen ),
    .io_diffCommits_info_26_v0Wen ( io_diffCommits_info_26_v0Wen ),
    .io_diffCommits_info_26_vlWen ( io_diffCommits_info_26_vlWen ),
    .io_diffCommits_info_27_ldest ( io_diffCommits_info_27_ldest ),
    .io_diffCommits_info_27_pdest ( io_diffCommits_info_27_pdest ),
    .io_diffCommits_info_27_rfWen ( io_diffCommits_info_27_rfWen ),
    .io_diffCommits_info_27_fpWen ( io_diffCommits_info_27_fpWen ),
    .io_diffCommits_info_27_vecWen ( io_diffCommits_info_27_vecWen ),
    .io_diffCommits_info_27_v0Wen ( io_diffCommits_info_27_v0Wen ),
    .io_diffCommits_info_27_vlWen ( io_diffCommits_info_27_vlWen ),
    .io_diffCommits_info_28_ldest ( io_diffCommits_info_28_ldest ),
    .io_diffCommits_info_28_pdest ( io_diffCommits_info_28_pdest ),
    .io_diffCommits_info_28_rfWen ( io_diffCommits_info_28_rfWen ),
    .io_diffCommits_info_28_fpWen ( io_diffCommits_info_28_fpWen ),
    .io_diffCommits_info_28_vecWen ( io_diffCommits_info_28_vecWen ),
    .io_diffCommits_info_28_v0Wen ( io_diffCommits_info_28_v0Wen ),
    .io_diffCommits_info_28_vlWen ( io_diffCommits_info_28_vlWen ),
    .io_diffCommits_info_29_ldest ( io_diffCommits_info_29_ldest ),
    .io_diffCommits_info_29_pdest ( io_diffCommits_info_29_pdest ),
    .io_diffCommits_info_29_rfWen ( io_diffCommits_info_29_rfWen ),
    .io_diffCommits_info_29_fpWen ( io_diffCommits_info_29_fpWen ),
    .io_diffCommits_info_29_vecWen ( io_diffCommits_info_29_vecWen ),
    .io_diffCommits_info_29_v0Wen ( io_diffCommits_info_29_v0Wen ),
    .io_diffCommits_info_29_vlWen ( io_diffCommits_info_29_vlWen ),
    .io_diffCommits_info_30_ldest ( io_diffCommits_info_30_ldest ),
    .io_diffCommits_info_30_pdest ( io_diffCommits_info_30_pdest ),
    .io_diffCommits_info_30_rfWen ( io_diffCommits_info_30_rfWen ),
    .io_diffCommits_info_30_fpWen ( io_diffCommits_info_30_fpWen ),
    .io_diffCommits_info_30_vecWen ( io_diffCommits_info_30_vecWen ),
    .io_diffCommits_info_30_v0Wen ( io_diffCommits_info_30_v0Wen ),
    .io_diffCommits_info_30_vlWen ( io_diffCommits_info_30_vlWen ),
    .io_diffCommits_info_31_ldest ( io_diffCommits_info_31_ldest ),
    .io_diffCommits_info_31_pdest ( io_diffCommits_info_31_pdest ),
    .io_diffCommits_info_31_rfWen ( io_diffCommits_info_31_rfWen ),
    .io_diffCommits_info_31_fpWen ( io_diffCommits_info_31_fpWen ),
    .io_diffCommits_info_31_vecWen ( io_diffCommits_info_31_vecWen ),
    .io_diffCommits_info_31_v0Wen ( io_diffCommits_info_31_v0Wen ),
    .io_diffCommits_info_31_vlWen ( io_diffCommits_info_31_vlWen ),
    .io_diffCommits_info_32_ldest ( io_diffCommits_info_32_ldest ),
    .io_diffCommits_info_32_pdest ( io_diffCommits_info_32_pdest ),
    .io_diffCommits_info_32_rfWen ( io_diffCommits_info_32_rfWen ),
    .io_diffCommits_info_32_fpWen ( io_diffCommits_info_32_fpWen ),
    .io_diffCommits_info_32_vecWen ( io_diffCommits_info_32_vecWen ),
    .io_diffCommits_info_32_v0Wen ( io_diffCommits_info_32_v0Wen ),
    .io_diffCommits_info_32_vlWen ( io_diffCommits_info_32_vlWen ),
    .io_diffCommits_info_33_ldest ( io_diffCommits_info_33_ldest ),
    .io_diffCommits_info_33_pdest ( io_diffCommits_info_33_pdest ),
    .io_diffCommits_info_33_rfWen ( io_diffCommits_info_33_rfWen ),
    .io_diffCommits_info_33_fpWen ( io_diffCommits_info_33_fpWen ),
    .io_diffCommits_info_33_vecWen ( io_diffCommits_info_33_vecWen ),
    .io_diffCommits_info_33_v0Wen ( io_diffCommits_info_33_v0Wen ),
    .io_diffCommits_info_33_vlWen ( io_diffCommits_info_33_vlWen ),
    .io_diffCommits_info_34_ldest ( io_diffCommits_info_34_ldest ),
    .io_diffCommits_info_34_pdest ( io_diffCommits_info_34_pdest ),
    .io_diffCommits_info_34_rfWen ( io_diffCommits_info_34_rfWen ),
    .io_diffCommits_info_34_fpWen ( io_diffCommits_info_34_fpWen ),
    .io_diffCommits_info_34_vecWen ( io_diffCommits_info_34_vecWen ),
    .io_diffCommits_info_34_v0Wen ( io_diffCommits_info_34_v0Wen ),
    .io_diffCommits_info_34_vlWen ( io_diffCommits_info_34_vlWen ),
    .io_diffCommits_info_35_ldest ( io_diffCommits_info_35_ldest ),
    .io_diffCommits_info_35_pdest ( io_diffCommits_info_35_pdest ),
    .io_diffCommits_info_35_rfWen ( io_diffCommits_info_35_rfWen ),
    .io_diffCommits_info_35_fpWen ( io_diffCommits_info_35_fpWen ),
    .io_diffCommits_info_35_vecWen ( io_diffCommits_info_35_vecWen ),
    .io_diffCommits_info_35_v0Wen ( io_diffCommits_info_35_v0Wen ),
    .io_diffCommits_info_35_vlWen ( io_diffCommits_info_35_vlWen ),
    .io_diffCommits_info_36_ldest ( io_diffCommits_info_36_ldest ),
    .io_diffCommits_info_36_pdest ( io_diffCommits_info_36_pdest ),
    .io_diffCommits_info_36_rfWen ( io_diffCommits_info_36_rfWen ),
    .io_diffCommits_info_36_fpWen ( io_diffCommits_info_36_fpWen ),
    .io_diffCommits_info_36_vecWen ( io_diffCommits_info_36_vecWen ),
    .io_diffCommits_info_36_v0Wen ( io_diffCommits_info_36_v0Wen ),
    .io_diffCommits_info_36_vlWen ( io_diffCommits_info_36_vlWen ),
    .io_diffCommits_info_37_ldest ( io_diffCommits_info_37_ldest ),
    .io_diffCommits_info_37_pdest ( io_diffCommits_info_37_pdest ),
    .io_diffCommits_info_37_rfWen ( io_diffCommits_info_37_rfWen ),
    .io_diffCommits_info_37_fpWen ( io_diffCommits_info_37_fpWen ),
    .io_diffCommits_info_37_vecWen ( io_diffCommits_info_37_vecWen ),
    .io_diffCommits_info_37_v0Wen ( io_diffCommits_info_37_v0Wen ),
    .io_diffCommits_info_37_vlWen ( io_diffCommits_info_37_vlWen ),
    .io_diffCommits_info_38_ldest ( io_diffCommits_info_38_ldest ),
    .io_diffCommits_info_38_pdest ( io_diffCommits_info_38_pdest ),
    .io_diffCommits_info_38_rfWen ( io_diffCommits_info_38_rfWen ),
    .io_diffCommits_info_38_fpWen ( io_diffCommits_info_38_fpWen ),
    .io_diffCommits_info_38_vecWen ( io_diffCommits_info_38_vecWen ),
    .io_diffCommits_info_38_v0Wen ( io_diffCommits_info_38_v0Wen ),
    .io_diffCommits_info_38_vlWen ( io_diffCommits_info_38_vlWen ),
    .io_diffCommits_info_39_ldest ( io_diffCommits_info_39_ldest ),
    .io_diffCommits_info_39_pdest ( io_diffCommits_info_39_pdest ),
    .io_diffCommits_info_39_rfWen ( io_diffCommits_info_39_rfWen ),
    .io_diffCommits_info_39_fpWen ( io_diffCommits_info_39_fpWen ),
    .io_diffCommits_info_39_vecWen ( io_diffCommits_info_39_vecWen ),
    .io_diffCommits_info_39_v0Wen ( io_diffCommits_info_39_v0Wen ),
    .io_diffCommits_info_39_vlWen ( io_diffCommits_info_39_vlWen ),
    .io_diffCommits_info_40_ldest ( io_diffCommits_info_40_ldest ),
    .io_diffCommits_info_40_pdest ( io_diffCommits_info_40_pdest ),
    .io_diffCommits_info_40_rfWen ( io_diffCommits_info_40_rfWen ),
    .io_diffCommits_info_40_fpWen ( io_diffCommits_info_40_fpWen ),
    .io_diffCommits_info_40_vecWen ( io_diffCommits_info_40_vecWen ),
    .io_diffCommits_info_40_v0Wen ( io_diffCommits_info_40_v0Wen ),
    .io_diffCommits_info_40_vlWen ( io_diffCommits_info_40_vlWen ),
    .io_diffCommits_info_41_ldest ( io_diffCommits_info_41_ldest ),
    .io_diffCommits_info_41_pdest ( io_diffCommits_info_41_pdest ),
    .io_diffCommits_info_41_rfWen ( io_diffCommits_info_41_rfWen ),
    .io_diffCommits_info_41_fpWen ( io_diffCommits_info_41_fpWen ),
    .io_diffCommits_info_41_vecWen ( io_diffCommits_info_41_vecWen ),
    .io_diffCommits_info_41_v0Wen ( io_diffCommits_info_41_v0Wen ),
    .io_diffCommits_info_41_vlWen ( io_diffCommits_info_41_vlWen ),
    .io_diffCommits_info_42_ldest ( io_diffCommits_info_42_ldest ),
    .io_diffCommits_info_42_pdest ( io_diffCommits_info_42_pdest ),
    .io_diffCommits_info_42_rfWen ( io_diffCommits_info_42_rfWen ),
    .io_diffCommits_info_42_fpWen ( io_diffCommits_info_42_fpWen ),
    .io_diffCommits_info_42_vecWen ( io_diffCommits_info_42_vecWen ),
    .io_diffCommits_info_42_v0Wen ( io_diffCommits_info_42_v0Wen ),
    .io_diffCommits_info_42_vlWen ( io_diffCommits_info_42_vlWen ),
    .io_diffCommits_info_43_ldest ( io_diffCommits_info_43_ldest ),
    .io_diffCommits_info_43_pdest ( io_diffCommits_info_43_pdest ),
    .io_diffCommits_info_43_rfWen ( io_diffCommits_info_43_rfWen ),
    .io_diffCommits_info_43_fpWen ( io_diffCommits_info_43_fpWen ),
    .io_diffCommits_info_43_vecWen ( io_diffCommits_info_43_vecWen ),
    .io_diffCommits_info_43_v0Wen ( io_diffCommits_info_43_v0Wen ),
    .io_diffCommits_info_43_vlWen ( io_diffCommits_info_43_vlWen ),
    .io_diffCommits_info_44_ldest ( io_diffCommits_info_44_ldest ),
    .io_diffCommits_info_44_pdest ( io_diffCommits_info_44_pdest ),
    .io_diffCommits_info_44_rfWen ( io_diffCommits_info_44_rfWen ),
    .io_diffCommits_info_44_fpWen ( io_diffCommits_info_44_fpWen ),
    .io_diffCommits_info_44_vecWen ( io_diffCommits_info_44_vecWen ),
    .io_diffCommits_info_44_v0Wen ( io_diffCommits_info_44_v0Wen ),
    .io_diffCommits_info_44_vlWen ( io_diffCommits_info_44_vlWen ),
    .io_diffCommits_info_45_ldest ( io_diffCommits_info_45_ldest ),
    .io_diffCommits_info_45_pdest ( io_diffCommits_info_45_pdest ),
    .io_diffCommits_info_45_rfWen ( io_diffCommits_info_45_rfWen ),
    .io_diffCommits_info_45_fpWen ( io_diffCommits_info_45_fpWen ),
    .io_diffCommits_info_45_vecWen ( io_diffCommits_info_45_vecWen ),
    .io_diffCommits_info_45_v0Wen ( io_diffCommits_info_45_v0Wen ),
    .io_diffCommits_info_45_vlWen ( io_diffCommits_info_45_vlWen ),
    .io_diffCommits_info_46_ldest ( io_diffCommits_info_46_ldest ),
    .io_diffCommits_info_46_pdest ( io_diffCommits_info_46_pdest ),
    .io_diffCommits_info_46_rfWen ( io_diffCommits_info_46_rfWen ),
    .io_diffCommits_info_46_fpWen ( io_diffCommits_info_46_fpWen ),
    .io_diffCommits_info_46_vecWen ( io_diffCommits_info_46_vecWen ),
    .io_diffCommits_info_46_v0Wen ( io_diffCommits_info_46_v0Wen ),
    .io_diffCommits_info_46_vlWen ( io_diffCommits_info_46_vlWen ),
    .io_diffCommits_info_47_ldest ( io_diffCommits_info_47_ldest ),
    .io_diffCommits_info_47_pdest ( io_diffCommits_info_47_pdest ),
    .io_diffCommits_info_47_rfWen ( io_diffCommits_info_47_rfWen ),
    .io_diffCommits_info_47_fpWen ( io_diffCommits_info_47_fpWen ),
    .io_diffCommits_info_47_vecWen ( io_diffCommits_info_47_vecWen ),
    .io_diffCommits_info_47_v0Wen ( io_diffCommits_info_47_v0Wen ),
    .io_diffCommits_info_47_vlWen ( io_diffCommits_info_47_vlWen ),
    .io_diffCommits_info_48_ldest ( io_diffCommits_info_48_ldest ),
    .io_diffCommits_info_48_pdest ( io_diffCommits_info_48_pdest ),
    .io_diffCommits_info_48_rfWen ( io_diffCommits_info_48_rfWen ),
    .io_diffCommits_info_48_fpWen ( io_diffCommits_info_48_fpWen ),
    .io_diffCommits_info_48_vecWen ( io_diffCommits_info_48_vecWen ),
    .io_diffCommits_info_48_v0Wen ( io_diffCommits_info_48_v0Wen ),
    .io_diffCommits_info_48_vlWen ( io_diffCommits_info_48_vlWen ),
    .io_diffCommits_info_49_ldest ( io_diffCommits_info_49_ldest ),
    .io_diffCommits_info_49_pdest ( io_diffCommits_info_49_pdest ),
    .io_diffCommits_info_49_rfWen ( io_diffCommits_info_49_rfWen ),
    .io_diffCommits_info_49_fpWen ( io_diffCommits_info_49_fpWen ),
    .io_diffCommits_info_49_vecWen ( io_diffCommits_info_49_vecWen ),
    .io_diffCommits_info_49_v0Wen ( io_diffCommits_info_49_v0Wen ),
    .io_diffCommits_info_49_vlWen ( io_diffCommits_info_49_vlWen ),
    .io_diffCommits_info_50_ldest ( io_diffCommits_info_50_ldest ),
    .io_diffCommits_info_50_pdest ( io_diffCommits_info_50_pdest ),
    .io_diffCommits_info_50_rfWen ( io_diffCommits_info_50_rfWen ),
    .io_diffCommits_info_50_fpWen ( io_diffCommits_info_50_fpWen ),
    .io_diffCommits_info_50_vecWen ( io_diffCommits_info_50_vecWen ),
    .io_diffCommits_info_50_v0Wen ( io_diffCommits_info_50_v0Wen ),
    .io_diffCommits_info_50_vlWen ( io_diffCommits_info_50_vlWen ),
    .io_diffCommits_info_51_ldest ( io_diffCommits_info_51_ldest ),
    .io_diffCommits_info_51_pdest ( io_diffCommits_info_51_pdest ),
    .io_diffCommits_info_51_rfWen ( io_diffCommits_info_51_rfWen ),
    .io_diffCommits_info_51_fpWen ( io_diffCommits_info_51_fpWen ),
    .io_diffCommits_info_51_vecWen ( io_diffCommits_info_51_vecWen ),
    .io_diffCommits_info_51_v0Wen ( io_diffCommits_info_51_v0Wen ),
    .io_diffCommits_info_51_vlWen ( io_diffCommits_info_51_vlWen ),
    .io_diffCommits_info_52_ldest ( io_diffCommits_info_52_ldest ),
    .io_diffCommits_info_52_pdest ( io_diffCommits_info_52_pdest ),
    .io_diffCommits_info_52_rfWen ( io_diffCommits_info_52_rfWen ),
    .io_diffCommits_info_52_fpWen ( io_diffCommits_info_52_fpWen ),
    .io_diffCommits_info_52_vecWen ( io_diffCommits_info_52_vecWen ),
    .io_diffCommits_info_52_v0Wen ( io_diffCommits_info_52_v0Wen ),
    .io_diffCommits_info_52_vlWen ( io_diffCommits_info_52_vlWen ),
    .io_diffCommits_info_53_ldest ( io_diffCommits_info_53_ldest ),
    .io_diffCommits_info_53_pdest ( io_diffCommits_info_53_pdest ),
    .io_diffCommits_info_53_rfWen ( io_diffCommits_info_53_rfWen ),
    .io_diffCommits_info_53_fpWen ( io_diffCommits_info_53_fpWen ),
    .io_diffCommits_info_53_vecWen ( io_diffCommits_info_53_vecWen ),
    .io_diffCommits_info_53_v0Wen ( io_diffCommits_info_53_v0Wen ),
    .io_diffCommits_info_53_vlWen ( io_diffCommits_info_53_vlWen ),
    .io_diffCommits_info_54_ldest ( io_diffCommits_info_54_ldest ),
    .io_diffCommits_info_54_pdest ( io_diffCommits_info_54_pdest ),
    .io_diffCommits_info_54_rfWen ( io_diffCommits_info_54_rfWen ),
    .io_diffCommits_info_54_fpWen ( io_diffCommits_info_54_fpWen ),
    .io_diffCommits_info_54_vecWen ( io_diffCommits_info_54_vecWen ),
    .io_diffCommits_info_54_v0Wen ( io_diffCommits_info_54_v0Wen ),
    .io_diffCommits_info_54_vlWen ( io_diffCommits_info_54_vlWen ),
    .io_diffCommits_info_55_ldest ( io_diffCommits_info_55_ldest ),
    .io_diffCommits_info_55_pdest ( io_diffCommits_info_55_pdest ),
    .io_diffCommits_info_55_rfWen ( io_diffCommits_info_55_rfWen ),
    .io_diffCommits_info_55_fpWen ( io_diffCommits_info_55_fpWen ),
    .io_diffCommits_info_55_vecWen ( io_diffCommits_info_55_vecWen ),
    .io_diffCommits_info_55_v0Wen ( io_diffCommits_info_55_v0Wen ),
    .io_diffCommits_info_55_vlWen ( io_diffCommits_info_55_vlWen ),
    .io_diffCommits_info_56_ldest ( io_diffCommits_info_56_ldest ),
    .io_diffCommits_info_56_pdest ( io_diffCommits_info_56_pdest ),
    .io_diffCommits_info_56_rfWen ( io_diffCommits_info_56_rfWen ),
    .io_diffCommits_info_56_fpWen ( io_diffCommits_info_56_fpWen ),
    .io_diffCommits_info_56_vecWen ( io_diffCommits_info_56_vecWen ),
    .io_diffCommits_info_56_v0Wen ( io_diffCommits_info_56_v0Wen ),
    .io_diffCommits_info_56_vlWen ( io_diffCommits_info_56_vlWen ),
    .io_diffCommits_info_57_ldest ( io_diffCommits_info_57_ldest ),
    .io_diffCommits_info_57_pdest ( io_diffCommits_info_57_pdest ),
    .io_diffCommits_info_57_rfWen ( io_diffCommits_info_57_rfWen ),
    .io_diffCommits_info_57_fpWen ( io_diffCommits_info_57_fpWen ),
    .io_diffCommits_info_57_vecWen ( io_diffCommits_info_57_vecWen ),
    .io_diffCommits_info_57_v0Wen ( io_diffCommits_info_57_v0Wen ),
    .io_diffCommits_info_57_vlWen ( io_diffCommits_info_57_vlWen ),
    .io_diffCommits_info_58_ldest ( io_diffCommits_info_58_ldest ),
    .io_diffCommits_info_58_pdest ( io_diffCommits_info_58_pdest ),
    .io_diffCommits_info_58_rfWen ( io_diffCommits_info_58_rfWen ),
    .io_diffCommits_info_58_fpWen ( io_diffCommits_info_58_fpWen ),
    .io_diffCommits_info_58_vecWen ( io_diffCommits_info_58_vecWen ),
    .io_diffCommits_info_58_v0Wen ( io_diffCommits_info_58_v0Wen ),
    .io_diffCommits_info_58_vlWen ( io_diffCommits_info_58_vlWen ),
    .io_diffCommits_info_59_ldest ( io_diffCommits_info_59_ldest ),
    .io_diffCommits_info_59_pdest ( io_diffCommits_info_59_pdest ),
    .io_diffCommits_info_59_rfWen ( io_diffCommits_info_59_rfWen ),
    .io_diffCommits_info_59_fpWen ( io_diffCommits_info_59_fpWen ),
    .io_diffCommits_info_59_vecWen ( io_diffCommits_info_59_vecWen ),
    .io_diffCommits_info_59_v0Wen ( io_diffCommits_info_59_v0Wen ),
    .io_diffCommits_info_59_vlWen ( io_diffCommits_info_59_vlWen ),
    .io_diffCommits_info_60_ldest ( io_diffCommits_info_60_ldest ),
    .io_diffCommits_info_60_pdest ( io_diffCommits_info_60_pdest ),
    .io_diffCommits_info_60_rfWen ( io_diffCommits_info_60_rfWen ),
    .io_diffCommits_info_60_fpWen ( io_diffCommits_info_60_fpWen ),
    .io_diffCommits_info_60_vecWen ( io_diffCommits_info_60_vecWen ),
    .io_diffCommits_info_60_v0Wen ( io_diffCommits_info_60_v0Wen ),
    .io_diffCommits_info_60_vlWen ( io_diffCommits_info_60_vlWen ),
    .io_diffCommits_info_61_ldest ( io_diffCommits_info_61_ldest ),
    .io_diffCommits_info_61_pdest ( io_diffCommits_info_61_pdest ),
    .io_diffCommits_info_61_rfWen ( io_diffCommits_info_61_rfWen ),
    .io_diffCommits_info_61_fpWen ( io_diffCommits_info_61_fpWen ),
    .io_diffCommits_info_61_vecWen ( io_diffCommits_info_61_vecWen ),
    .io_diffCommits_info_61_v0Wen ( io_diffCommits_info_61_v0Wen ),
    .io_diffCommits_info_61_vlWen ( io_diffCommits_info_61_vlWen ),
    .io_diffCommits_info_62_ldest ( io_diffCommits_info_62_ldest ),
    .io_diffCommits_info_62_pdest ( io_diffCommits_info_62_pdest ),
    .io_diffCommits_info_62_rfWen ( io_diffCommits_info_62_rfWen ),
    .io_diffCommits_info_62_fpWen ( io_diffCommits_info_62_fpWen ),
    .io_diffCommits_info_62_vecWen ( io_diffCommits_info_62_vecWen ),
    .io_diffCommits_info_62_v0Wen ( io_diffCommits_info_62_v0Wen ),
    .io_diffCommits_info_62_vlWen ( io_diffCommits_info_62_vlWen ),
    .io_diffCommits_info_63_ldest ( io_diffCommits_info_63_ldest ),
    .io_diffCommits_info_63_pdest ( io_diffCommits_info_63_pdest ),
    .io_diffCommits_info_63_rfWen ( io_diffCommits_info_63_rfWen ),
    .io_diffCommits_info_63_fpWen ( io_diffCommits_info_63_fpWen ),
    .io_diffCommits_info_63_vecWen ( io_diffCommits_info_63_vecWen ),
    .io_diffCommits_info_63_v0Wen ( io_diffCommits_info_63_v0Wen ),
    .io_diffCommits_info_63_vlWen ( io_diffCommits_info_63_vlWen ),
    .io_diffCommits_info_64_ldest ( io_diffCommits_info_64_ldest ),
    .io_diffCommits_info_64_pdest ( io_diffCommits_info_64_pdest ),
    .io_diffCommits_info_64_rfWen ( io_diffCommits_info_64_rfWen ),
    .io_diffCommits_info_64_fpWen ( io_diffCommits_info_64_fpWen ),
    .io_diffCommits_info_64_vecWen ( io_diffCommits_info_64_vecWen ),
    .io_diffCommits_info_64_v0Wen ( io_diffCommits_info_64_v0Wen ),
    .io_diffCommits_info_64_vlWen ( io_diffCommits_info_64_vlWen ),
    .io_diffCommits_info_65_ldest ( io_diffCommits_info_65_ldest ),
    .io_diffCommits_info_65_pdest ( io_diffCommits_info_65_pdest ),
    .io_diffCommits_info_65_rfWen ( io_diffCommits_info_65_rfWen ),
    .io_diffCommits_info_65_fpWen ( io_diffCommits_info_65_fpWen ),
    .io_diffCommits_info_65_vecWen ( io_diffCommits_info_65_vecWen ),
    .io_diffCommits_info_65_v0Wen ( io_diffCommits_info_65_v0Wen ),
    .io_diffCommits_info_65_vlWen ( io_diffCommits_info_65_vlWen ),
    .io_diffCommits_info_66_ldest ( io_diffCommits_info_66_ldest ),
    .io_diffCommits_info_66_pdest ( io_diffCommits_info_66_pdest ),
    .io_diffCommits_info_66_rfWen ( io_diffCommits_info_66_rfWen ),
    .io_diffCommits_info_66_fpWen ( io_diffCommits_info_66_fpWen ),
    .io_diffCommits_info_66_vecWen ( io_diffCommits_info_66_vecWen ),
    .io_diffCommits_info_66_v0Wen ( io_diffCommits_info_66_v0Wen ),
    .io_diffCommits_info_66_vlWen ( io_diffCommits_info_66_vlWen ),
    .io_diffCommits_info_67_ldest ( io_diffCommits_info_67_ldest ),
    .io_diffCommits_info_67_pdest ( io_diffCommits_info_67_pdest ),
    .io_diffCommits_info_67_rfWen ( io_diffCommits_info_67_rfWen ),
    .io_diffCommits_info_67_fpWen ( io_diffCommits_info_67_fpWen ),
    .io_diffCommits_info_67_vecWen ( io_diffCommits_info_67_vecWen ),
    .io_diffCommits_info_67_v0Wen ( io_diffCommits_info_67_v0Wen ),
    .io_diffCommits_info_67_vlWen ( io_diffCommits_info_67_vlWen ),
    .io_diffCommits_info_68_ldest ( io_diffCommits_info_68_ldest ),
    .io_diffCommits_info_68_pdest ( io_diffCommits_info_68_pdest ),
    .io_diffCommits_info_68_rfWen ( io_diffCommits_info_68_rfWen ),
    .io_diffCommits_info_68_fpWen ( io_diffCommits_info_68_fpWen ),
    .io_diffCommits_info_68_vecWen ( io_diffCommits_info_68_vecWen ),
    .io_diffCommits_info_68_v0Wen ( io_diffCommits_info_68_v0Wen ),
    .io_diffCommits_info_68_vlWen ( io_diffCommits_info_68_vlWen ),
    .io_diffCommits_info_69_ldest ( io_diffCommits_info_69_ldest ),
    .io_diffCommits_info_69_pdest ( io_diffCommits_info_69_pdest ),
    .io_diffCommits_info_69_rfWen ( io_diffCommits_info_69_rfWen ),
    .io_diffCommits_info_69_fpWen ( io_diffCommits_info_69_fpWen ),
    .io_diffCommits_info_69_vecWen ( io_diffCommits_info_69_vecWen ),
    .io_diffCommits_info_69_v0Wen ( io_diffCommits_info_69_v0Wen ),
    .io_diffCommits_info_69_vlWen ( io_diffCommits_info_69_vlWen ),
    .io_diffCommits_info_70_ldest ( io_diffCommits_info_70_ldest ),
    .io_diffCommits_info_70_pdest ( io_diffCommits_info_70_pdest ),
    .io_diffCommits_info_70_rfWen ( io_diffCommits_info_70_rfWen ),
    .io_diffCommits_info_70_fpWen ( io_diffCommits_info_70_fpWen ),
    .io_diffCommits_info_70_vecWen ( io_diffCommits_info_70_vecWen ),
    .io_diffCommits_info_70_v0Wen ( io_diffCommits_info_70_v0Wen ),
    .io_diffCommits_info_70_vlWen ( io_diffCommits_info_70_vlWen ),
    .io_diffCommits_info_71_ldest ( io_diffCommits_info_71_ldest ),
    .io_diffCommits_info_71_pdest ( io_diffCommits_info_71_pdest ),
    .io_diffCommits_info_71_rfWen ( io_diffCommits_info_71_rfWen ),
    .io_diffCommits_info_71_fpWen ( io_diffCommits_info_71_fpWen ),
    .io_diffCommits_info_71_vecWen ( io_diffCommits_info_71_vecWen ),
    .io_diffCommits_info_71_v0Wen ( io_diffCommits_info_71_v0Wen ),
    .io_diffCommits_info_71_vlWen ( io_diffCommits_info_71_vlWen ),
    .io_diffCommits_info_72_ldest ( io_diffCommits_info_72_ldest ),
    .io_diffCommits_info_72_pdest ( io_diffCommits_info_72_pdest ),
    .io_diffCommits_info_72_rfWen ( io_diffCommits_info_72_rfWen ),
    .io_diffCommits_info_72_fpWen ( io_diffCommits_info_72_fpWen ),
    .io_diffCommits_info_72_vecWen ( io_diffCommits_info_72_vecWen ),
    .io_diffCommits_info_72_v0Wen ( io_diffCommits_info_72_v0Wen ),
    .io_diffCommits_info_72_vlWen ( io_diffCommits_info_72_vlWen ),
    .io_diffCommits_info_73_ldest ( io_diffCommits_info_73_ldest ),
    .io_diffCommits_info_73_pdest ( io_diffCommits_info_73_pdest ),
    .io_diffCommits_info_73_rfWen ( io_diffCommits_info_73_rfWen ),
    .io_diffCommits_info_73_fpWen ( io_diffCommits_info_73_fpWen ),
    .io_diffCommits_info_73_vecWen ( io_diffCommits_info_73_vecWen ),
    .io_diffCommits_info_73_v0Wen ( io_diffCommits_info_73_v0Wen ),
    .io_diffCommits_info_73_vlWen ( io_diffCommits_info_73_vlWen ),
    .io_diffCommits_info_74_ldest ( io_diffCommits_info_74_ldest ),
    .io_diffCommits_info_74_pdest ( io_diffCommits_info_74_pdest ),
    .io_diffCommits_info_74_rfWen ( io_diffCommits_info_74_rfWen ),
    .io_diffCommits_info_74_fpWen ( io_diffCommits_info_74_fpWen ),
    .io_diffCommits_info_74_vecWen ( io_diffCommits_info_74_vecWen ),
    .io_diffCommits_info_74_v0Wen ( io_diffCommits_info_74_v0Wen ),
    .io_diffCommits_info_74_vlWen ( io_diffCommits_info_74_vlWen ),
    .io_diffCommits_info_75_ldest ( io_diffCommits_info_75_ldest ),
    .io_diffCommits_info_75_pdest ( io_diffCommits_info_75_pdest ),
    .io_diffCommits_info_75_rfWen ( io_diffCommits_info_75_rfWen ),
    .io_diffCommits_info_75_fpWen ( io_diffCommits_info_75_fpWen ),
    .io_diffCommits_info_75_vecWen ( io_diffCommits_info_75_vecWen ),
    .io_diffCommits_info_75_v0Wen ( io_diffCommits_info_75_v0Wen ),
    .io_diffCommits_info_75_vlWen ( io_diffCommits_info_75_vlWen ),
    .io_diffCommits_info_76_ldest ( io_diffCommits_info_76_ldest ),
    .io_diffCommits_info_76_pdest ( io_diffCommits_info_76_pdest ),
    .io_diffCommits_info_76_rfWen ( io_diffCommits_info_76_rfWen ),
    .io_diffCommits_info_76_fpWen ( io_diffCommits_info_76_fpWen ),
    .io_diffCommits_info_76_vecWen ( io_diffCommits_info_76_vecWen ),
    .io_diffCommits_info_76_v0Wen ( io_diffCommits_info_76_v0Wen ),
    .io_diffCommits_info_76_vlWen ( io_diffCommits_info_76_vlWen ),
    .io_diffCommits_info_77_ldest ( io_diffCommits_info_77_ldest ),
    .io_diffCommits_info_77_pdest ( io_diffCommits_info_77_pdest ),
    .io_diffCommits_info_77_rfWen ( io_diffCommits_info_77_rfWen ),
    .io_diffCommits_info_77_fpWen ( io_diffCommits_info_77_fpWen ),
    .io_diffCommits_info_77_vecWen ( io_diffCommits_info_77_vecWen ),
    .io_diffCommits_info_77_v0Wen ( io_diffCommits_info_77_v0Wen ),
    .io_diffCommits_info_77_vlWen ( io_diffCommits_info_77_vlWen ),
    .io_diffCommits_info_78_ldest ( io_diffCommits_info_78_ldest ),
    .io_diffCommits_info_78_pdest ( io_diffCommits_info_78_pdest ),
    .io_diffCommits_info_78_rfWen ( io_diffCommits_info_78_rfWen ),
    .io_diffCommits_info_78_fpWen ( io_diffCommits_info_78_fpWen ),
    .io_diffCommits_info_78_vecWen ( io_diffCommits_info_78_vecWen ),
    .io_diffCommits_info_78_v0Wen ( io_diffCommits_info_78_v0Wen ),
    .io_diffCommits_info_78_vlWen ( io_diffCommits_info_78_vlWen ),
    .io_diffCommits_info_79_ldest ( io_diffCommits_info_79_ldest ),
    .io_diffCommits_info_79_pdest ( io_diffCommits_info_79_pdest ),
    .io_diffCommits_info_79_rfWen ( io_diffCommits_info_79_rfWen ),
    .io_diffCommits_info_79_fpWen ( io_diffCommits_info_79_fpWen ),
    .io_diffCommits_info_79_vecWen ( io_diffCommits_info_79_vecWen ),
    .io_diffCommits_info_79_v0Wen ( io_diffCommits_info_79_v0Wen ),
    .io_diffCommits_info_79_vlWen ( io_diffCommits_info_79_vlWen ),
    .io_diffCommits_info_80_ldest ( io_diffCommits_info_80_ldest ),
    .io_diffCommits_info_80_pdest ( io_diffCommits_info_80_pdest ),
    .io_diffCommits_info_80_rfWen ( io_diffCommits_info_80_rfWen ),
    .io_diffCommits_info_80_fpWen ( io_diffCommits_info_80_fpWen ),
    .io_diffCommits_info_80_vecWen ( io_diffCommits_info_80_vecWen ),
    .io_diffCommits_info_80_v0Wen ( io_diffCommits_info_80_v0Wen ),
    .io_diffCommits_info_80_vlWen ( io_diffCommits_info_80_vlWen ),
    .io_diffCommits_info_81_ldest ( io_diffCommits_info_81_ldest ),
    .io_diffCommits_info_81_pdest ( io_diffCommits_info_81_pdest ),
    .io_diffCommits_info_81_rfWen ( io_diffCommits_info_81_rfWen ),
    .io_diffCommits_info_81_fpWen ( io_diffCommits_info_81_fpWen ),
    .io_diffCommits_info_81_vecWen ( io_diffCommits_info_81_vecWen ),
    .io_diffCommits_info_81_v0Wen ( io_diffCommits_info_81_v0Wen ),
    .io_diffCommits_info_81_vlWen ( io_diffCommits_info_81_vlWen ),
    .io_diffCommits_info_82_ldest ( io_diffCommits_info_82_ldest ),
    .io_diffCommits_info_82_pdest ( io_diffCommits_info_82_pdest ),
    .io_diffCommits_info_82_rfWen ( io_diffCommits_info_82_rfWen ),
    .io_diffCommits_info_82_fpWen ( io_diffCommits_info_82_fpWen ),
    .io_diffCommits_info_82_vecWen ( io_diffCommits_info_82_vecWen ),
    .io_diffCommits_info_82_v0Wen ( io_diffCommits_info_82_v0Wen ),
    .io_diffCommits_info_82_vlWen ( io_diffCommits_info_82_vlWen ),
    .io_diffCommits_info_83_ldest ( io_diffCommits_info_83_ldest ),
    .io_diffCommits_info_83_pdest ( io_diffCommits_info_83_pdest ),
    .io_diffCommits_info_83_rfWen ( io_diffCommits_info_83_rfWen ),
    .io_diffCommits_info_83_fpWen ( io_diffCommits_info_83_fpWen ),
    .io_diffCommits_info_83_vecWen ( io_diffCommits_info_83_vecWen ),
    .io_diffCommits_info_83_v0Wen ( io_diffCommits_info_83_v0Wen ),
    .io_diffCommits_info_83_vlWen ( io_diffCommits_info_83_vlWen ),
    .io_diffCommits_info_84_ldest ( io_diffCommits_info_84_ldest ),
    .io_diffCommits_info_84_pdest ( io_diffCommits_info_84_pdest ),
    .io_diffCommits_info_84_rfWen ( io_diffCommits_info_84_rfWen ),
    .io_diffCommits_info_84_fpWen ( io_diffCommits_info_84_fpWen ),
    .io_diffCommits_info_84_vecWen ( io_diffCommits_info_84_vecWen ),
    .io_diffCommits_info_84_v0Wen ( io_diffCommits_info_84_v0Wen ),
    .io_diffCommits_info_84_vlWen ( io_diffCommits_info_84_vlWen ),
    .io_diffCommits_info_85_ldest ( io_diffCommits_info_85_ldest ),
    .io_diffCommits_info_85_pdest ( io_diffCommits_info_85_pdest ),
    .io_diffCommits_info_85_rfWen ( io_diffCommits_info_85_rfWen ),
    .io_diffCommits_info_85_fpWen ( io_diffCommits_info_85_fpWen ),
    .io_diffCommits_info_85_vecWen ( io_diffCommits_info_85_vecWen ),
    .io_diffCommits_info_85_v0Wen ( io_diffCommits_info_85_v0Wen ),
    .io_diffCommits_info_85_vlWen ( io_diffCommits_info_85_vlWen ),
    .io_diffCommits_info_86_ldest ( io_diffCommits_info_86_ldest ),
    .io_diffCommits_info_86_pdest ( io_diffCommits_info_86_pdest ),
    .io_diffCommits_info_86_rfWen ( io_diffCommits_info_86_rfWen ),
    .io_diffCommits_info_86_fpWen ( io_diffCommits_info_86_fpWen ),
    .io_diffCommits_info_86_vecWen ( io_diffCommits_info_86_vecWen ),
    .io_diffCommits_info_86_v0Wen ( io_diffCommits_info_86_v0Wen ),
    .io_diffCommits_info_86_vlWen ( io_diffCommits_info_86_vlWen ),
    .io_diffCommits_info_87_ldest ( io_diffCommits_info_87_ldest ),
    .io_diffCommits_info_87_pdest ( io_diffCommits_info_87_pdest ),
    .io_diffCommits_info_87_rfWen ( io_diffCommits_info_87_rfWen ),
    .io_diffCommits_info_87_fpWen ( io_diffCommits_info_87_fpWen ),
    .io_diffCommits_info_87_vecWen ( io_diffCommits_info_87_vecWen ),
    .io_diffCommits_info_87_v0Wen ( io_diffCommits_info_87_v0Wen ),
    .io_diffCommits_info_87_vlWen ( io_diffCommits_info_87_vlWen ),
    .io_diffCommits_info_88_ldest ( io_diffCommits_info_88_ldest ),
    .io_diffCommits_info_88_pdest ( io_diffCommits_info_88_pdest ),
    .io_diffCommits_info_88_rfWen ( io_diffCommits_info_88_rfWen ),
    .io_diffCommits_info_88_fpWen ( io_diffCommits_info_88_fpWen ),
    .io_diffCommits_info_88_vecWen ( io_diffCommits_info_88_vecWen ),
    .io_diffCommits_info_88_v0Wen ( io_diffCommits_info_88_v0Wen ),
    .io_diffCommits_info_88_vlWen ( io_diffCommits_info_88_vlWen ),
    .io_diffCommits_info_89_ldest ( io_diffCommits_info_89_ldest ),
    .io_diffCommits_info_89_pdest ( io_diffCommits_info_89_pdest ),
    .io_diffCommits_info_89_rfWen ( io_diffCommits_info_89_rfWen ),
    .io_diffCommits_info_89_fpWen ( io_diffCommits_info_89_fpWen ),
    .io_diffCommits_info_89_vecWen ( io_diffCommits_info_89_vecWen ),
    .io_diffCommits_info_89_v0Wen ( io_diffCommits_info_89_v0Wen ),
    .io_diffCommits_info_89_vlWen ( io_diffCommits_info_89_vlWen ),
    .io_diffCommits_info_90_ldest ( io_diffCommits_info_90_ldest ),
    .io_diffCommits_info_90_pdest ( io_diffCommits_info_90_pdest ),
    .io_diffCommits_info_90_rfWen ( io_diffCommits_info_90_rfWen ),
    .io_diffCommits_info_90_fpWen ( io_diffCommits_info_90_fpWen ),
    .io_diffCommits_info_90_vecWen ( io_diffCommits_info_90_vecWen ),
    .io_diffCommits_info_90_v0Wen ( io_diffCommits_info_90_v0Wen ),
    .io_diffCommits_info_90_vlWen ( io_diffCommits_info_90_vlWen ),
    .io_diffCommits_info_91_ldest ( io_diffCommits_info_91_ldest ),
    .io_diffCommits_info_91_pdest ( io_diffCommits_info_91_pdest ),
    .io_diffCommits_info_91_rfWen ( io_diffCommits_info_91_rfWen ),
    .io_diffCommits_info_91_fpWen ( io_diffCommits_info_91_fpWen ),
    .io_diffCommits_info_91_vecWen ( io_diffCommits_info_91_vecWen ),
    .io_diffCommits_info_91_v0Wen ( io_diffCommits_info_91_v0Wen ),
    .io_diffCommits_info_91_vlWen ( io_diffCommits_info_91_vlWen ),
    .io_diffCommits_info_92_ldest ( io_diffCommits_info_92_ldest ),
    .io_diffCommits_info_92_pdest ( io_diffCommits_info_92_pdest ),
    .io_diffCommits_info_92_rfWen ( io_diffCommits_info_92_rfWen ),
    .io_diffCommits_info_92_fpWen ( io_diffCommits_info_92_fpWen ),
    .io_diffCommits_info_92_vecWen ( io_diffCommits_info_92_vecWen ),
    .io_diffCommits_info_92_v0Wen ( io_diffCommits_info_92_v0Wen ),
    .io_diffCommits_info_92_vlWen ( io_diffCommits_info_92_vlWen ),
    .io_diffCommits_info_93_ldest ( io_diffCommits_info_93_ldest ),
    .io_diffCommits_info_93_pdest ( io_diffCommits_info_93_pdest ),
    .io_diffCommits_info_93_rfWen ( io_diffCommits_info_93_rfWen ),
    .io_diffCommits_info_93_fpWen ( io_diffCommits_info_93_fpWen ),
    .io_diffCommits_info_93_vecWen ( io_diffCommits_info_93_vecWen ),
    .io_diffCommits_info_93_v0Wen ( io_diffCommits_info_93_v0Wen ),
    .io_diffCommits_info_93_vlWen ( io_diffCommits_info_93_vlWen ),
    .io_diffCommits_info_94_ldest ( io_diffCommits_info_94_ldest ),
    .io_diffCommits_info_94_pdest ( io_diffCommits_info_94_pdest ),
    .io_diffCommits_info_94_rfWen ( io_diffCommits_info_94_rfWen ),
    .io_diffCommits_info_94_fpWen ( io_diffCommits_info_94_fpWen ),
    .io_diffCommits_info_94_vecWen ( io_diffCommits_info_94_vecWen ),
    .io_diffCommits_info_94_v0Wen ( io_diffCommits_info_94_v0Wen ),
    .io_diffCommits_info_94_vlWen ( io_diffCommits_info_94_vlWen ),
    .io_diffCommits_info_95_ldest ( io_diffCommits_info_95_ldest ),
    .io_diffCommits_info_95_pdest ( io_diffCommits_info_95_pdest ),
    .io_diffCommits_info_95_rfWen ( io_diffCommits_info_95_rfWen ),
    .io_diffCommits_info_95_fpWen ( io_diffCommits_info_95_fpWen ),
    .io_diffCommits_info_95_vecWen ( io_diffCommits_info_95_vecWen ),
    .io_diffCommits_info_95_v0Wen ( io_diffCommits_info_95_v0Wen ),
    .io_diffCommits_info_95_vlWen ( io_diffCommits_info_95_vlWen ),
    .io_diffCommits_info_96_ldest ( io_diffCommits_info_96_ldest ),
    .io_diffCommits_info_96_pdest ( io_diffCommits_info_96_pdest ),
    .io_diffCommits_info_96_rfWen ( io_diffCommits_info_96_rfWen ),
    .io_diffCommits_info_96_fpWen ( io_diffCommits_info_96_fpWen ),
    .io_diffCommits_info_96_vecWen ( io_diffCommits_info_96_vecWen ),
    .io_diffCommits_info_96_v0Wen ( io_diffCommits_info_96_v0Wen ),
    .io_diffCommits_info_96_vlWen ( io_diffCommits_info_96_vlWen ),
    .io_diffCommits_info_97_ldest ( io_diffCommits_info_97_ldest ),
    .io_diffCommits_info_97_pdest ( io_diffCommits_info_97_pdest ),
    .io_diffCommits_info_97_rfWen ( io_diffCommits_info_97_rfWen ),
    .io_diffCommits_info_97_fpWen ( io_diffCommits_info_97_fpWen ),
    .io_diffCommits_info_97_vecWen ( io_diffCommits_info_97_vecWen ),
    .io_diffCommits_info_97_v0Wen ( io_diffCommits_info_97_v0Wen ),
    .io_diffCommits_info_97_vlWen ( io_diffCommits_info_97_vlWen ),
    .io_diffCommits_info_98_ldest ( io_diffCommits_info_98_ldest ),
    .io_diffCommits_info_98_pdest ( io_diffCommits_info_98_pdest ),
    .io_diffCommits_info_98_rfWen ( io_diffCommits_info_98_rfWen ),
    .io_diffCommits_info_98_fpWen ( io_diffCommits_info_98_fpWen ),
    .io_diffCommits_info_98_vecWen ( io_diffCommits_info_98_vecWen ),
    .io_diffCommits_info_98_v0Wen ( io_diffCommits_info_98_v0Wen ),
    .io_diffCommits_info_98_vlWen ( io_diffCommits_info_98_vlWen ),
    .io_diffCommits_info_99_ldest ( io_diffCommits_info_99_ldest ),
    .io_diffCommits_info_99_pdest ( io_diffCommits_info_99_pdest ),
    .io_diffCommits_info_99_rfWen ( io_diffCommits_info_99_rfWen ),
    .io_diffCommits_info_99_fpWen ( io_diffCommits_info_99_fpWen ),
    .io_diffCommits_info_99_vecWen ( io_diffCommits_info_99_vecWen ),
    .io_diffCommits_info_99_v0Wen ( io_diffCommits_info_99_v0Wen ),
    .io_diffCommits_info_99_vlWen ( io_diffCommits_info_99_vlWen ),
    .io_diffCommits_info_100_ldest ( io_diffCommits_info_100_ldest ),
    .io_diffCommits_info_100_pdest ( io_diffCommits_info_100_pdest ),
    .io_diffCommits_info_100_rfWen ( io_diffCommits_info_100_rfWen ),
    .io_diffCommits_info_100_fpWen ( io_diffCommits_info_100_fpWen ),
    .io_diffCommits_info_100_vecWen ( io_diffCommits_info_100_vecWen ),
    .io_diffCommits_info_100_v0Wen ( io_diffCommits_info_100_v0Wen ),
    .io_diffCommits_info_100_vlWen ( io_diffCommits_info_100_vlWen ),
    .io_diffCommits_info_101_ldest ( io_diffCommits_info_101_ldest ),
    .io_diffCommits_info_101_pdest ( io_diffCommits_info_101_pdest ),
    .io_diffCommits_info_101_rfWen ( io_diffCommits_info_101_rfWen ),
    .io_diffCommits_info_101_fpWen ( io_diffCommits_info_101_fpWen ),
    .io_diffCommits_info_101_vecWen ( io_diffCommits_info_101_vecWen ),
    .io_diffCommits_info_101_v0Wen ( io_diffCommits_info_101_v0Wen ),
    .io_diffCommits_info_101_vlWen ( io_diffCommits_info_101_vlWen ),
    .io_diffCommits_info_102_ldest ( io_diffCommits_info_102_ldest ),
    .io_diffCommits_info_102_pdest ( io_diffCommits_info_102_pdest ),
    .io_diffCommits_info_102_rfWen ( io_diffCommits_info_102_rfWen ),
    .io_diffCommits_info_102_fpWen ( io_diffCommits_info_102_fpWen ),
    .io_diffCommits_info_102_vecWen ( io_diffCommits_info_102_vecWen ),
    .io_diffCommits_info_102_v0Wen ( io_diffCommits_info_102_v0Wen ),
    .io_diffCommits_info_102_vlWen ( io_diffCommits_info_102_vlWen ),
    .io_diffCommits_info_103_ldest ( io_diffCommits_info_103_ldest ),
    .io_diffCommits_info_103_pdest ( io_diffCommits_info_103_pdest ),
    .io_diffCommits_info_103_rfWen ( io_diffCommits_info_103_rfWen ),
    .io_diffCommits_info_103_fpWen ( io_diffCommits_info_103_fpWen ),
    .io_diffCommits_info_103_vecWen ( io_diffCommits_info_103_vecWen ),
    .io_diffCommits_info_103_v0Wen ( io_diffCommits_info_103_v0Wen ),
    .io_diffCommits_info_103_vlWen ( io_diffCommits_info_103_vlWen ),
    .io_diffCommits_info_104_ldest ( io_diffCommits_info_104_ldest ),
    .io_diffCommits_info_104_pdest ( io_diffCommits_info_104_pdest ),
    .io_diffCommits_info_104_rfWen ( io_diffCommits_info_104_rfWen ),
    .io_diffCommits_info_104_fpWen ( io_diffCommits_info_104_fpWen ),
    .io_diffCommits_info_104_vecWen ( io_diffCommits_info_104_vecWen ),
    .io_diffCommits_info_104_v0Wen ( io_diffCommits_info_104_v0Wen ),
    .io_diffCommits_info_104_vlWen ( io_diffCommits_info_104_vlWen ),
    .io_diffCommits_info_105_ldest ( io_diffCommits_info_105_ldest ),
    .io_diffCommits_info_105_pdest ( io_diffCommits_info_105_pdest ),
    .io_diffCommits_info_105_rfWen ( io_diffCommits_info_105_rfWen ),
    .io_diffCommits_info_105_fpWen ( io_diffCommits_info_105_fpWen ),
    .io_diffCommits_info_105_vecWen ( io_diffCommits_info_105_vecWen ),
    .io_diffCommits_info_105_v0Wen ( io_diffCommits_info_105_v0Wen ),
    .io_diffCommits_info_105_vlWen ( io_diffCommits_info_105_vlWen ),
    .io_diffCommits_info_106_ldest ( io_diffCommits_info_106_ldest ),
    .io_diffCommits_info_106_pdest ( io_diffCommits_info_106_pdest ),
    .io_diffCommits_info_106_rfWen ( io_diffCommits_info_106_rfWen ),
    .io_diffCommits_info_106_fpWen ( io_diffCommits_info_106_fpWen ),
    .io_diffCommits_info_106_vecWen ( io_diffCommits_info_106_vecWen ),
    .io_diffCommits_info_106_v0Wen ( io_diffCommits_info_106_v0Wen ),
    .io_diffCommits_info_106_vlWen ( io_diffCommits_info_106_vlWen ),
    .io_diffCommits_info_107_ldest ( io_diffCommits_info_107_ldest ),
    .io_diffCommits_info_107_pdest ( io_diffCommits_info_107_pdest ),
    .io_diffCommits_info_107_rfWen ( io_diffCommits_info_107_rfWen ),
    .io_diffCommits_info_107_fpWen ( io_diffCommits_info_107_fpWen ),
    .io_diffCommits_info_107_vecWen ( io_diffCommits_info_107_vecWen ),
    .io_diffCommits_info_107_v0Wen ( io_diffCommits_info_107_v0Wen ),
    .io_diffCommits_info_107_vlWen ( io_diffCommits_info_107_vlWen ),
    .io_diffCommits_info_108_ldest ( io_diffCommits_info_108_ldest ),
    .io_diffCommits_info_108_pdest ( io_diffCommits_info_108_pdest ),
    .io_diffCommits_info_108_rfWen ( io_diffCommits_info_108_rfWen ),
    .io_diffCommits_info_108_fpWen ( io_diffCommits_info_108_fpWen ),
    .io_diffCommits_info_108_vecWen ( io_diffCommits_info_108_vecWen ),
    .io_diffCommits_info_108_v0Wen ( io_diffCommits_info_108_v0Wen ),
    .io_diffCommits_info_108_vlWen ( io_diffCommits_info_108_vlWen ),
    .io_diffCommits_info_109_ldest ( io_diffCommits_info_109_ldest ),
    .io_diffCommits_info_109_pdest ( io_diffCommits_info_109_pdest ),
    .io_diffCommits_info_109_rfWen ( io_diffCommits_info_109_rfWen ),
    .io_diffCommits_info_109_fpWen ( io_diffCommits_info_109_fpWen ),
    .io_diffCommits_info_109_vecWen ( io_diffCommits_info_109_vecWen ),
    .io_diffCommits_info_109_v0Wen ( io_diffCommits_info_109_v0Wen ),
    .io_diffCommits_info_109_vlWen ( io_diffCommits_info_109_vlWen ),
    .io_diffCommits_info_110_ldest ( io_diffCommits_info_110_ldest ),
    .io_diffCommits_info_110_pdest ( io_diffCommits_info_110_pdest ),
    .io_diffCommits_info_110_rfWen ( io_diffCommits_info_110_rfWen ),
    .io_diffCommits_info_110_fpWen ( io_diffCommits_info_110_fpWen ),
    .io_diffCommits_info_110_vecWen ( io_diffCommits_info_110_vecWen ),
    .io_diffCommits_info_110_v0Wen ( io_diffCommits_info_110_v0Wen ),
    .io_diffCommits_info_110_vlWen ( io_diffCommits_info_110_vlWen ),
    .io_diffCommits_info_111_ldest ( io_diffCommits_info_111_ldest ),
    .io_diffCommits_info_111_pdest ( io_diffCommits_info_111_pdest ),
    .io_diffCommits_info_111_rfWen ( io_diffCommits_info_111_rfWen ),
    .io_diffCommits_info_111_fpWen ( io_diffCommits_info_111_fpWen ),
    .io_diffCommits_info_111_vecWen ( io_diffCommits_info_111_vecWen ),
    .io_diffCommits_info_111_v0Wen ( io_diffCommits_info_111_v0Wen ),
    .io_diffCommits_info_111_vlWen ( io_diffCommits_info_111_vlWen ),
    .io_diffCommits_info_112_ldest ( io_diffCommits_info_112_ldest ),
    .io_diffCommits_info_112_pdest ( io_diffCommits_info_112_pdest ),
    .io_diffCommits_info_112_rfWen ( io_diffCommits_info_112_rfWen ),
    .io_diffCommits_info_112_fpWen ( io_diffCommits_info_112_fpWen ),
    .io_diffCommits_info_112_vecWen ( io_diffCommits_info_112_vecWen ),
    .io_diffCommits_info_112_v0Wen ( io_diffCommits_info_112_v0Wen ),
    .io_diffCommits_info_112_vlWen ( io_diffCommits_info_112_vlWen ),
    .io_diffCommits_info_113_ldest ( io_diffCommits_info_113_ldest ),
    .io_diffCommits_info_113_pdest ( io_diffCommits_info_113_pdest ),
    .io_diffCommits_info_113_rfWen ( io_diffCommits_info_113_rfWen ),
    .io_diffCommits_info_113_fpWen ( io_diffCommits_info_113_fpWen ),
    .io_diffCommits_info_113_vecWen ( io_diffCommits_info_113_vecWen ),
    .io_diffCommits_info_113_v0Wen ( io_diffCommits_info_113_v0Wen ),
    .io_diffCommits_info_113_vlWen ( io_diffCommits_info_113_vlWen ),
    .io_diffCommits_info_114_ldest ( io_diffCommits_info_114_ldest ),
    .io_diffCommits_info_114_pdest ( io_diffCommits_info_114_pdest ),
    .io_diffCommits_info_114_rfWen ( io_diffCommits_info_114_rfWen ),
    .io_diffCommits_info_114_fpWen ( io_diffCommits_info_114_fpWen ),
    .io_diffCommits_info_114_vecWen ( io_diffCommits_info_114_vecWen ),
    .io_diffCommits_info_114_v0Wen ( io_diffCommits_info_114_v0Wen ),
    .io_diffCommits_info_114_vlWen ( io_diffCommits_info_114_vlWen ),
    .io_diffCommits_info_115_ldest ( io_diffCommits_info_115_ldest ),
    .io_diffCommits_info_115_pdest ( io_diffCommits_info_115_pdest ),
    .io_diffCommits_info_115_rfWen ( io_diffCommits_info_115_rfWen ),
    .io_diffCommits_info_115_fpWen ( io_diffCommits_info_115_fpWen ),
    .io_diffCommits_info_115_vecWen ( io_diffCommits_info_115_vecWen ),
    .io_diffCommits_info_115_v0Wen ( io_diffCommits_info_115_v0Wen ),
    .io_diffCommits_info_115_vlWen ( io_diffCommits_info_115_vlWen ),
    .io_diffCommits_info_116_ldest ( io_diffCommits_info_116_ldest ),
    .io_diffCommits_info_116_pdest ( io_diffCommits_info_116_pdest ),
    .io_diffCommits_info_116_rfWen ( io_diffCommits_info_116_rfWen ),
    .io_diffCommits_info_116_fpWen ( io_diffCommits_info_116_fpWen ),
    .io_diffCommits_info_116_vecWen ( io_diffCommits_info_116_vecWen ),
    .io_diffCommits_info_116_v0Wen ( io_diffCommits_info_116_v0Wen ),
    .io_diffCommits_info_116_vlWen ( io_diffCommits_info_116_vlWen ),
    .io_diffCommits_info_117_ldest ( io_diffCommits_info_117_ldest ),
    .io_diffCommits_info_117_pdest ( io_diffCommits_info_117_pdest ),
    .io_diffCommits_info_117_rfWen ( io_diffCommits_info_117_rfWen ),
    .io_diffCommits_info_117_fpWen ( io_diffCommits_info_117_fpWen ),
    .io_diffCommits_info_117_vecWen ( io_diffCommits_info_117_vecWen ),
    .io_diffCommits_info_117_v0Wen ( io_diffCommits_info_117_v0Wen ),
    .io_diffCommits_info_117_vlWen ( io_diffCommits_info_117_vlWen ),
    .io_diffCommits_info_118_ldest ( io_diffCommits_info_118_ldest ),
    .io_diffCommits_info_118_pdest ( io_diffCommits_info_118_pdest ),
    .io_diffCommits_info_118_rfWen ( io_diffCommits_info_118_rfWen ),
    .io_diffCommits_info_118_fpWen ( io_diffCommits_info_118_fpWen ),
    .io_diffCommits_info_118_vecWen ( io_diffCommits_info_118_vecWen ),
    .io_diffCommits_info_118_v0Wen ( io_diffCommits_info_118_v0Wen ),
    .io_diffCommits_info_118_vlWen ( io_diffCommits_info_118_vlWen ),
    .io_diffCommits_info_119_ldest ( io_diffCommits_info_119_ldest ),
    .io_diffCommits_info_119_pdest ( io_diffCommits_info_119_pdest ),
    .io_diffCommits_info_119_rfWen ( io_diffCommits_info_119_rfWen ),
    .io_diffCommits_info_119_fpWen ( io_diffCommits_info_119_fpWen ),
    .io_diffCommits_info_119_vecWen ( io_diffCommits_info_119_vecWen ),
    .io_diffCommits_info_119_v0Wen ( io_diffCommits_info_119_v0Wen ),
    .io_diffCommits_info_119_vlWen ( io_diffCommits_info_119_vlWen ),
    .io_diffCommits_info_120_ldest ( io_diffCommits_info_120_ldest ),
    .io_diffCommits_info_120_pdest ( io_diffCommits_info_120_pdest ),
    .io_diffCommits_info_120_rfWen ( io_diffCommits_info_120_rfWen ),
    .io_diffCommits_info_120_fpWen ( io_diffCommits_info_120_fpWen ),
    .io_diffCommits_info_120_vecWen ( io_diffCommits_info_120_vecWen ),
    .io_diffCommits_info_120_v0Wen ( io_diffCommits_info_120_v0Wen ),
    .io_diffCommits_info_120_vlWen ( io_diffCommits_info_120_vlWen ),
    .io_diffCommits_info_121_ldest ( io_diffCommits_info_121_ldest ),
    .io_diffCommits_info_121_pdest ( io_diffCommits_info_121_pdest ),
    .io_diffCommits_info_121_rfWen ( io_diffCommits_info_121_rfWen ),
    .io_diffCommits_info_121_fpWen ( io_diffCommits_info_121_fpWen ),
    .io_diffCommits_info_121_vecWen ( io_diffCommits_info_121_vecWen ),
    .io_diffCommits_info_121_v0Wen ( io_diffCommits_info_121_v0Wen ),
    .io_diffCommits_info_121_vlWen ( io_diffCommits_info_121_vlWen ),
    .io_diffCommits_info_122_ldest ( io_diffCommits_info_122_ldest ),
    .io_diffCommits_info_122_pdest ( io_diffCommits_info_122_pdest ),
    .io_diffCommits_info_122_rfWen ( io_diffCommits_info_122_rfWen ),
    .io_diffCommits_info_122_fpWen ( io_diffCommits_info_122_fpWen ),
    .io_diffCommits_info_122_vecWen ( io_diffCommits_info_122_vecWen ),
    .io_diffCommits_info_122_v0Wen ( io_diffCommits_info_122_v0Wen ),
    .io_diffCommits_info_122_vlWen ( io_diffCommits_info_122_vlWen ),
    .io_diffCommits_info_123_ldest ( io_diffCommits_info_123_ldest ),
    .io_diffCommits_info_123_pdest ( io_diffCommits_info_123_pdest ),
    .io_diffCommits_info_123_rfWen ( io_diffCommits_info_123_rfWen ),
    .io_diffCommits_info_123_fpWen ( io_diffCommits_info_123_fpWen ),
    .io_diffCommits_info_123_vecWen ( io_diffCommits_info_123_vecWen ),
    .io_diffCommits_info_123_v0Wen ( io_diffCommits_info_123_v0Wen ),
    .io_diffCommits_info_123_vlWen ( io_diffCommits_info_123_vlWen ),
    .io_diffCommits_info_124_ldest ( io_diffCommits_info_124_ldest ),
    .io_diffCommits_info_124_pdest ( io_diffCommits_info_124_pdest ),
    .io_diffCommits_info_124_rfWen ( io_diffCommits_info_124_rfWen ),
    .io_diffCommits_info_124_fpWen ( io_diffCommits_info_124_fpWen ),
    .io_diffCommits_info_124_vecWen ( io_diffCommits_info_124_vecWen ),
    .io_diffCommits_info_124_v0Wen ( io_diffCommits_info_124_v0Wen ),
    .io_diffCommits_info_124_vlWen ( io_diffCommits_info_124_vlWen ),
    .io_diffCommits_info_125_ldest ( io_diffCommits_info_125_ldest ),
    .io_diffCommits_info_125_pdest ( io_diffCommits_info_125_pdest ),
    .io_diffCommits_info_125_rfWen ( io_diffCommits_info_125_rfWen ),
    .io_diffCommits_info_125_fpWen ( io_diffCommits_info_125_fpWen ),
    .io_diffCommits_info_125_vecWen ( io_diffCommits_info_125_vecWen ),
    .io_diffCommits_info_125_v0Wen ( io_diffCommits_info_125_v0Wen ),
    .io_diffCommits_info_125_vlWen ( io_diffCommits_info_125_vlWen ),
    .io_diffCommits_info_126_ldest ( io_diffCommits_info_126_ldest ),
    .io_diffCommits_info_126_pdest ( io_diffCommits_info_126_pdest ),
    .io_diffCommits_info_126_rfWen ( io_diffCommits_info_126_rfWen ),
    .io_diffCommits_info_126_fpWen ( io_diffCommits_info_126_fpWen ),
    .io_diffCommits_info_126_vecWen ( io_diffCommits_info_126_vecWen ),
    .io_diffCommits_info_126_v0Wen ( io_diffCommits_info_126_v0Wen ),
    .io_diffCommits_info_126_vlWen ( io_diffCommits_info_126_vlWen ),
    .io_diffCommits_info_127_ldest ( io_diffCommits_info_127_ldest ),
    .io_diffCommits_info_127_pdest ( io_diffCommits_info_127_pdest ),
    .io_diffCommits_info_127_rfWen ( io_diffCommits_info_127_rfWen ),
    .io_diffCommits_info_127_fpWen ( io_diffCommits_info_127_fpWen ),
    .io_diffCommits_info_127_vecWen ( io_diffCommits_info_127_vecWen ),
    .io_diffCommits_info_127_v0Wen ( io_diffCommits_info_127_v0Wen ),
    .io_diffCommits_info_127_vlWen ( io_diffCommits_info_127_vlWen ),
    .io_diffCommits_info_128_ldest ( io_diffCommits_info_128_ldest ),
    .io_diffCommits_info_128_pdest ( io_diffCommits_info_128_pdest ),
    .io_diffCommits_info_128_rfWen ( io_diffCommits_info_128_rfWen ),
    .io_diffCommits_info_128_fpWen ( io_diffCommits_info_128_fpWen ),
    .io_diffCommits_info_128_vecWen ( io_diffCommits_info_128_vecWen ),
    .io_diffCommits_info_128_v0Wen ( io_diffCommits_info_128_v0Wen ),
    .io_diffCommits_info_128_vlWen ( io_diffCommits_info_128_vlWen ),
    .io_diffCommits_info_129_ldest ( io_diffCommits_info_129_ldest ),
    .io_diffCommits_info_129_pdest ( io_diffCommits_info_129_pdest ),
    .io_diffCommits_info_129_rfWen ( io_diffCommits_info_129_rfWen ),
    .io_diffCommits_info_129_fpWen ( io_diffCommits_info_129_fpWen ),
    .io_diffCommits_info_129_vecWen ( io_diffCommits_info_129_vecWen ),
    .io_diffCommits_info_129_v0Wen ( io_diffCommits_info_129_v0Wen ),
    .io_diffCommits_info_129_vlWen ( io_diffCommits_info_129_vlWen ),
    .io_diffCommits_info_130_ldest ( io_diffCommits_info_130_ldest ),
    .io_diffCommits_info_130_pdest ( io_diffCommits_info_130_pdest ),
    .io_diffCommits_info_130_rfWen ( io_diffCommits_info_130_rfWen ),
    .io_diffCommits_info_130_fpWen ( io_diffCommits_info_130_fpWen ),
    .io_diffCommits_info_130_vecWen ( io_diffCommits_info_130_vecWen ),
    .io_diffCommits_info_130_v0Wen ( io_diffCommits_info_130_v0Wen ),
    .io_diffCommits_info_130_vlWen ( io_diffCommits_info_130_vlWen ),
    .io_diffCommits_info_131_ldest ( io_diffCommits_info_131_ldest ),
    .io_diffCommits_info_131_pdest ( io_diffCommits_info_131_pdest ),
    .io_diffCommits_info_131_rfWen ( io_diffCommits_info_131_rfWen ),
    .io_diffCommits_info_131_fpWen ( io_diffCommits_info_131_fpWen ),
    .io_diffCommits_info_131_vecWen ( io_diffCommits_info_131_vecWen ),
    .io_diffCommits_info_131_v0Wen ( io_diffCommits_info_131_v0Wen ),
    .io_diffCommits_info_131_vlWen ( io_diffCommits_info_131_vlWen ),
    .io_diffCommits_info_132_ldest ( io_diffCommits_info_132_ldest ),
    .io_diffCommits_info_132_pdest ( io_diffCommits_info_132_pdest ),
    .io_diffCommits_info_132_rfWen ( io_diffCommits_info_132_rfWen ),
    .io_diffCommits_info_132_fpWen ( io_diffCommits_info_132_fpWen ),
    .io_diffCommits_info_132_vecWen ( io_diffCommits_info_132_vecWen ),
    .io_diffCommits_info_132_v0Wen ( io_diffCommits_info_132_v0Wen ),
    .io_diffCommits_info_132_vlWen ( io_diffCommits_info_132_vlWen ),
    .io_diffCommits_info_133_ldest ( io_diffCommits_info_133_ldest ),
    .io_diffCommits_info_133_pdest ( io_diffCommits_info_133_pdest ),
    .io_diffCommits_info_133_rfWen ( io_diffCommits_info_133_rfWen ),
    .io_diffCommits_info_133_fpWen ( io_diffCommits_info_133_fpWen ),
    .io_diffCommits_info_133_vecWen ( io_diffCommits_info_133_vecWen ),
    .io_diffCommits_info_133_v0Wen ( io_diffCommits_info_133_v0Wen ),
    .io_diffCommits_info_133_vlWen ( io_diffCommits_info_133_vlWen ),
    .io_diffCommits_info_134_ldest ( io_diffCommits_info_134_ldest ),
    .io_diffCommits_info_134_pdest ( io_diffCommits_info_134_pdest ),
    .io_diffCommits_info_134_rfWen ( io_diffCommits_info_134_rfWen ),
    .io_diffCommits_info_134_fpWen ( io_diffCommits_info_134_fpWen ),
    .io_diffCommits_info_134_vecWen ( io_diffCommits_info_134_vecWen ),
    .io_diffCommits_info_134_v0Wen ( io_diffCommits_info_134_v0Wen ),
    .io_diffCommits_info_134_vlWen ( io_diffCommits_info_134_vlWen ),
    .io_diffCommits_info_135_ldest ( io_diffCommits_info_135_ldest ),
    .io_diffCommits_info_135_pdest ( io_diffCommits_info_135_pdest ),
    .io_diffCommits_info_135_rfWen ( io_diffCommits_info_135_rfWen ),
    .io_diffCommits_info_135_fpWen ( io_diffCommits_info_135_fpWen ),
    .io_diffCommits_info_135_vecWen ( io_diffCommits_info_135_vecWen ),
    .io_diffCommits_info_135_v0Wen ( io_diffCommits_info_135_v0Wen ),
    .io_diffCommits_info_135_vlWen ( io_diffCommits_info_135_vlWen ),
    .io_diffCommits_info_136_ldest ( io_diffCommits_info_136_ldest ),
    .io_diffCommits_info_136_pdest ( io_diffCommits_info_136_pdest ),
    .io_diffCommits_info_136_rfWen ( io_diffCommits_info_136_rfWen ),
    .io_diffCommits_info_136_fpWen ( io_diffCommits_info_136_fpWen ),
    .io_diffCommits_info_136_vecWen ( io_diffCommits_info_136_vecWen ),
    .io_diffCommits_info_136_v0Wen ( io_diffCommits_info_136_v0Wen ),
    .io_diffCommits_info_136_vlWen ( io_diffCommits_info_136_vlWen ),
    .io_diffCommits_info_137_ldest ( io_diffCommits_info_137_ldest ),
    .io_diffCommits_info_137_pdest ( io_diffCommits_info_137_pdest ),
    .io_diffCommits_info_137_rfWen ( io_diffCommits_info_137_rfWen ),
    .io_diffCommits_info_137_fpWen ( io_diffCommits_info_137_fpWen ),
    .io_diffCommits_info_137_vecWen ( io_diffCommits_info_137_vecWen ),
    .io_diffCommits_info_137_v0Wen ( io_diffCommits_info_137_v0Wen ),
    .io_diffCommits_info_137_vlWen ( io_diffCommits_info_137_vlWen ),
    .io_diffCommits_info_138_ldest ( io_diffCommits_info_138_ldest ),
    .io_diffCommits_info_138_pdest ( io_diffCommits_info_138_pdest ),
    .io_diffCommits_info_138_rfWen ( io_diffCommits_info_138_rfWen ),
    .io_diffCommits_info_138_fpWen ( io_diffCommits_info_138_fpWen ),
    .io_diffCommits_info_138_vecWen ( io_diffCommits_info_138_vecWen ),
    .io_diffCommits_info_138_v0Wen ( io_diffCommits_info_138_v0Wen ),
    .io_diffCommits_info_138_vlWen ( io_diffCommits_info_138_vlWen ),
    .io_diffCommits_info_139_ldest ( io_diffCommits_info_139_ldest ),
    .io_diffCommits_info_139_pdest ( io_diffCommits_info_139_pdest ),
    .io_diffCommits_info_139_rfWen ( io_diffCommits_info_139_rfWen ),
    .io_diffCommits_info_139_fpWen ( io_diffCommits_info_139_fpWen ),
    .io_diffCommits_info_139_vecWen ( io_diffCommits_info_139_vecWen ),
    .io_diffCommits_info_139_v0Wen ( io_diffCommits_info_139_v0Wen ),
    .io_diffCommits_info_139_vlWen ( io_diffCommits_info_139_vlWen ),
    .io_diffCommits_info_140_ldest ( io_diffCommits_info_140_ldest ),
    .io_diffCommits_info_140_pdest ( io_diffCommits_info_140_pdest ),
    .io_diffCommits_info_140_rfWen ( io_diffCommits_info_140_rfWen ),
    .io_diffCommits_info_140_fpWen ( io_diffCommits_info_140_fpWen ),
    .io_diffCommits_info_140_vecWen ( io_diffCommits_info_140_vecWen ),
    .io_diffCommits_info_140_v0Wen ( io_diffCommits_info_140_v0Wen ),
    .io_diffCommits_info_140_vlWen ( io_diffCommits_info_140_vlWen ),
    .io_diffCommits_info_141_ldest ( io_diffCommits_info_141_ldest ),
    .io_diffCommits_info_141_pdest ( io_diffCommits_info_141_pdest ),
    .io_diffCommits_info_141_rfWen ( io_diffCommits_info_141_rfWen ),
    .io_diffCommits_info_141_fpWen ( io_diffCommits_info_141_fpWen ),
    .io_diffCommits_info_141_vecWen ( io_diffCommits_info_141_vecWen ),
    .io_diffCommits_info_141_v0Wen ( io_diffCommits_info_141_v0Wen ),
    .io_diffCommits_info_141_vlWen ( io_diffCommits_info_141_vlWen ),
    .io_diffCommits_info_142_ldest ( io_diffCommits_info_142_ldest ),
    .io_diffCommits_info_142_pdest ( io_diffCommits_info_142_pdest ),
    .io_diffCommits_info_142_rfWen ( io_diffCommits_info_142_rfWen ),
    .io_diffCommits_info_142_fpWen ( io_diffCommits_info_142_fpWen ),
    .io_diffCommits_info_142_vecWen ( io_diffCommits_info_142_vecWen ),
    .io_diffCommits_info_142_v0Wen ( io_diffCommits_info_142_v0Wen ),
    .io_diffCommits_info_142_vlWen ( io_diffCommits_info_142_vlWen ),
    .io_diffCommits_info_143_ldest ( io_diffCommits_info_143_ldest ),
    .io_diffCommits_info_143_pdest ( io_diffCommits_info_143_pdest ),
    .io_diffCommits_info_143_rfWen ( io_diffCommits_info_143_rfWen ),
    .io_diffCommits_info_143_fpWen ( io_diffCommits_info_143_fpWen ),
    .io_diffCommits_info_143_vecWen ( io_diffCommits_info_143_vecWen ),
    .io_diffCommits_info_143_v0Wen ( io_diffCommits_info_143_v0Wen ),
    .io_diffCommits_info_143_vlWen ( io_diffCommits_info_143_vlWen ),
    .io_diffCommits_info_144_ldest ( io_diffCommits_info_144_ldest ),
    .io_diffCommits_info_144_pdest ( io_diffCommits_info_144_pdest ),
    .io_diffCommits_info_144_rfWen ( io_diffCommits_info_144_rfWen ),
    .io_diffCommits_info_144_fpWen ( io_diffCommits_info_144_fpWen ),
    .io_diffCommits_info_144_vecWen ( io_diffCommits_info_144_vecWen ),
    .io_diffCommits_info_144_v0Wen ( io_diffCommits_info_144_v0Wen ),
    .io_diffCommits_info_144_vlWen ( io_diffCommits_info_144_vlWen ),
    .io_diffCommits_info_145_ldest ( io_diffCommits_info_145_ldest ),
    .io_diffCommits_info_145_pdest ( io_diffCommits_info_145_pdest ),
    .io_diffCommits_info_145_rfWen ( io_diffCommits_info_145_rfWen ),
    .io_diffCommits_info_145_fpWen ( io_diffCommits_info_145_fpWen ),
    .io_diffCommits_info_145_vecWen ( io_diffCommits_info_145_vecWen ),
    .io_diffCommits_info_145_v0Wen ( io_diffCommits_info_145_v0Wen ),
    .io_diffCommits_info_145_vlWen ( io_diffCommits_info_145_vlWen ),
    .io_diffCommits_info_146_ldest ( io_diffCommits_info_146_ldest ),
    .io_diffCommits_info_146_pdest ( io_diffCommits_info_146_pdest ),
    .io_diffCommits_info_146_rfWen ( io_diffCommits_info_146_rfWen ),
    .io_diffCommits_info_146_fpWen ( io_diffCommits_info_146_fpWen ),
    .io_diffCommits_info_146_vecWen ( io_diffCommits_info_146_vecWen ),
    .io_diffCommits_info_146_v0Wen ( io_diffCommits_info_146_v0Wen ),
    .io_diffCommits_info_146_vlWen ( io_diffCommits_info_146_vlWen ),
    .io_diffCommits_info_147_ldest ( io_diffCommits_info_147_ldest ),
    .io_diffCommits_info_147_pdest ( io_diffCommits_info_147_pdest ),
    .io_diffCommits_info_147_rfWen ( io_diffCommits_info_147_rfWen ),
    .io_diffCommits_info_147_fpWen ( io_diffCommits_info_147_fpWen ),
    .io_diffCommits_info_147_vecWen ( io_diffCommits_info_147_vecWen ),
    .io_diffCommits_info_147_v0Wen ( io_diffCommits_info_147_v0Wen ),
    .io_diffCommits_info_147_vlWen ( io_diffCommits_info_147_vlWen ),
    .io_diffCommits_info_148_ldest ( io_diffCommits_info_148_ldest ),
    .io_diffCommits_info_148_pdest ( io_diffCommits_info_148_pdest ),
    .io_diffCommits_info_148_rfWen ( io_diffCommits_info_148_rfWen ),
    .io_diffCommits_info_148_fpWen ( io_diffCommits_info_148_fpWen ),
    .io_diffCommits_info_148_vecWen ( io_diffCommits_info_148_vecWen ),
    .io_diffCommits_info_148_v0Wen ( io_diffCommits_info_148_v0Wen ),
    .io_diffCommits_info_148_vlWen ( io_diffCommits_info_148_vlWen ),
    .io_diffCommits_info_149_ldest ( io_diffCommits_info_149_ldest ),
    .io_diffCommits_info_149_pdest ( io_diffCommits_info_149_pdest ),
    .io_diffCommits_info_149_rfWen ( io_diffCommits_info_149_rfWen ),
    .io_diffCommits_info_149_fpWen ( io_diffCommits_info_149_fpWen ),
    .io_diffCommits_info_149_vecWen ( io_diffCommits_info_149_vecWen ),
    .io_diffCommits_info_149_v0Wen ( io_diffCommits_info_149_v0Wen ),
    .io_diffCommits_info_149_vlWen ( io_diffCommits_info_149_vlWen ),
    .io_diffCommits_info_150_ldest ( io_diffCommits_info_150_ldest ),
    .io_diffCommits_info_150_pdest ( io_diffCommits_info_150_pdest ),
    .io_diffCommits_info_150_rfWen ( io_diffCommits_info_150_rfWen ),
    .io_diffCommits_info_150_fpWen ( io_diffCommits_info_150_fpWen ),
    .io_diffCommits_info_150_vecWen ( io_diffCommits_info_150_vecWen ),
    .io_diffCommits_info_150_v0Wen ( io_diffCommits_info_150_v0Wen ),
    .io_diffCommits_info_150_vlWen ( io_diffCommits_info_150_vlWen ),
    .io_diffCommits_info_151_ldest ( io_diffCommits_info_151_ldest ),
    .io_diffCommits_info_151_pdest ( io_diffCommits_info_151_pdest ),
    .io_diffCommits_info_151_rfWen ( io_diffCommits_info_151_rfWen ),
    .io_diffCommits_info_151_fpWen ( io_diffCommits_info_151_fpWen ),
    .io_diffCommits_info_151_vecWen ( io_diffCommits_info_151_vecWen ),
    .io_diffCommits_info_151_v0Wen ( io_diffCommits_info_151_v0Wen ),
    .io_diffCommits_info_151_vlWen ( io_diffCommits_info_151_vlWen ),
    .io_diffCommits_info_152_ldest ( io_diffCommits_info_152_ldest ),
    .io_diffCommits_info_152_pdest ( io_diffCommits_info_152_pdest ),
    .io_diffCommits_info_152_rfWen ( io_diffCommits_info_152_rfWen ),
    .io_diffCommits_info_152_fpWen ( io_diffCommits_info_152_fpWen ),
    .io_diffCommits_info_152_vecWen ( io_diffCommits_info_152_vecWen ),
    .io_diffCommits_info_152_v0Wen ( io_diffCommits_info_152_v0Wen ),
    .io_diffCommits_info_152_vlWen ( io_diffCommits_info_152_vlWen ),
    .io_diffCommits_info_153_ldest ( io_diffCommits_info_153_ldest ),
    .io_diffCommits_info_153_pdest ( io_diffCommits_info_153_pdest ),
    .io_diffCommits_info_153_rfWen ( io_diffCommits_info_153_rfWen ),
    .io_diffCommits_info_153_fpWen ( io_diffCommits_info_153_fpWen ),
    .io_diffCommits_info_153_vecWen ( io_diffCommits_info_153_vecWen ),
    .io_diffCommits_info_153_v0Wen ( io_diffCommits_info_153_v0Wen ),
    .io_diffCommits_info_153_vlWen ( io_diffCommits_info_153_vlWen ),
    .io_diffCommits_info_154_ldest ( io_diffCommits_info_154_ldest ),
    .io_diffCommits_info_154_pdest ( io_diffCommits_info_154_pdest ),
    .io_diffCommits_info_154_rfWen ( io_diffCommits_info_154_rfWen ),
    .io_diffCommits_info_154_fpWen ( io_diffCommits_info_154_fpWen ),
    .io_diffCommits_info_154_vecWen ( io_diffCommits_info_154_vecWen ),
    .io_diffCommits_info_154_v0Wen ( io_diffCommits_info_154_v0Wen ),
    .io_diffCommits_info_154_vlWen ( io_diffCommits_info_154_vlWen ),
    .io_diffCommits_info_155_ldest ( io_diffCommits_info_155_ldest ),
    .io_diffCommits_info_155_pdest ( io_diffCommits_info_155_pdest ),
    .io_diffCommits_info_155_rfWen ( io_diffCommits_info_155_rfWen ),
    .io_diffCommits_info_155_fpWen ( io_diffCommits_info_155_fpWen ),
    .io_diffCommits_info_155_vecWen ( io_diffCommits_info_155_vecWen ),
    .io_diffCommits_info_155_v0Wen ( io_diffCommits_info_155_v0Wen ),
    .io_diffCommits_info_155_vlWen ( io_diffCommits_info_155_vlWen ),
    .io_diffCommits_info_156_ldest ( io_diffCommits_info_156_ldest ),
    .io_diffCommits_info_156_pdest ( io_diffCommits_info_156_pdest ),
    .io_diffCommits_info_156_rfWen ( io_diffCommits_info_156_rfWen ),
    .io_diffCommits_info_156_fpWen ( io_diffCommits_info_156_fpWen ),
    .io_diffCommits_info_156_vecWen ( io_diffCommits_info_156_vecWen ),
    .io_diffCommits_info_156_v0Wen ( io_diffCommits_info_156_v0Wen ),
    .io_diffCommits_info_156_vlWen ( io_diffCommits_info_156_vlWen ),
    .io_diffCommits_info_157_ldest ( io_diffCommits_info_157_ldest ),
    .io_diffCommits_info_157_pdest ( io_diffCommits_info_157_pdest ),
    .io_diffCommits_info_157_rfWen ( io_diffCommits_info_157_rfWen ),
    .io_diffCommits_info_157_fpWen ( io_diffCommits_info_157_fpWen ),
    .io_diffCommits_info_157_vecWen ( io_diffCommits_info_157_vecWen ),
    .io_diffCommits_info_157_v0Wen ( io_diffCommits_info_157_v0Wen ),
    .io_diffCommits_info_157_vlWen ( io_diffCommits_info_157_vlWen ),
    .io_diffCommits_info_158_ldest ( io_diffCommits_info_158_ldest ),
    .io_diffCommits_info_158_pdest ( io_diffCommits_info_158_pdest ),
    .io_diffCommits_info_158_rfWen ( io_diffCommits_info_158_rfWen ),
    .io_diffCommits_info_158_fpWen ( io_diffCommits_info_158_fpWen ),
    .io_diffCommits_info_158_vecWen ( io_diffCommits_info_158_vecWen ),
    .io_diffCommits_info_158_v0Wen ( io_diffCommits_info_158_v0Wen ),
    .io_diffCommits_info_158_vlWen ( io_diffCommits_info_158_vlWen ),
    .io_diffCommits_info_159_ldest ( io_diffCommits_info_159_ldest ),
    .io_diffCommits_info_159_pdest ( io_diffCommits_info_159_pdest ),
    .io_diffCommits_info_159_rfWen ( io_diffCommits_info_159_rfWen ),
    .io_diffCommits_info_159_fpWen ( io_diffCommits_info_159_fpWen ),
    .io_diffCommits_info_159_vecWen ( io_diffCommits_info_159_vecWen ),
    .io_diffCommits_info_159_v0Wen ( io_diffCommits_info_159_v0Wen ),
    .io_diffCommits_info_159_vlWen ( io_diffCommits_info_159_vlWen ),
    .io_diffCommits_info_160_ldest ( io_diffCommits_info_160_ldest ),
    .io_diffCommits_info_160_pdest ( io_diffCommits_info_160_pdest ),
    .io_diffCommits_info_160_rfWen ( io_diffCommits_info_160_rfWen ),
    .io_diffCommits_info_160_fpWen ( io_diffCommits_info_160_fpWen ),
    .io_diffCommits_info_160_vecWen ( io_diffCommits_info_160_vecWen ),
    .io_diffCommits_info_160_v0Wen ( io_diffCommits_info_160_v0Wen ),
    .io_diffCommits_info_160_vlWen ( io_diffCommits_info_160_vlWen ),
    .io_diffCommits_info_161_ldest ( io_diffCommits_info_161_ldest ),
    .io_diffCommits_info_161_pdest ( io_diffCommits_info_161_pdest ),
    .io_diffCommits_info_161_rfWen ( io_diffCommits_info_161_rfWen ),
    .io_diffCommits_info_161_fpWen ( io_diffCommits_info_161_fpWen ),
    .io_diffCommits_info_161_vecWen ( io_diffCommits_info_161_vecWen ),
    .io_diffCommits_info_161_v0Wen ( io_diffCommits_info_161_v0Wen ),
    .io_diffCommits_info_161_vlWen ( io_diffCommits_info_161_vlWen ),
    .io_diffCommits_info_162_ldest ( io_diffCommits_info_162_ldest ),
    .io_diffCommits_info_162_pdest ( io_diffCommits_info_162_pdest ),
    .io_diffCommits_info_162_rfWen ( io_diffCommits_info_162_rfWen ),
    .io_diffCommits_info_162_fpWen ( io_diffCommits_info_162_fpWen ),
    .io_diffCommits_info_162_vecWen ( io_diffCommits_info_162_vecWen ),
    .io_diffCommits_info_162_v0Wen ( io_diffCommits_info_162_v0Wen ),
    .io_diffCommits_info_162_vlWen ( io_diffCommits_info_162_vlWen ),
    .io_diffCommits_info_163_ldest ( io_diffCommits_info_163_ldest ),
    .io_diffCommits_info_163_pdest ( io_diffCommits_info_163_pdest ),
    .io_diffCommits_info_163_rfWen ( io_diffCommits_info_163_rfWen ),
    .io_diffCommits_info_163_fpWen ( io_diffCommits_info_163_fpWen ),
    .io_diffCommits_info_163_vecWen ( io_diffCommits_info_163_vecWen ),
    .io_diffCommits_info_163_v0Wen ( io_diffCommits_info_163_v0Wen ),
    .io_diffCommits_info_163_vlWen ( io_diffCommits_info_163_vlWen ),
    .io_diffCommits_info_164_ldest ( io_diffCommits_info_164_ldest ),
    .io_diffCommits_info_164_pdest ( io_diffCommits_info_164_pdest ),
    .io_diffCommits_info_164_rfWen ( io_diffCommits_info_164_rfWen ),
    .io_diffCommits_info_164_fpWen ( io_diffCommits_info_164_fpWen ),
    .io_diffCommits_info_164_vecWen ( io_diffCommits_info_164_vecWen ),
    .io_diffCommits_info_164_v0Wen ( io_diffCommits_info_164_v0Wen ),
    .io_diffCommits_info_164_vlWen ( io_diffCommits_info_164_vlWen ),
    .io_diffCommits_info_165_ldest ( io_diffCommits_info_165_ldest ),
    .io_diffCommits_info_165_pdest ( io_diffCommits_info_165_pdest ),
    .io_diffCommits_info_165_rfWen ( io_diffCommits_info_165_rfWen ),
    .io_diffCommits_info_165_fpWen ( io_diffCommits_info_165_fpWen ),
    .io_diffCommits_info_165_vecWen ( io_diffCommits_info_165_vecWen ),
    .io_diffCommits_info_165_v0Wen ( io_diffCommits_info_165_v0Wen ),
    .io_diffCommits_info_165_vlWen ( io_diffCommits_info_165_vlWen ),
    .io_diffCommits_info_166_ldest ( io_diffCommits_info_166_ldest ),
    .io_diffCommits_info_166_pdest ( io_diffCommits_info_166_pdest ),
    .io_diffCommits_info_166_rfWen ( io_diffCommits_info_166_rfWen ),
    .io_diffCommits_info_166_fpWen ( io_diffCommits_info_166_fpWen ),
    .io_diffCommits_info_166_vecWen ( io_diffCommits_info_166_vecWen ),
    .io_diffCommits_info_166_v0Wen ( io_diffCommits_info_166_v0Wen ),
    .io_diffCommits_info_166_vlWen ( io_diffCommits_info_166_vlWen ),
    .io_diffCommits_info_167_ldest ( io_diffCommits_info_167_ldest ),
    .io_diffCommits_info_167_pdest ( io_diffCommits_info_167_pdest ),
    .io_diffCommits_info_167_rfWen ( io_diffCommits_info_167_rfWen ),
    .io_diffCommits_info_167_fpWen ( io_diffCommits_info_167_fpWen ),
    .io_diffCommits_info_167_vecWen ( io_diffCommits_info_167_vecWen ),
    .io_diffCommits_info_167_v0Wen ( io_diffCommits_info_167_v0Wen ),
    .io_diffCommits_info_167_vlWen ( io_diffCommits_info_167_vlWen ),
    .io_diffCommits_info_168_ldest ( io_diffCommits_info_168_ldest ),
    .io_diffCommits_info_168_pdest ( io_diffCommits_info_168_pdest ),
    .io_diffCommits_info_168_rfWen ( io_diffCommits_info_168_rfWen ),
    .io_diffCommits_info_168_fpWen ( io_diffCommits_info_168_fpWen ),
    .io_diffCommits_info_168_vecWen ( io_diffCommits_info_168_vecWen ),
    .io_diffCommits_info_168_v0Wen ( io_diffCommits_info_168_v0Wen ),
    .io_diffCommits_info_168_vlWen ( io_diffCommits_info_168_vlWen ),
    .io_diffCommits_info_169_ldest ( io_diffCommits_info_169_ldest ),
    .io_diffCommits_info_169_pdest ( io_diffCommits_info_169_pdest ),
    .io_diffCommits_info_169_rfWen ( io_diffCommits_info_169_rfWen ),
    .io_diffCommits_info_169_fpWen ( io_diffCommits_info_169_fpWen ),
    .io_diffCommits_info_169_vecWen ( io_diffCommits_info_169_vecWen ),
    .io_diffCommits_info_169_v0Wen ( io_diffCommits_info_169_v0Wen ),
    .io_diffCommits_info_169_vlWen ( io_diffCommits_info_169_vlWen ),
    .io_diffCommits_info_170_ldest ( io_diffCommits_info_170_ldest ),
    .io_diffCommits_info_170_pdest ( io_diffCommits_info_170_pdest ),
    .io_diffCommits_info_170_rfWen ( io_diffCommits_info_170_rfWen ),
    .io_diffCommits_info_170_fpWen ( io_diffCommits_info_170_fpWen ),
    .io_diffCommits_info_170_vecWen ( io_diffCommits_info_170_vecWen ),
    .io_diffCommits_info_170_v0Wen ( io_diffCommits_info_170_v0Wen ),
    .io_diffCommits_info_170_vlWen ( io_diffCommits_info_170_vlWen ),
    .io_diffCommits_info_171_ldest ( io_diffCommits_info_171_ldest ),
    .io_diffCommits_info_171_pdest ( io_diffCommits_info_171_pdest ),
    .io_diffCommits_info_171_rfWen ( io_diffCommits_info_171_rfWen ),
    .io_diffCommits_info_171_fpWen ( io_diffCommits_info_171_fpWen ),
    .io_diffCommits_info_171_vecWen ( io_diffCommits_info_171_vecWen ),
    .io_diffCommits_info_171_v0Wen ( io_diffCommits_info_171_v0Wen ),
    .io_diffCommits_info_171_vlWen ( io_diffCommits_info_171_vlWen ),
    .io_diffCommits_info_172_ldest ( io_diffCommits_info_172_ldest ),
    .io_diffCommits_info_172_pdest ( io_diffCommits_info_172_pdest ),
    .io_diffCommits_info_172_rfWen ( io_diffCommits_info_172_rfWen ),
    .io_diffCommits_info_172_fpWen ( io_diffCommits_info_172_fpWen ),
    .io_diffCommits_info_172_vecWen ( io_diffCommits_info_172_vecWen ),
    .io_diffCommits_info_172_v0Wen ( io_diffCommits_info_172_v0Wen ),
    .io_diffCommits_info_172_vlWen ( io_diffCommits_info_172_vlWen ),
    .io_diffCommits_info_173_ldest ( io_diffCommits_info_173_ldest ),
    .io_diffCommits_info_173_pdest ( io_diffCommits_info_173_pdest ),
    .io_diffCommits_info_173_rfWen ( io_diffCommits_info_173_rfWen ),
    .io_diffCommits_info_173_fpWen ( io_diffCommits_info_173_fpWen ),
    .io_diffCommits_info_173_vecWen ( io_diffCommits_info_173_vecWen ),
    .io_diffCommits_info_173_v0Wen ( io_diffCommits_info_173_v0Wen ),
    .io_diffCommits_info_173_vlWen ( io_diffCommits_info_173_vlWen ),
    .io_diffCommits_info_174_ldest ( io_diffCommits_info_174_ldest ),
    .io_diffCommits_info_174_pdest ( io_diffCommits_info_174_pdest ),
    .io_diffCommits_info_174_rfWen ( io_diffCommits_info_174_rfWen ),
    .io_diffCommits_info_174_fpWen ( io_diffCommits_info_174_fpWen ),
    .io_diffCommits_info_174_vecWen ( io_diffCommits_info_174_vecWen ),
    .io_diffCommits_info_174_v0Wen ( io_diffCommits_info_174_v0Wen ),
    .io_diffCommits_info_174_vlWen ( io_diffCommits_info_174_vlWen ),
    .io_diffCommits_info_175_ldest ( io_diffCommits_info_175_ldest ),
    .io_diffCommits_info_175_pdest ( io_diffCommits_info_175_pdest ),
    .io_diffCommits_info_175_rfWen ( io_diffCommits_info_175_rfWen ),
    .io_diffCommits_info_175_fpWen ( io_diffCommits_info_175_fpWen ),
    .io_diffCommits_info_175_vecWen ( io_diffCommits_info_175_vecWen ),
    .io_diffCommits_info_175_v0Wen ( io_diffCommits_info_175_v0Wen ),
    .io_diffCommits_info_175_vlWen ( io_diffCommits_info_175_vlWen ),
    .io_diffCommits_info_176_ldest ( io_diffCommits_info_176_ldest ),
    .io_diffCommits_info_176_pdest ( io_diffCommits_info_176_pdest ),
    .io_diffCommits_info_176_rfWen ( io_diffCommits_info_176_rfWen ),
    .io_diffCommits_info_176_fpWen ( io_diffCommits_info_176_fpWen ),
    .io_diffCommits_info_176_vecWen ( io_diffCommits_info_176_vecWen ),
    .io_diffCommits_info_176_v0Wen ( io_diffCommits_info_176_v0Wen ),
    .io_diffCommits_info_176_vlWen ( io_diffCommits_info_176_vlWen ),
    .io_diffCommits_info_177_ldest ( io_diffCommits_info_177_ldest ),
    .io_diffCommits_info_177_pdest ( io_diffCommits_info_177_pdest ),
    .io_diffCommits_info_177_rfWen ( io_diffCommits_info_177_rfWen ),
    .io_diffCommits_info_177_fpWen ( io_diffCommits_info_177_fpWen ),
    .io_diffCommits_info_177_vecWen ( io_diffCommits_info_177_vecWen ),
    .io_diffCommits_info_177_v0Wen ( io_diffCommits_info_177_v0Wen ),
    .io_diffCommits_info_177_vlWen ( io_diffCommits_info_177_vlWen ),
    .io_diffCommits_info_178_ldest ( io_diffCommits_info_178_ldest ),
    .io_diffCommits_info_178_pdest ( io_diffCommits_info_178_pdest ),
    .io_diffCommits_info_178_rfWen ( io_diffCommits_info_178_rfWen ),
    .io_diffCommits_info_178_fpWen ( io_diffCommits_info_178_fpWen ),
    .io_diffCommits_info_178_vecWen ( io_diffCommits_info_178_vecWen ),
    .io_diffCommits_info_178_v0Wen ( io_diffCommits_info_178_v0Wen ),
    .io_diffCommits_info_178_vlWen ( io_diffCommits_info_178_vlWen ),
    .io_diffCommits_info_179_ldest ( io_diffCommits_info_179_ldest ),
    .io_diffCommits_info_179_pdest ( io_diffCommits_info_179_pdest ),
    .io_diffCommits_info_179_rfWen ( io_diffCommits_info_179_rfWen ),
    .io_diffCommits_info_179_fpWen ( io_diffCommits_info_179_fpWen ),
    .io_diffCommits_info_179_vecWen ( io_diffCommits_info_179_vecWen ),
    .io_diffCommits_info_179_v0Wen ( io_diffCommits_info_179_v0Wen ),
    .io_diffCommits_info_179_vlWen ( io_diffCommits_info_179_vlWen ),
    .io_diffCommits_info_180_ldest ( io_diffCommits_info_180_ldest ),
    .io_diffCommits_info_180_pdest ( io_diffCommits_info_180_pdest ),
    .io_diffCommits_info_180_rfWen ( io_diffCommits_info_180_rfWen ),
    .io_diffCommits_info_180_fpWen ( io_diffCommits_info_180_fpWen ),
    .io_diffCommits_info_180_vecWen ( io_diffCommits_info_180_vecWen ),
    .io_diffCommits_info_180_v0Wen ( io_diffCommits_info_180_v0Wen ),
    .io_diffCommits_info_180_vlWen ( io_diffCommits_info_180_vlWen ),
    .io_diffCommits_info_181_ldest ( io_diffCommits_info_181_ldest ),
    .io_diffCommits_info_181_pdest ( io_diffCommits_info_181_pdest ),
    .io_diffCommits_info_181_rfWen ( io_diffCommits_info_181_rfWen ),
    .io_diffCommits_info_181_fpWen ( io_diffCommits_info_181_fpWen ),
    .io_diffCommits_info_181_vecWen ( io_diffCommits_info_181_vecWen ),
    .io_diffCommits_info_181_v0Wen ( io_diffCommits_info_181_v0Wen ),
    .io_diffCommits_info_181_vlWen ( io_diffCommits_info_181_vlWen ),
    .io_diffCommits_info_182_ldest ( io_diffCommits_info_182_ldest ),
    .io_diffCommits_info_182_pdest ( io_diffCommits_info_182_pdest ),
    .io_diffCommits_info_182_rfWen ( io_diffCommits_info_182_rfWen ),
    .io_diffCommits_info_182_fpWen ( io_diffCommits_info_182_fpWen ),
    .io_diffCommits_info_182_vecWen ( io_diffCommits_info_182_vecWen ),
    .io_diffCommits_info_182_v0Wen ( io_diffCommits_info_182_v0Wen ),
    .io_diffCommits_info_182_vlWen ( io_diffCommits_info_182_vlWen ),
    .io_diffCommits_info_183_ldest ( io_diffCommits_info_183_ldest ),
    .io_diffCommits_info_183_pdest ( io_diffCommits_info_183_pdest ),
    .io_diffCommits_info_183_rfWen ( io_diffCommits_info_183_rfWen ),
    .io_diffCommits_info_183_fpWen ( io_diffCommits_info_183_fpWen ),
    .io_diffCommits_info_183_vecWen ( io_diffCommits_info_183_vecWen ),
    .io_diffCommits_info_183_v0Wen ( io_diffCommits_info_183_v0Wen ),
    .io_diffCommits_info_183_vlWen ( io_diffCommits_info_183_vlWen ),
    .io_diffCommits_info_184_ldest ( io_diffCommits_info_184_ldest ),
    .io_diffCommits_info_184_pdest ( io_diffCommits_info_184_pdest ),
    .io_diffCommits_info_184_rfWen ( io_diffCommits_info_184_rfWen ),
    .io_diffCommits_info_184_fpWen ( io_diffCommits_info_184_fpWen ),
    .io_diffCommits_info_184_vecWen ( io_diffCommits_info_184_vecWen ),
    .io_diffCommits_info_184_v0Wen ( io_diffCommits_info_184_v0Wen ),
    .io_diffCommits_info_184_vlWen ( io_diffCommits_info_184_vlWen ),
    .io_diffCommits_info_185_ldest ( io_diffCommits_info_185_ldest ),
    .io_diffCommits_info_185_pdest ( io_diffCommits_info_185_pdest ),
    .io_diffCommits_info_185_rfWen ( io_diffCommits_info_185_rfWen ),
    .io_diffCommits_info_185_fpWen ( io_diffCommits_info_185_fpWen ),
    .io_diffCommits_info_185_vecWen ( io_diffCommits_info_185_vecWen ),
    .io_diffCommits_info_185_v0Wen ( io_diffCommits_info_185_v0Wen ),
    .io_diffCommits_info_185_vlWen ( io_diffCommits_info_185_vlWen ),
    .io_diffCommits_info_186_ldest ( io_diffCommits_info_186_ldest ),
    .io_diffCommits_info_186_pdest ( io_diffCommits_info_186_pdest ),
    .io_diffCommits_info_186_rfWen ( io_diffCommits_info_186_rfWen ),
    .io_diffCommits_info_186_fpWen ( io_diffCommits_info_186_fpWen ),
    .io_diffCommits_info_186_vecWen ( io_diffCommits_info_186_vecWen ),
    .io_diffCommits_info_186_v0Wen ( io_diffCommits_info_186_v0Wen ),
    .io_diffCommits_info_186_vlWen ( io_diffCommits_info_186_vlWen ),
    .io_diffCommits_info_187_ldest ( io_diffCommits_info_187_ldest ),
    .io_diffCommits_info_187_pdest ( io_diffCommits_info_187_pdest ),
    .io_diffCommits_info_187_rfWen ( io_diffCommits_info_187_rfWen ),
    .io_diffCommits_info_187_fpWen ( io_diffCommits_info_187_fpWen ),
    .io_diffCommits_info_187_vecWen ( io_diffCommits_info_187_vecWen ),
    .io_diffCommits_info_187_v0Wen ( io_diffCommits_info_187_v0Wen ),
    .io_diffCommits_info_187_vlWen ( io_diffCommits_info_187_vlWen ),
    .io_diffCommits_info_188_ldest ( io_diffCommits_info_188_ldest ),
    .io_diffCommits_info_188_pdest ( io_diffCommits_info_188_pdest ),
    .io_diffCommits_info_188_rfWen ( io_diffCommits_info_188_rfWen ),
    .io_diffCommits_info_188_fpWen ( io_diffCommits_info_188_fpWen ),
    .io_diffCommits_info_188_vecWen ( io_diffCommits_info_188_vecWen ),
    .io_diffCommits_info_188_v0Wen ( io_diffCommits_info_188_v0Wen ),
    .io_diffCommits_info_188_vlWen ( io_diffCommits_info_188_vlWen ),
    .io_diffCommits_info_189_ldest ( io_diffCommits_info_189_ldest ),
    .io_diffCommits_info_189_pdest ( io_diffCommits_info_189_pdest ),
    .io_diffCommits_info_189_rfWen ( io_diffCommits_info_189_rfWen ),
    .io_diffCommits_info_189_fpWen ( io_diffCommits_info_189_fpWen ),
    .io_diffCommits_info_189_vecWen ( io_diffCommits_info_189_vecWen ),
    .io_diffCommits_info_189_v0Wen ( io_diffCommits_info_189_v0Wen ),
    .io_diffCommits_info_189_vlWen ( io_diffCommits_info_189_vlWen ),
    .io_diffCommits_info_190_ldest ( io_diffCommits_info_190_ldest ),
    .io_diffCommits_info_190_pdest ( io_diffCommits_info_190_pdest ),
    .io_diffCommits_info_190_rfWen ( io_diffCommits_info_190_rfWen ),
    .io_diffCommits_info_190_fpWen ( io_diffCommits_info_190_fpWen ),
    .io_diffCommits_info_190_vecWen ( io_diffCommits_info_190_vecWen ),
    .io_diffCommits_info_190_v0Wen ( io_diffCommits_info_190_v0Wen ),
    .io_diffCommits_info_190_vlWen ( io_diffCommits_info_190_vlWen ),
    .io_diffCommits_info_191_ldest ( io_diffCommits_info_191_ldest ),
    .io_diffCommits_info_191_pdest ( io_diffCommits_info_191_pdest ),
    .io_diffCommits_info_191_rfWen ( io_diffCommits_info_191_rfWen ),
    .io_diffCommits_info_191_fpWen ( io_diffCommits_info_191_fpWen ),
    .io_diffCommits_info_191_vecWen ( io_diffCommits_info_191_vecWen ),
    .io_diffCommits_info_191_v0Wen ( io_diffCommits_info_191_v0Wen ),
    .io_diffCommits_info_191_vlWen ( io_diffCommits_info_191_vlWen ),
    .io_diffCommits_info_192_ldest ( io_diffCommits_info_192_ldest ),
    .io_diffCommits_info_192_pdest ( io_diffCommits_info_192_pdest ),
    .io_diffCommits_info_192_rfWen ( io_diffCommits_info_192_rfWen ),
    .io_diffCommits_info_192_fpWen ( io_diffCommits_info_192_fpWen ),
    .io_diffCommits_info_192_vecWen ( io_diffCommits_info_192_vecWen ),
    .io_diffCommits_info_192_v0Wen ( io_diffCommits_info_192_v0Wen ),
    .io_diffCommits_info_192_vlWen ( io_diffCommits_info_192_vlWen ),
    .io_diffCommits_info_193_ldest ( io_diffCommits_info_193_ldest ),
    .io_diffCommits_info_193_pdest ( io_diffCommits_info_193_pdest ),
    .io_diffCommits_info_193_rfWen ( io_diffCommits_info_193_rfWen ),
    .io_diffCommits_info_193_fpWen ( io_diffCommits_info_193_fpWen ),
    .io_diffCommits_info_193_vecWen ( io_diffCommits_info_193_vecWen ),
    .io_diffCommits_info_193_v0Wen ( io_diffCommits_info_193_v0Wen ),
    .io_diffCommits_info_193_vlWen ( io_diffCommits_info_193_vlWen ),
    .io_diffCommits_info_194_ldest ( io_diffCommits_info_194_ldest ),
    .io_diffCommits_info_194_pdest ( io_diffCommits_info_194_pdest ),
    .io_diffCommits_info_194_rfWen ( io_diffCommits_info_194_rfWen ),
    .io_diffCommits_info_194_fpWen ( io_diffCommits_info_194_fpWen ),
    .io_diffCommits_info_194_vecWen ( io_diffCommits_info_194_vecWen ),
    .io_diffCommits_info_194_v0Wen ( io_diffCommits_info_194_v0Wen ),
    .io_diffCommits_info_194_vlWen ( io_diffCommits_info_194_vlWen ),
    .io_diffCommits_info_195_ldest ( io_diffCommits_info_195_ldest ),
    .io_diffCommits_info_195_pdest ( io_diffCommits_info_195_pdest ),
    .io_diffCommits_info_195_rfWen ( io_diffCommits_info_195_rfWen ),
    .io_diffCommits_info_195_fpWen ( io_diffCommits_info_195_fpWen ),
    .io_diffCommits_info_195_vecWen ( io_diffCommits_info_195_vecWen ),
    .io_diffCommits_info_195_v0Wen ( io_diffCommits_info_195_v0Wen ),
    .io_diffCommits_info_195_vlWen ( io_diffCommits_info_195_vlWen ),
    .io_diffCommits_info_196_ldest ( io_diffCommits_info_196_ldest ),
    .io_diffCommits_info_196_pdest ( io_diffCommits_info_196_pdest ),
    .io_diffCommits_info_196_rfWen ( io_diffCommits_info_196_rfWen ),
    .io_diffCommits_info_196_fpWen ( io_diffCommits_info_196_fpWen ),
    .io_diffCommits_info_196_vecWen ( io_diffCommits_info_196_vecWen ),
    .io_diffCommits_info_196_v0Wen ( io_diffCommits_info_196_v0Wen ),
    .io_diffCommits_info_196_vlWen ( io_diffCommits_info_196_vlWen ),
    .io_diffCommits_info_197_ldest ( io_diffCommits_info_197_ldest ),
    .io_diffCommits_info_197_pdest ( io_diffCommits_info_197_pdest ),
    .io_diffCommits_info_197_rfWen ( io_diffCommits_info_197_rfWen ),
    .io_diffCommits_info_197_fpWen ( io_diffCommits_info_197_fpWen ),
    .io_diffCommits_info_197_vecWen ( io_diffCommits_info_197_vecWen ),
    .io_diffCommits_info_197_v0Wen ( io_diffCommits_info_197_v0Wen ),
    .io_diffCommits_info_197_vlWen ( io_diffCommits_info_197_vlWen ),
    .io_diffCommits_info_198_ldest ( io_diffCommits_info_198_ldest ),
    .io_diffCommits_info_198_pdest ( io_diffCommits_info_198_pdest ),
    .io_diffCommits_info_198_rfWen ( io_diffCommits_info_198_rfWen ),
    .io_diffCommits_info_198_fpWen ( io_diffCommits_info_198_fpWen ),
    .io_diffCommits_info_198_vecWen ( io_diffCommits_info_198_vecWen ),
    .io_diffCommits_info_198_v0Wen ( io_diffCommits_info_198_v0Wen ),
    .io_diffCommits_info_198_vlWen ( io_diffCommits_info_198_vlWen ),
    .io_diffCommits_info_199_ldest ( io_diffCommits_info_199_ldest ),
    .io_diffCommits_info_199_pdest ( io_diffCommits_info_199_pdest ),
    .io_diffCommits_info_199_rfWen ( io_diffCommits_info_199_rfWen ),
    .io_diffCommits_info_199_fpWen ( io_diffCommits_info_199_fpWen ),
    .io_diffCommits_info_199_vecWen ( io_diffCommits_info_199_vecWen ),
    .io_diffCommits_info_199_v0Wen ( io_diffCommits_info_199_v0Wen ),
    .io_diffCommits_info_199_vlWen ( io_diffCommits_info_199_vlWen ),
    .io_diffCommits_info_200_ldest ( io_diffCommits_info_200_ldest ),
    .io_diffCommits_info_200_pdest ( io_diffCommits_info_200_pdest ),
    .io_diffCommits_info_200_rfWen ( io_diffCommits_info_200_rfWen ),
    .io_diffCommits_info_200_fpWen ( io_diffCommits_info_200_fpWen ),
    .io_diffCommits_info_200_vecWen ( io_diffCommits_info_200_vecWen ),
    .io_diffCommits_info_200_v0Wen ( io_diffCommits_info_200_v0Wen ),
    .io_diffCommits_info_200_vlWen ( io_diffCommits_info_200_vlWen ),
    .io_diffCommits_info_201_ldest ( io_diffCommits_info_201_ldest ),
    .io_diffCommits_info_201_pdest ( io_diffCommits_info_201_pdest ),
    .io_diffCommits_info_201_rfWen ( io_diffCommits_info_201_rfWen ),
    .io_diffCommits_info_201_fpWen ( io_diffCommits_info_201_fpWen ),
    .io_diffCommits_info_201_vecWen ( io_diffCommits_info_201_vecWen ),
    .io_diffCommits_info_201_v0Wen ( io_diffCommits_info_201_v0Wen ),
    .io_diffCommits_info_201_vlWen ( io_diffCommits_info_201_vlWen ),
    .io_diffCommits_info_202_ldest ( io_diffCommits_info_202_ldest ),
    .io_diffCommits_info_202_pdest ( io_diffCommits_info_202_pdest ),
    .io_diffCommits_info_202_rfWen ( io_diffCommits_info_202_rfWen ),
    .io_diffCommits_info_202_fpWen ( io_diffCommits_info_202_fpWen ),
    .io_diffCommits_info_202_vecWen ( io_diffCommits_info_202_vecWen ),
    .io_diffCommits_info_202_v0Wen ( io_diffCommits_info_202_v0Wen ),
    .io_diffCommits_info_202_vlWen ( io_diffCommits_info_202_vlWen ),
    .io_diffCommits_info_203_ldest ( io_diffCommits_info_203_ldest ),
    .io_diffCommits_info_203_pdest ( io_diffCommits_info_203_pdest ),
    .io_diffCommits_info_203_rfWen ( io_diffCommits_info_203_rfWen ),
    .io_diffCommits_info_203_fpWen ( io_diffCommits_info_203_fpWen ),
    .io_diffCommits_info_203_vecWen ( io_diffCommits_info_203_vecWen ),
    .io_diffCommits_info_203_v0Wen ( io_diffCommits_info_203_v0Wen ),
    .io_diffCommits_info_203_vlWen ( io_diffCommits_info_203_vlWen ),
    .io_diffCommits_info_204_ldest ( io_diffCommits_info_204_ldest ),
    .io_diffCommits_info_204_pdest ( io_diffCommits_info_204_pdest ),
    .io_diffCommits_info_204_rfWen ( io_diffCommits_info_204_rfWen ),
    .io_diffCommits_info_204_fpWen ( io_diffCommits_info_204_fpWen ),
    .io_diffCommits_info_204_vecWen ( io_diffCommits_info_204_vecWen ),
    .io_diffCommits_info_204_v0Wen ( io_diffCommits_info_204_v0Wen ),
    .io_diffCommits_info_204_vlWen ( io_diffCommits_info_204_vlWen ),
    .io_diffCommits_info_205_ldest ( io_diffCommits_info_205_ldest ),
    .io_diffCommits_info_205_pdest ( io_diffCommits_info_205_pdest ),
    .io_diffCommits_info_205_rfWen ( io_diffCommits_info_205_rfWen ),
    .io_diffCommits_info_205_fpWen ( io_diffCommits_info_205_fpWen ),
    .io_diffCommits_info_205_vecWen ( io_diffCommits_info_205_vecWen ),
    .io_diffCommits_info_205_v0Wen ( io_diffCommits_info_205_v0Wen ),
    .io_diffCommits_info_205_vlWen ( io_diffCommits_info_205_vlWen ),
    .io_diffCommits_info_206_ldest ( io_diffCommits_info_206_ldest ),
    .io_diffCommits_info_206_pdest ( io_diffCommits_info_206_pdest ),
    .io_diffCommits_info_206_rfWen ( io_diffCommits_info_206_rfWen ),
    .io_diffCommits_info_206_fpWen ( io_diffCommits_info_206_fpWen ),
    .io_diffCommits_info_206_vecWen ( io_diffCommits_info_206_vecWen ),
    .io_diffCommits_info_206_v0Wen ( io_diffCommits_info_206_v0Wen ),
    .io_diffCommits_info_206_vlWen ( io_diffCommits_info_206_vlWen ),
    .io_diffCommits_info_207_ldest ( io_diffCommits_info_207_ldest ),
    .io_diffCommits_info_207_pdest ( io_diffCommits_info_207_pdest ),
    .io_diffCommits_info_207_rfWen ( io_diffCommits_info_207_rfWen ),
    .io_diffCommits_info_207_fpWen ( io_diffCommits_info_207_fpWen ),
    .io_diffCommits_info_207_vecWen ( io_diffCommits_info_207_vecWen ),
    .io_diffCommits_info_207_v0Wen ( io_diffCommits_info_207_v0Wen ),
    .io_diffCommits_info_207_vlWen ( io_diffCommits_info_207_vlWen ),
    .io_diffCommits_info_208_ldest ( io_diffCommits_info_208_ldest ),
    .io_diffCommits_info_208_pdest ( io_diffCommits_info_208_pdest ),
    .io_diffCommits_info_208_rfWen ( io_diffCommits_info_208_rfWen ),
    .io_diffCommits_info_208_fpWen ( io_diffCommits_info_208_fpWen ),
    .io_diffCommits_info_208_vecWen ( io_diffCommits_info_208_vecWen ),
    .io_diffCommits_info_208_v0Wen ( io_diffCommits_info_208_v0Wen ),
    .io_diffCommits_info_208_vlWen ( io_diffCommits_info_208_vlWen ),
    .io_diffCommits_info_209_ldest ( io_diffCommits_info_209_ldest ),
    .io_diffCommits_info_209_pdest ( io_diffCommits_info_209_pdest ),
    .io_diffCommits_info_209_rfWen ( io_diffCommits_info_209_rfWen ),
    .io_diffCommits_info_209_fpWen ( io_diffCommits_info_209_fpWen ),
    .io_diffCommits_info_209_vecWen ( io_diffCommits_info_209_vecWen ),
    .io_diffCommits_info_209_v0Wen ( io_diffCommits_info_209_v0Wen ),
    .io_diffCommits_info_209_vlWen ( io_diffCommits_info_209_vlWen ),
    .io_diffCommits_info_210_ldest ( io_diffCommits_info_210_ldest ),
    .io_diffCommits_info_210_pdest ( io_diffCommits_info_210_pdest ),
    .io_diffCommits_info_210_rfWen ( io_diffCommits_info_210_rfWen ),
    .io_diffCommits_info_210_fpWen ( io_diffCommits_info_210_fpWen ),
    .io_diffCommits_info_210_vecWen ( io_diffCommits_info_210_vecWen ),
    .io_diffCommits_info_210_v0Wen ( io_diffCommits_info_210_v0Wen ),
    .io_diffCommits_info_210_vlWen ( io_diffCommits_info_210_vlWen ),
    .io_diffCommits_info_211_ldest ( io_diffCommits_info_211_ldest ),
    .io_diffCommits_info_211_pdest ( io_diffCommits_info_211_pdest ),
    .io_diffCommits_info_211_rfWen ( io_diffCommits_info_211_rfWen ),
    .io_diffCommits_info_211_fpWen ( io_diffCommits_info_211_fpWen ),
    .io_diffCommits_info_211_vecWen ( io_diffCommits_info_211_vecWen ),
    .io_diffCommits_info_211_v0Wen ( io_diffCommits_info_211_v0Wen ),
    .io_diffCommits_info_211_vlWen ( io_diffCommits_info_211_vlWen ),
    .io_diffCommits_info_212_ldest ( io_diffCommits_info_212_ldest ),
    .io_diffCommits_info_212_pdest ( io_diffCommits_info_212_pdest ),
    .io_diffCommits_info_212_rfWen ( io_diffCommits_info_212_rfWen ),
    .io_diffCommits_info_212_fpWen ( io_diffCommits_info_212_fpWen ),
    .io_diffCommits_info_212_vecWen ( io_diffCommits_info_212_vecWen ),
    .io_diffCommits_info_212_v0Wen ( io_diffCommits_info_212_v0Wen ),
    .io_diffCommits_info_212_vlWen ( io_diffCommits_info_212_vlWen ),
    .io_diffCommits_info_213_ldest ( io_diffCommits_info_213_ldest ),
    .io_diffCommits_info_213_pdest ( io_diffCommits_info_213_pdest ),
    .io_diffCommits_info_213_rfWen ( io_diffCommits_info_213_rfWen ),
    .io_diffCommits_info_213_fpWen ( io_diffCommits_info_213_fpWen ),
    .io_diffCommits_info_213_vecWen ( io_diffCommits_info_213_vecWen ),
    .io_diffCommits_info_213_v0Wen ( io_diffCommits_info_213_v0Wen ),
    .io_diffCommits_info_213_vlWen ( io_diffCommits_info_213_vlWen ),
    .io_diffCommits_info_214_ldest ( io_diffCommits_info_214_ldest ),
    .io_diffCommits_info_214_pdest ( io_diffCommits_info_214_pdest ),
    .io_diffCommits_info_214_rfWen ( io_diffCommits_info_214_rfWen ),
    .io_diffCommits_info_214_fpWen ( io_diffCommits_info_214_fpWen ),
    .io_diffCommits_info_214_vecWen ( io_diffCommits_info_214_vecWen ),
    .io_diffCommits_info_214_v0Wen ( io_diffCommits_info_214_v0Wen ),
    .io_diffCommits_info_214_vlWen ( io_diffCommits_info_214_vlWen ),
    .io_diffCommits_info_215_ldest ( io_diffCommits_info_215_ldest ),
    .io_diffCommits_info_215_pdest ( io_diffCommits_info_215_pdest ),
    .io_diffCommits_info_215_rfWen ( io_diffCommits_info_215_rfWen ),
    .io_diffCommits_info_215_fpWen ( io_diffCommits_info_215_fpWen ),
    .io_diffCommits_info_215_vecWen ( io_diffCommits_info_215_vecWen ),
    .io_diffCommits_info_215_v0Wen ( io_diffCommits_info_215_v0Wen ),
    .io_diffCommits_info_215_vlWen ( io_diffCommits_info_215_vlWen ),
    .io_diffCommits_info_216_ldest ( io_diffCommits_info_216_ldest ),
    .io_diffCommits_info_216_pdest ( io_diffCommits_info_216_pdest ),
    .io_diffCommits_info_216_rfWen ( io_diffCommits_info_216_rfWen ),
    .io_diffCommits_info_216_fpWen ( io_diffCommits_info_216_fpWen ),
    .io_diffCommits_info_216_vecWen ( io_diffCommits_info_216_vecWen ),
    .io_diffCommits_info_216_v0Wen ( io_diffCommits_info_216_v0Wen ),
    .io_diffCommits_info_216_vlWen ( io_diffCommits_info_216_vlWen ),
    .io_diffCommits_info_217_ldest ( io_diffCommits_info_217_ldest ),
    .io_diffCommits_info_217_pdest ( io_diffCommits_info_217_pdest ),
    .io_diffCommits_info_217_rfWen ( io_diffCommits_info_217_rfWen ),
    .io_diffCommits_info_217_fpWen ( io_diffCommits_info_217_fpWen ),
    .io_diffCommits_info_217_vecWen ( io_diffCommits_info_217_vecWen ),
    .io_diffCommits_info_217_v0Wen ( io_diffCommits_info_217_v0Wen ),
    .io_diffCommits_info_217_vlWen ( io_diffCommits_info_217_vlWen ),
    .io_diffCommits_info_218_ldest ( io_diffCommits_info_218_ldest ),
    .io_diffCommits_info_218_pdest ( io_diffCommits_info_218_pdest ),
    .io_diffCommits_info_218_rfWen ( io_diffCommits_info_218_rfWen ),
    .io_diffCommits_info_218_fpWen ( io_diffCommits_info_218_fpWen ),
    .io_diffCommits_info_218_vecWen ( io_diffCommits_info_218_vecWen ),
    .io_diffCommits_info_218_v0Wen ( io_diffCommits_info_218_v0Wen ),
    .io_diffCommits_info_218_vlWen ( io_diffCommits_info_218_vlWen ),
    .io_diffCommits_info_219_ldest ( io_diffCommits_info_219_ldest ),
    .io_diffCommits_info_219_pdest ( io_diffCommits_info_219_pdest ),
    .io_diffCommits_info_219_rfWen ( io_diffCommits_info_219_rfWen ),
    .io_diffCommits_info_219_fpWen ( io_diffCommits_info_219_fpWen ),
    .io_diffCommits_info_219_vecWen ( io_diffCommits_info_219_vecWen ),
    .io_diffCommits_info_219_v0Wen ( io_diffCommits_info_219_v0Wen ),
    .io_diffCommits_info_219_vlWen ( io_diffCommits_info_219_vlWen ),
    .io_diffCommits_info_220_ldest ( io_diffCommits_info_220_ldest ),
    .io_diffCommits_info_220_pdest ( io_diffCommits_info_220_pdest ),
    .io_diffCommits_info_220_rfWen ( io_diffCommits_info_220_rfWen ),
    .io_diffCommits_info_220_fpWen ( io_diffCommits_info_220_fpWen ),
    .io_diffCommits_info_220_vecWen ( io_diffCommits_info_220_vecWen ),
    .io_diffCommits_info_220_v0Wen ( io_diffCommits_info_220_v0Wen ),
    .io_diffCommits_info_220_vlWen ( io_diffCommits_info_220_vlWen ),
    .io_diffCommits_info_221_ldest ( io_diffCommits_info_221_ldest ),
    .io_diffCommits_info_221_pdest ( io_diffCommits_info_221_pdest ),
    .io_diffCommits_info_221_rfWen ( io_diffCommits_info_221_rfWen ),
    .io_diffCommits_info_221_fpWen ( io_diffCommits_info_221_fpWen ),
    .io_diffCommits_info_221_vecWen ( io_diffCommits_info_221_vecWen ),
    .io_diffCommits_info_221_v0Wen ( io_diffCommits_info_221_v0Wen ),
    .io_diffCommits_info_221_vlWen ( io_diffCommits_info_221_vlWen ),
    .io_diffCommits_info_222_ldest ( io_diffCommits_info_222_ldest ),
    .io_diffCommits_info_222_pdest ( io_diffCommits_info_222_pdest ),
    .io_diffCommits_info_222_rfWen ( io_diffCommits_info_222_rfWen ),
    .io_diffCommits_info_222_fpWen ( io_diffCommits_info_222_fpWen ),
    .io_diffCommits_info_222_vecWen ( io_diffCommits_info_222_vecWen ),
    .io_diffCommits_info_222_v0Wen ( io_diffCommits_info_222_v0Wen ),
    .io_diffCommits_info_222_vlWen ( io_diffCommits_info_222_vlWen ),
    .io_diffCommits_info_223_ldest ( io_diffCommits_info_223_ldest ),
    .io_diffCommits_info_223_pdest ( io_diffCommits_info_223_pdest ),
    .io_diffCommits_info_223_rfWen ( io_diffCommits_info_223_rfWen ),
    .io_diffCommits_info_223_fpWen ( io_diffCommits_info_223_fpWen ),
    .io_diffCommits_info_223_vecWen ( io_diffCommits_info_223_vecWen ),
    .io_diffCommits_info_223_v0Wen ( io_diffCommits_info_223_v0Wen ),
    .io_diffCommits_info_223_vlWen ( io_diffCommits_info_223_vlWen ),
    .io_diffCommits_info_224_ldest ( io_diffCommits_info_224_ldest ),
    .io_diffCommits_info_224_pdest ( io_diffCommits_info_224_pdest ),
    .io_diffCommits_info_224_rfWen ( io_diffCommits_info_224_rfWen ),
    .io_diffCommits_info_224_fpWen ( io_diffCommits_info_224_fpWen ),
    .io_diffCommits_info_224_vecWen ( io_diffCommits_info_224_vecWen ),
    .io_diffCommits_info_224_v0Wen ( io_diffCommits_info_224_v0Wen ),
    .io_diffCommits_info_224_vlWen ( io_diffCommits_info_224_vlWen ),
    .io_diffCommits_info_225_ldest ( io_diffCommits_info_225_ldest ),
    .io_diffCommits_info_225_pdest ( io_diffCommits_info_225_pdest ),
    .io_diffCommits_info_225_rfWen ( io_diffCommits_info_225_rfWen ),
    .io_diffCommits_info_225_fpWen ( io_diffCommits_info_225_fpWen ),
    .io_diffCommits_info_225_vecWen ( io_diffCommits_info_225_vecWen ),
    .io_diffCommits_info_225_v0Wen ( io_diffCommits_info_225_v0Wen ),
    .io_diffCommits_info_225_vlWen ( io_diffCommits_info_225_vlWen ),
    .io_diffCommits_info_226_ldest ( io_diffCommits_info_226_ldest ),
    .io_diffCommits_info_226_pdest ( io_diffCommits_info_226_pdest ),
    .io_diffCommits_info_226_rfWen ( io_diffCommits_info_226_rfWen ),
    .io_diffCommits_info_226_fpWen ( io_diffCommits_info_226_fpWen ),
    .io_diffCommits_info_226_vecWen ( io_diffCommits_info_226_vecWen ),
    .io_diffCommits_info_226_v0Wen ( io_diffCommits_info_226_v0Wen ),
    .io_diffCommits_info_226_vlWen ( io_diffCommits_info_226_vlWen ),
    .io_diffCommits_info_227_ldest ( io_diffCommits_info_227_ldest ),
    .io_diffCommits_info_227_pdest ( io_diffCommits_info_227_pdest ),
    .io_diffCommits_info_227_rfWen ( io_diffCommits_info_227_rfWen ),
    .io_diffCommits_info_227_fpWen ( io_diffCommits_info_227_fpWen ),
    .io_diffCommits_info_227_vecWen ( io_diffCommits_info_227_vecWen ),
    .io_diffCommits_info_227_v0Wen ( io_diffCommits_info_227_v0Wen ),
    .io_diffCommits_info_227_vlWen ( io_diffCommits_info_227_vlWen ),
    .io_diffCommits_info_228_ldest ( io_diffCommits_info_228_ldest ),
    .io_diffCommits_info_228_pdest ( io_diffCommits_info_228_pdest ),
    .io_diffCommits_info_228_rfWen ( io_diffCommits_info_228_rfWen ),
    .io_diffCommits_info_228_fpWen ( io_diffCommits_info_228_fpWen ),
    .io_diffCommits_info_228_vecWen ( io_diffCommits_info_228_vecWen ),
    .io_diffCommits_info_228_v0Wen ( io_diffCommits_info_228_v0Wen ),
    .io_diffCommits_info_228_vlWen ( io_diffCommits_info_228_vlWen ),
    .io_diffCommits_info_229_ldest ( io_diffCommits_info_229_ldest ),
    .io_diffCommits_info_229_pdest ( io_diffCommits_info_229_pdest ),
    .io_diffCommits_info_229_rfWen ( io_diffCommits_info_229_rfWen ),
    .io_diffCommits_info_229_fpWen ( io_diffCommits_info_229_fpWen ),
    .io_diffCommits_info_229_vecWen ( io_diffCommits_info_229_vecWen ),
    .io_diffCommits_info_229_v0Wen ( io_diffCommits_info_229_v0Wen ),
    .io_diffCommits_info_229_vlWen ( io_diffCommits_info_229_vlWen ),
    .io_diffCommits_info_230_ldest ( io_diffCommits_info_230_ldest ),
    .io_diffCommits_info_230_pdest ( io_diffCommits_info_230_pdest ),
    .io_diffCommits_info_230_rfWen ( io_diffCommits_info_230_rfWen ),
    .io_diffCommits_info_230_fpWen ( io_diffCommits_info_230_fpWen ),
    .io_diffCommits_info_230_vecWen ( io_diffCommits_info_230_vecWen ),
    .io_diffCommits_info_230_v0Wen ( io_diffCommits_info_230_v0Wen ),
    .io_diffCommits_info_230_vlWen ( io_diffCommits_info_230_vlWen ),
    .io_diffCommits_info_231_ldest ( io_diffCommits_info_231_ldest ),
    .io_diffCommits_info_231_pdest ( io_diffCommits_info_231_pdest ),
    .io_diffCommits_info_231_rfWen ( io_diffCommits_info_231_rfWen ),
    .io_diffCommits_info_231_fpWen ( io_diffCommits_info_231_fpWen ),
    .io_diffCommits_info_231_vecWen ( io_diffCommits_info_231_vecWen ),
    .io_diffCommits_info_231_v0Wen ( io_diffCommits_info_231_v0Wen ),
    .io_diffCommits_info_231_vlWen ( io_diffCommits_info_231_vlWen ),
    .io_diffCommits_info_232_ldest ( io_diffCommits_info_232_ldest ),
    .io_diffCommits_info_232_pdest ( io_diffCommits_info_232_pdest ),
    .io_diffCommits_info_232_rfWen ( io_diffCommits_info_232_rfWen ),
    .io_diffCommits_info_232_fpWen ( io_diffCommits_info_232_fpWen ),
    .io_diffCommits_info_232_vecWen ( io_diffCommits_info_232_vecWen ),
    .io_diffCommits_info_232_v0Wen ( io_diffCommits_info_232_v0Wen ),
    .io_diffCommits_info_232_vlWen ( io_diffCommits_info_232_vlWen ),
    .io_diffCommits_info_233_ldest ( io_diffCommits_info_233_ldest ),
    .io_diffCommits_info_233_pdest ( io_diffCommits_info_233_pdest ),
    .io_diffCommits_info_233_rfWen ( io_diffCommits_info_233_rfWen ),
    .io_diffCommits_info_233_fpWen ( io_diffCommits_info_233_fpWen ),
    .io_diffCommits_info_233_vecWen ( io_diffCommits_info_233_vecWen ),
    .io_diffCommits_info_233_v0Wen ( io_diffCommits_info_233_v0Wen ),
    .io_diffCommits_info_233_vlWen ( io_diffCommits_info_233_vlWen ),
    .io_diffCommits_info_234_ldest ( io_diffCommits_info_234_ldest ),
    .io_diffCommits_info_234_pdest ( io_diffCommits_info_234_pdest ),
    .io_diffCommits_info_234_rfWen ( io_diffCommits_info_234_rfWen ),
    .io_diffCommits_info_234_fpWen ( io_diffCommits_info_234_fpWen ),
    .io_diffCommits_info_234_vecWen ( io_diffCommits_info_234_vecWen ),
    .io_diffCommits_info_234_v0Wen ( io_diffCommits_info_234_v0Wen ),
    .io_diffCommits_info_234_vlWen ( io_diffCommits_info_234_vlWen ),
    .io_diffCommits_info_235_ldest ( io_diffCommits_info_235_ldest ),
    .io_diffCommits_info_235_pdest ( io_diffCommits_info_235_pdest ),
    .io_diffCommits_info_235_rfWen ( io_diffCommits_info_235_rfWen ),
    .io_diffCommits_info_235_fpWen ( io_diffCommits_info_235_fpWen ),
    .io_diffCommits_info_235_vecWen ( io_diffCommits_info_235_vecWen ),
    .io_diffCommits_info_235_v0Wen ( io_diffCommits_info_235_v0Wen ),
    .io_diffCommits_info_235_vlWen ( io_diffCommits_info_235_vlWen ),
    .io_diffCommits_info_236_ldest ( io_diffCommits_info_236_ldest ),
    .io_diffCommits_info_236_pdest ( io_diffCommits_info_236_pdest ),
    .io_diffCommits_info_236_rfWen ( io_diffCommits_info_236_rfWen ),
    .io_diffCommits_info_236_fpWen ( io_diffCommits_info_236_fpWen ),
    .io_diffCommits_info_236_vecWen ( io_diffCommits_info_236_vecWen ),
    .io_diffCommits_info_236_v0Wen ( io_diffCommits_info_236_v0Wen ),
    .io_diffCommits_info_236_vlWen ( io_diffCommits_info_236_vlWen ),
    .io_diffCommits_info_237_ldest ( io_diffCommits_info_237_ldest ),
    .io_diffCommits_info_237_pdest ( io_diffCommits_info_237_pdest ),
    .io_diffCommits_info_237_rfWen ( io_diffCommits_info_237_rfWen ),
    .io_diffCommits_info_237_fpWen ( io_diffCommits_info_237_fpWen ),
    .io_diffCommits_info_237_vecWen ( io_diffCommits_info_237_vecWen ),
    .io_diffCommits_info_237_v0Wen ( io_diffCommits_info_237_v0Wen ),
    .io_diffCommits_info_237_vlWen ( io_diffCommits_info_237_vlWen ),
    .io_diffCommits_info_238_ldest ( io_diffCommits_info_238_ldest ),
    .io_diffCommits_info_238_pdest ( io_diffCommits_info_238_pdest ),
    .io_diffCommits_info_238_rfWen ( io_diffCommits_info_238_rfWen ),
    .io_diffCommits_info_238_fpWen ( io_diffCommits_info_238_fpWen ),
    .io_diffCommits_info_238_vecWen ( io_diffCommits_info_238_vecWen ),
    .io_diffCommits_info_238_v0Wen ( io_diffCommits_info_238_v0Wen ),
    .io_diffCommits_info_238_vlWen ( io_diffCommits_info_238_vlWen ),
    .io_diffCommits_info_239_ldest ( io_diffCommits_info_239_ldest ),
    .io_diffCommits_info_239_pdest ( io_diffCommits_info_239_pdest ),
    .io_diffCommits_info_239_rfWen ( io_diffCommits_info_239_rfWen ),
    .io_diffCommits_info_239_fpWen ( io_diffCommits_info_239_fpWen ),
    .io_diffCommits_info_239_vecWen ( io_diffCommits_info_239_vecWen ),
    .io_diffCommits_info_239_v0Wen ( io_diffCommits_info_239_v0Wen ),
    .io_diffCommits_info_239_vlWen ( io_diffCommits_info_239_vlWen ),
    .io_diffCommits_info_240_ldest ( io_diffCommits_info_240_ldest ),
    .io_diffCommits_info_240_pdest ( io_diffCommits_info_240_pdest ),
    .io_diffCommits_info_240_rfWen ( io_diffCommits_info_240_rfWen ),
    .io_diffCommits_info_240_fpWen ( io_diffCommits_info_240_fpWen ),
    .io_diffCommits_info_240_vecWen ( io_diffCommits_info_240_vecWen ),
    .io_diffCommits_info_240_v0Wen ( io_diffCommits_info_240_v0Wen ),
    .io_diffCommits_info_240_vlWen ( io_diffCommits_info_240_vlWen ),
    .io_diffCommits_info_241_ldest ( io_diffCommits_info_241_ldest ),
    .io_diffCommits_info_241_pdest ( io_diffCommits_info_241_pdest ),
    .io_diffCommits_info_241_rfWen ( io_diffCommits_info_241_rfWen ),
    .io_diffCommits_info_241_fpWen ( io_diffCommits_info_241_fpWen ),
    .io_diffCommits_info_241_vecWen ( io_diffCommits_info_241_vecWen ),
    .io_diffCommits_info_241_v0Wen ( io_diffCommits_info_241_v0Wen ),
    .io_diffCommits_info_241_vlWen ( io_diffCommits_info_241_vlWen ),
    .io_diffCommits_info_242_ldest ( io_diffCommits_info_242_ldest ),
    .io_diffCommits_info_242_pdest ( io_diffCommits_info_242_pdest ),
    .io_diffCommits_info_242_rfWen ( io_diffCommits_info_242_rfWen ),
    .io_diffCommits_info_242_fpWen ( io_diffCommits_info_242_fpWen ),
    .io_diffCommits_info_242_vecWen ( io_diffCommits_info_242_vecWen ),
    .io_diffCommits_info_242_v0Wen ( io_diffCommits_info_242_v0Wen ),
    .io_diffCommits_info_242_vlWen ( io_diffCommits_info_242_vlWen ),
    .io_diffCommits_info_243_ldest ( io_diffCommits_info_243_ldest ),
    .io_diffCommits_info_243_pdest ( io_diffCommits_info_243_pdest ),
    .io_diffCommits_info_243_rfWen ( io_diffCommits_info_243_rfWen ),
    .io_diffCommits_info_243_fpWen ( io_diffCommits_info_243_fpWen ),
    .io_diffCommits_info_243_vecWen ( io_diffCommits_info_243_vecWen ),
    .io_diffCommits_info_243_v0Wen ( io_diffCommits_info_243_v0Wen ),
    .io_diffCommits_info_243_vlWen ( io_diffCommits_info_243_vlWen ),
    .io_diffCommits_info_244_ldest ( io_diffCommits_info_244_ldest ),
    .io_diffCommits_info_244_pdest ( io_diffCommits_info_244_pdest ),
    .io_diffCommits_info_244_rfWen ( io_diffCommits_info_244_rfWen ),
    .io_diffCommits_info_244_fpWen ( io_diffCommits_info_244_fpWen ),
    .io_diffCommits_info_244_vecWen ( io_diffCommits_info_244_vecWen ),
    .io_diffCommits_info_244_v0Wen ( io_diffCommits_info_244_v0Wen ),
    .io_diffCommits_info_244_vlWen ( io_diffCommits_info_244_vlWen ),
    .io_diffCommits_info_245_ldest ( io_diffCommits_info_245_ldest ),
    .io_diffCommits_info_245_pdest ( io_diffCommits_info_245_pdest ),
    .io_diffCommits_info_245_rfWen ( io_diffCommits_info_245_rfWen ),
    .io_diffCommits_info_245_fpWen ( io_diffCommits_info_245_fpWen ),
    .io_diffCommits_info_245_vecWen ( io_diffCommits_info_245_vecWen ),
    .io_diffCommits_info_245_v0Wen ( io_diffCommits_info_245_v0Wen ),
    .io_diffCommits_info_245_vlWen ( io_diffCommits_info_245_vlWen ),
    .io_diffCommits_info_246_ldest ( io_diffCommits_info_246_ldest ),
    .io_diffCommits_info_246_pdest ( io_diffCommits_info_246_pdest ),
    .io_diffCommits_info_246_rfWen ( io_diffCommits_info_246_rfWen ),
    .io_diffCommits_info_246_fpWen ( io_diffCommits_info_246_fpWen ),
    .io_diffCommits_info_246_vecWen ( io_diffCommits_info_246_vecWen ),
    .io_diffCommits_info_246_v0Wen ( io_diffCommits_info_246_v0Wen ),
    .io_diffCommits_info_246_vlWen ( io_diffCommits_info_246_vlWen ),
    .io_diffCommits_info_247_ldest ( io_diffCommits_info_247_ldest ),
    .io_diffCommits_info_247_pdest ( io_diffCommits_info_247_pdest ),
    .io_diffCommits_info_247_rfWen ( io_diffCommits_info_247_rfWen ),
    .io_diffCommits_info_247_fpWen ( io_diffCommits_info_247_fpWen ),
    .io_diffCommits_info_247_vecWen ( io_diffCommits_info_247_vecWen ),
    .io_diffCommits_info_247_v0Wen ( io_diffCommits_info_247_v0Wen ),
    .io_diffCommits_info_247_vlWen ( io_diffCommits_info_247_vlWen ),
    .io_diffCommits_info_248_ldest ( io_diffCommits_info_248_ldest ),
    .io_diffCommits_info_248_pdest ( io_diffCommits_info_248_pdest ),
    .io_diffCommits_info_248_rfWen ( io_diffCommits_info_248_rfWen ),
    .io_diffCommits_info_248_fpWen ( io_diffCommits_info_248_fpWen ),
    .io_diffCommits_info_248_vecWen ( io_diffCommits_info_248_vecWen ),
    .io_diffCommits_info_248_v0Wen ( io_diffCommits_info_248_v0Wen ),
    .io_diffCommits_info_248_vlWen ( io_diffCommits_info_248_vlWen ),
    .io_diffCommits_info_249_ldest ( io_diffCommits_info_249_ldest ),
    .io_diffCommits_info_249_pdest ( io_diffCommits_info_249_pdest ),
    .io_diffCommits_info_249_rfWen ( io_diffCommits_info_249_rfWen ),
    .io_diffCommits_info_249_fpWen ( io_diffCommits_info_249_fpWen ),
    .io_diffCommits_info_249_vecWen ( io_diffCommits_info_249_vecWen ),
    .io_diffCommits_info_249_v0Wen ( io_diffCommits_info_249_v0Wen ),
    .io_diffCommits_info_249_vlWen ( io_diffCommits_info_249_vlWen ),
    .io_diffCommits_info_250_ldest ( io_diffCommits_info_250_ldest ),
    .io_diffCommits_info_250_pdest ( io_diffCommits_info_250_pdest ),
    .io_diffCommits_info_250_rfWen ( io_diffCommits_info_250_rfWen ),
    .io_diffCommits_info_250_fpWen ( io_diffCommits_info_250_fpWen ),
    .io_diffCommits_info_250_vecWen ( io_diffCommits_info_250_vecWen ),
    .io_diffCommits_info_250_v0Wen ( io_diffCommits_info_250_v0Wen ),
    .io_diffCommits_info_250_vlWen ( io_diffCommits_info_250_vlWen ),
    .io_diffCommits_info_251_ldest ( io_diffCommits_info_251_ldest ),
    .io_diffCommits_info_251_pdest ( io_diffCommits_info_251_pdest ),
    .io_diffCommits_info_251_rfWen ( io_diffCommits_info_251_rfWen ),
    .io_diffCommits_info_251_fpWen ( io_diffCommits_info_251_fpWen ),
    .io_diffCommits_info_251_vecWen ( io_diffCommits_info_251_vecWen ),
    .io_diffCommits_info_251_v0Wen ( io_diffCommits_info_251_v0Wen ),
    .io_diffCommits_info_251_vlWen ( io_diffCommits_info_251_vlWen ),
    .io_diffCommits_info_252_ldest ( io_diffCommits_info_252_ldest ),
    .io_diffCommits_info_252_pdest ( io_diffCommits_info_252_pdest ),
    .io_diffCommits_info_252_rfWen ( io_diffCommits_info_252_rfWen ),
    .io_diffCommits_info_252_fpWen ( io_diffCommits_info_252_fpWen ),
    .io_diffCommits_info_252_vecWen ( io_diffCommits_info_252_vecWen ),
    .io_diffCommits_info_252_v0Wen ( io_diffCommits_info_252_v0Wen ),
    .io_diffCommits_info_252_vlWen ( io_diffCommits_info_252_vlWen ),
    .io_diffCommits_info_253_ldest ( io_diffCommits_info_253_ldest ),
    .io_diffCommits_info_253_pdest ( io_diffCommits_info_253_pdest ),
    .io_diffCommits_info_253_rfWen ( io_diffCommits_info_253_rfWen ),
    .io_diffCommits_info_253_fpWen ( io_diffCommits_info_253_fpWen ),
    .io_diffCommits_info_253_vecWen ( io_diffCommits_info_253_vecWen ),
    .io_diffCommits_info_253_v0Wen ( io_diffCommits_info_253_v0Wen ),
    .io_diffCommits_info_253_vlWen ( io_diffCommits_info_253_vlWen ),
    .io_diffCommits_info_254_ldest ( io_diffCommits_info_254_ldest ),
    .io_diffCommits_info_254_pdest ( io_diffCommits_info_254_pdest ),
    .io_diffCommits_info_254_rfWen ( io_diffCommits_info_254_rfWen ),
    .io_diffCommits_info_254_fpWen ( io_diffCommits_info_254_fpWen ),
    .io_diffCommits_info_254_vecWen ( io_diffCommits_info_254_vecWen ),
    .io_diffCommits_info_254_v0Wen ( io_diffCommits_info_254_v0Wen ),
    .io_diffCommits_info_254_vlWen ( io_diffCommits_info_254_vlWen ),
    .io_diffCommits_info_255_ldest ( io_diffCommits_info_255_ldest ),
    .io_diffCommits_info_255_pdest ( io_diffCommits_info_255_pdest ),
    .io_diffCommits_info_256_ldest ( io_diffCommits_info_256_ldest ),
    .io_diffCommits_info_256_pdest ( io_diffCommits_info_256_pdest ),
    .io_diffCommits_info_257_ldest ( io_diffCommits_info_257_ldest ),
    .io_diffCommits_info_257_pdest ( io_diffCommits_info_257_pdest ),
    .io_diffCommits_info_258_ldest ( io_diffCommits_info_258_ldest ),
    .io_diffCommits_info_258_pdest ( io_diffCommits_info_258_pdest ),
    .io_diffCommits_info_259_ldest ( io_diffCommits_info_259_ldest ),
    .io_diffCommits_info_259_pdest ( io_diffCommits_info_259_pdest ),
    .io_diffCommits_info_260_ldest ( io_diffCommits_info_260_ldest ),
    .io_diffCommits_info_260_pdest ( io_diffCommits_info_260_pdest ),
    .io_diffCommits_info_261_ldest ( io_diffCommits_info_261_ldest ),
    .io_diffCommits_info_261_pdest ( io_diffCommits_info_261_pdest ),
    .io_diffCommits_info_262_ldest ( io_diffCommits_info_262_ldest ),
    .io_diffCommits_info_262_pdest ( io_diffCommits_info_262_pdest ),
    .io_diffCommits_info_263_ldest ( io_diffCommits_info_263_ldest ),
    .io_diffCommits_info_263_pdest ( io_diffCommits_info_263_pdest ),
    .io_diffCommits_info_264_ldest ( io_diffCommits_info_264_ldest ),
    .io_diffCommits_info_264_pdest ( io_diffCommits_info_264_pdest ),
    .io_diffCommits_info_265_ldest ( io_diffCommits_info_265_ldest ),
    .io_diffCommits_info_265_pdest ( io_diffCommits_info_265_pdest ),
    .io_diffCommits_info_266_ldest ( io_diffCommits_info_266_ldest ),
    .io_diffCommits_info_266_pdest ( io_diffCommits_info_266_pdest ),
    .io_diffCommits_info_267_ldest ( io_diffCommits_info_267_ldest ),
    .io_diffCommits_info_267_pdest ( io_diffCommits_info_267_pdest ),
    .io_diffCommits_info_268_ldest ( io_diffCommits_info_268_ldest ),
    .io_diffCommits_info_268_pdest ( io_diffCommits_info_268_pdest ),
    .io_diffCommits_info_269_ldest ( io_diffCommits_info_269_ldest ),
    .io_diffCommits_info_269_pdest ( io_diffCommits_info_269_pdest ),
    .io_diffCommits_info_270_ldest ( io_diffCommits_info_270_ldest ),
    .io_diffCommits_info_270_pdest ( io_diffCommits_info_270_pdest ),
    .io_diffCommits_info_271_ldest ( io_diffCommits_info_271_ldest ),
    .io_diffCommits_info_271_pdest ( io_diffCommits_info_271_pdest ),
    .io_diffCommits_info_272_ldest ( io_diffCommits_info_272_ldest ),
    .io_diffCommits_info_272_pdest ( io_diffCommits_info_272_pdest ),
    .io_diffCommits_info_273_ldest ( io_diffCommits_info_273_ldest ),
    .io_diffCommits_info_273_pdest ( io_diffCommits_info_273_pdest ),
    .io_diffCommits_info_274_ldest ( io_diffCommits_info_274_ldest ),
    .io_diffCommits_info_274_pdest ( io_diffCommits_info_274_pdest ),
    .io_diffCommits_info_275_ldest ( io_diffCommits_info_275_ldest ),
    .io_diffCommits_info_275_pdest ( io_diffCommits_info_275_pdest ),
    .io_diffCommits_info_276_ldest ( io_diffCommits_info_276_ldest ),
    .io_diffCommits_info_276_pdest ( io_diffCommits_info_276_pdest ),
    .io_diffCommits_info_277_ldest ( io_diffCommits_info_277_ldest ),
    .io_diffCommits_info_277_pdest ( io_diffCommits_info_277_pdest ),
    .io_diffCommits_info_278_ldest ( io_diffCommits_info_278_ldest ),
    .io_diffCommits_info_278_pdest ( io_diffCommits_info_278_pdest ),
    .io_diffCommits_info_279_ldest ( io_diffCommits_info_279_ldest ),
    .io_diffCommits_info_279_pdest ( io_diffCommits_info_279_pdest ),
    .io_diffCommits_info_280_ldest ( io_diffCommits_info_280_ldest ),
    .io_diffCommits_info_280_pdest ( io_diffCommits_info_280_pdest ),
    .io_diffCommits_info_281_ldest ( io_diffCommits_info_281_ldest ),
    .io_diffCommits_info_281_pdest ( io_diffCommits_info_281_pdest ),
    .io_diffCommits_info_282_ldest ( io_diffCommits_info_282_ldest ),
    .io_diffCommits_info_282_pdest ( io_diffCommits_info_282_pdest ),
    .io_diffCommits_info_283_ldest ( io_diffCommits_info_283_ldest ),
    .io_diffCommits_info_283_pdest ( io_diffCommits_info_283_pdest ),
    .io_diffCommits_info_284_ldest ( io_diffCommits_info_284_ldest ),
    .io_diffCommits_info_284_pdest ( io_diffCommits_info_284_pdest ),
    .io_diffCommits_info_285_ldest ( io_diffCommits_info_285_ldest ),
    .io_diffCommits_info_285_pdest ( io_diffCommits_info_285_pdest ),
    .io_diffCommits_info_286_ldest ( io_diffCommits_info_286_ldest ),
    .io_diffCommits_info_286_pdest ( io_diffCommits_info_286_pdest ),
    .io_diffCommits_info_287_ldest ( io_diffCommits_info_287_ldest ),
    .io_diffCommits_info_287_pdest ( io_diffCommits_info_287_pdest ),
    .io_diffCommits_info_288_ldest ( io_diffCommits_info_288_ldest ),
    .io_diffCommits_info_288_pdest ( io_diffCommits_info_288_pdest ),
    .io_diffCommits_info_289_ldest ( io_diffCommits_info_289_ldest ),
    .io_diffCommits_info_289_pdest ( io_diffCommits_info_289_pdest ),
    .io_diffCommits_info_290_ldest ( io_diffCommits_info_290_ldest ),
    .io_diffCommits_info_290_pdest ( io_diffCommits_info_290_pdest ),
    .io_diffCommits_info_291_ldest ( io_diffCommits_info_291_ldest ),
    .io_diffCommits_info_291_pdest ( io_diffCommits_info_291_pdest ),
    .io_diffCommits_info_292_ldest ( io_diffCommits_info_292_ldest ),
    .io_diffCommits_info_292_pdest ( io_diffCommits_info_292_pdest ),
    .io_diffCommits_info_293_ldest ( io_diffCommits_info_293_ldest ),
    .io_diffCommits_info_293_pdest ( io_diffCommits_info_293_pdest ),
    .io_diffCommits_info_294_ldest ( io_diffCommits_info_294_ldest ),
    .io_diffCommits_info_294_pdest ( io_diffCommits_info_294_pdest ),
    .io_diffCommits_info_295_ldest ( io_diffCommits_info_295_ldest ),
    .io_diffCommits_info_295_pdest ( io_diffCommits_info_295_pdest ),
    .io_diffCommits_info_296_ldest ( io_diffCommits_info_296_ldest ),
    .io_diffCommits_info_296_pdest ( io_diffCommits_info_296_pdest ),
    .io_diffCommits_info_297_ldest ( io_diffCommits_info_297_ldest ),
    .io_diffCommits_info_297_pdest ( io_diffCommits_info_297_pdest ),
    .io_diffCommits_info_298_ldest ( io_diffCommits_info_298_ldest ),
    .io_diffCommits_info_298_pdest ( io_diffCommits_info_298_pdest ),
    .io_diffCommits_info_299_ldest ( io_diffCommits_info_299_ldest ),
    .io_diffCommits_info_299_pdest ( io_diffCommits_info_299_pdest ),
    .io_diffCommits_info_300_ldest ( io_diffCommits_info_300_ldest ),
    .io_diffCommits_info_300_pdest ( io_diffCommits_info_300_pdest ),
    .io_diffCommits_info_301_ldest ( io_diffCommits_info_301_ldest ),
    .io_diffCommits_info_301_pdest ( io_diffCommits_info_301_pdest ),
    .io_diffCommits_info_302_ldest ( io_diffCommits_info_302_ldest ),
    .io_diffCommits_info_302_pdest ( io_diffCommits_info_302_pdest ),
    .io_diffCommits_info_303_ldest ( io_diffCommits_info_303_ldest ),
    .io_diffCommits_info_303_pdest ( io_diffCommits_info_303_pdest ),
    .io_diffCommits_info_304_ldest ( io_diffCommits_info_304_ldest ),
    .io_diffCommits_info_304_pdest ( io_diffCommits_info_304_pdest ),
    .io_diffCommits_info_305_ldest ( io_diffCommits_info_305_ldest ),
    .io_diffCommits_info_305_pdest ( io_diffCommits_info_305_pdest ),
    .io_diffCommits_info_306_ldest ( io_diffCommits_info_306_ldest ),
    .io_diffCommits_info_306_pdest ( io_diffCommits_info_306_pdest ),
    .io_diffCommits_info_307_ldest ( io_diffCommits_info_307_ldest ),
    .io_diffCommits_info_307_pdest ( io_diffCommits_info_307_pdest ),
    .io_diffCommits_info_308_ldest ( io_diffCommits_info_308_ldest ),
    .io_diffCommits_info_308_pdest ( io_diffCommits_info_308_pdest ),
    .io_diffCommits_info_309_ldest ( io_diffCommits_info_309_ldest ),
    .io_diffCommits_info_309_pdest ( io_diffCommits_info_309_pdest ),
    .io_diffCommits_info_310_ldest ( io_diffCommits_info_310_ldest ),
    .io_diffCommits_info_310_pdest ( io_diffCommits_info_310_pdest ),
    .io_diffCommits_info_311_ldest ( io_diffCommits_info_311_ldest ),
    .io_diffCommits_info_311_pdest ( io_diffCommits_info_311_pdest ),
    .io_diffCommits_info_312_ldest ( io_diffCommits_info_312_ldest ),
    .io_diffCommits_info_312_pdest ( io_diffCommits_info_312_pdest ),
    .io_diffCommits_info_313_ldest ( io_diffCommits_info_313_ldest ),
    .io_diffCommits_info_313_pdest ( io_diffCommits_info_313_pdest ),
    .io_diffCommits_info_314_ldest ( io_diffCommits_info_314_ldest ),
    .io_diffCommits_info_314_pdest ( io_diffCommits_info_314_pdest ),
    .io_diffCommits_info_315_ldest ( io_diffCommits_info_315_ldest ),
    .io_diffCommits_info_315_pdest ( io_diffCommits_info_315_pdest ),
    .io_diffCommits_info_316_ldest ( io_diffCommits_info_316_ldest ),
    .io_diffCommits_info_316_pdest ( io_diffCommits_info_316_pdest ),
    .io_diffCommits_info_317_ldest ( io_diffCommits_info_317_ldest ),
    .io_diffCommits_info_317_pdest ( io_diffCommits_info_317_pdest ),
    .io_diffCommits_info_318_ldest ( io_diffCommits_info_318_ldest ),
    .io_diffCommits_info_318_pdest ( io_diffCommits_info_318_pdest ),
    .io_diffCommits_info_319_ldest ( io_diffCommits_info_319_ldest ),
    .io_diffCommits_info_319_pdest ( io_diffCommits_info_319_pdest ),
    .io_diffCommits_info_320_ldest ( io_diffCommits_info_320_ldest ),
    .io_diffCommits_info_320_pdest ( io_diffCommits_info_320_pdest ),
    .io_diffCommits_info_321_ldest ( io_diffCommits_info_321_ldest ),
    .io_diffCommits_info_321_pdest ( io_diffCommits_info_321_pdest ),
    .io_diffCommits_info_322_ldest ( io_diffCommits_info_322_ldest ),
    .io_diffCommits_info_322_pdest ( io_diffCommits_info_322_pdest ),
    .io_diffCommits_info_323_ldest ( io_diffCommits_info_323_ldest ),
    .io_diffCommits_info_323_pdest ( io_diffCommits_info_323_pdest ),
    .io_diffCommits_info_324_ldest ( io_diffCommits_info_324_ldest ),
    .io_diffCommits_info_324_pdest ( io_diffCommits_info_324_pdest ),
    .io_diffCommits_info_325_ldest ( io_diffCommits_info_325_ldest ),
    .io_diffCommits_info_325_pdest ( io_diffCommits_info_325_pdest ),
    .io_diffCommits_info_326_ldest ( io_diffCommits_info_326_ldest ),
    .io_diffCommits_info_326_pdest ( io_diffCommits_info_326_pdest ),
    .io_diffCommits_info_327_ldest ( io_diffCommits_info_327_ldest ),
    .io_diffCommits_info_327_pdest ( io_diffCommits_info_327_pdest ),
    .io_diffCommits_info_328_ldest ( io_diffCommits_info_328_ldest ),
    .io_diffCommits_info_328_pdest ( io_diffCommits_info_328_pdest ),
    .io_diffCommits_info_329_ldest ( io_diffCommits_info_329_ldest ),
    .io_diffCommits_info_329_pdest ( io_diffCommits_info_329_pdest ),
    .io_diffCommits_info_330_ldest ( io_diffCommits_info_330_ldest ),
    .io_diffCommits_info_330_pdest ( io_diffCommits_info_330_pdest ),
    .io_diffCommits_info_331_ldest ( io_diffCommits_info_331_ldest ),
    .io_diffCommits_info_331_pdest ( io_diffCommits_info_331_pdest ),
    .io_diffCommits_info_332_ldest ( io_diffCommits_info_332_ldest ),
    .io_diffCommits_info_332_pdest ( io_diffCommits_info_332_pdest ),
    .io_diffCommits_info_333_ldest ( io_diffCommits_info_333_ldest ),
    .io_diffCommits_info_333_pdest ( io_diffCommits_info_333_pdest ),
    .io_diffCommits_info_334_ldest ( io_diffCommits_info_334_ldest ),
    .io_diffCommits_info_334_pdest ( io_diffCommits_info_334_pdest ),
    .io_diffCommits_info_335_ldest ( io_diffCommits_info_335_ldest ),
    .io_diffCommits_info_335_pdest ( io_diffCommits_info_335_pdest ),
    .io_diffCommits_info_336_ldest ( io_diffCommits_info_336_ldest ),
    .io_diffCommits_info_336_pdest ( io_diffCommits_info_336_pdest ),
    .io_diffCommits_info_337_ldest ( io_diffCommits_info_337_ldest ),
    .io_diffCommits_info_337_pdest ( io_diffCommits_info_337_pdest ),
    .io_diffCommits_info_338_ldest ( io_diffCommits_info_338_ldest ),
    .io_diffCommits_info_338_pdest ( io_diffCommits_info_338_pdest ),
    .io_diffCommits_info_339_ldest ( io_diffCommits_info_339_ldest ),
    .io_diffCommits_info_339_pdest ( io_diffCommits_info_339_pdest ),
    .io_diffCommits_info_340_ldest ( io_diffCommits_info_340_ldest ),
    .io_diffCommits_info_340_pdest ( io_diffCommits_info_340_pdest ),
    .io_diffCommits_info_341_ldest ( io_diffCommits_info_341_ldest ),
    .io_diffCommits_info_341_pdest ( io_diffCommits_info_341_pdest ),
    .io_diffCommits_info_342_ldest ( io_diffCommits_info_342_ldest ),
    .io_diffCommits_info_342_pdest ( io_diffCommits_info_342_pdest ),
    .io_diffCommits_info_343_ldest ( io_diffCommits_info_343_ldest ),
    .io_diffCommits_info_343_pdest ( io_diffCommits_info_343_pdest ),
    .io_diffCommits_info_344_ldest ( io_diffCommits_info_344_ldest ),
    .io_diffCommits_info_344_pdest ( io_diffCommits_info_344_pdest ),
    .io_diffCommits_info_345_ldest ( io_diffCommits_info_345_ldest ),
    .io_diffCommits_info_345_pdest ( io_diffCommits_info_345_pdest ),
    .io_diffCommits_info_346_ldest ( io_diffCommits_info_346_ldest ),
    .io_diffCommits_info_346_pdest ( io_diffCommits_info_346_pdest ),
    .io_diffCommits_info_347_ldest ( io_diffCommits_info_347_ldest ),
    .io_diffCommits_info_347_pdest ( io_diffCommits_info_347_pdest ),
    .io_diffCommits_info_348_ldest ( io_diffCommits_info_348_ldest ),
    .io_diffCommits_info_348_pdest ( io_diffCommits_info_348_pdest ),
    .io_diffCommits_info_349_ldest ( io_diffCommits_info_349_ldest ),
    .io_diffCommits_info_349_pdest ( io_diffCommits_info_349_pdest ),
    .io_diffCommits_info_350_ldest ( io_diffCommits_info_350_ldest ),
    .io_diffCommits_info_350_pdest ( io_diffCommits_info_350_pdest ),
    .io_diffCommits_info_351_ldest ( io_diffCommits_info_351_ldest ),
    .io_diffCommits_info_351_pdest ( io_diffCommits_info_351_pdest ),
    .io_diffCommits_info_352_ldest ( io_diffCommits_info_352_ldest ),
    .io_diffCommits_info_352_pdest ( io_diffCommits_info_352_pdest ),
    .io_diffCommits_info_353_ldest ( io_diffCommits_info_353_ldest ),
    .io_diffCommits_info_353_pdest ( io_diffCommits_info_353_pdest ),
    .io_diffCommits_info_354_ldest ( io_diffCommits_info_354_ldest ),
    .io_diffCommits_info_354_pdest ( io_diffCommits_info_354_pdest ),
    .io_diffCommits_info_355_ldest ( io_diffCommits_info_355_ldest ),
    .io_diffCommits_info_355_pdest ( io_diffCommits_info_355_pdest ),
    .io_diffCommits_info_356_ldest ( io_diffCommits_info_356_ldest ),
    .io_diffCommits_info_356_pdest ( io_diffCommits_info_356_pdest ),
    .io_diffCommits_info_357_ldest ( io_diffCommits_info_357_ldest ),
    .io_diffCommits_info_357_pdest ( io_diffCommits_info_357_pdest ),
    .io_diffCommits_info_358_ldest ( io_diffCommits_info_358_ldest ),
    .io_diffCommits_info_358_pdest ( io_diffCommits_info_358_pdest ),
    .io_diffCommits_info_359_ldest ( io_diffCommits_info_359_ldest ),
    .io_diffCommits_info_359_pdest ( io_diffCommits_info_359_pdest ),
    .io_diffCommits_info_360_ldest ( io_diffCommits_info_360_ldest ),
    .io_diffCommits_info_360_pdest ( io_diffCommits_info_360_pdest ),
    .io_diffCommits_info_361_ldest ( io_diffCommits_info_361_ldest ),
    .io_diffCommits_info_361_pdest ( io_diffCommits_info_361_pdest ),
    .io_diffCommits_info_362_ldest ( io_diffCommits_info_362_ldest ),
    .io_diffCommits_info_362_pdest ( io_diffCommits_info_362_pdest ),
    .io_diffCommits_info_363_ldest ( io_diffCommits_info_363_ldest ),
    .io_diffCommits_info_363_pdest ( io_diffCommits_info_363_pdest ),
    .io_diffCommits_info_364_ldest ( io_diffCommits_info_364_ldest ),
    .io_diffCommits_info_364_pdest ( io_diffCommits_info_364_pdest ),
    .io_diffCommits_info_365_ldest ( io_diffCommits_info_365_ldest ),
    .io_diffCommits_info_365_pdest ( io_diffCommits_info_365_pdest ),
    .io_diffCommits_info_366_ldest ( io_diffCommits_info_366_ldest ),
    .io_diffCommits_info_366_pdest ( io_diffCommits_info_366_pdest ),
    .io_diffCommits_info_367_ldest ( io_diffCommits_info_367_ldest ),
    .io_diffCommits_info_367_pdest ( io_diffCommits_info_367_pdest ),
    .io_diffCommits_info_368_ldest ( io_diffCommits_info_368_ldest ),
    .io_diffCommits_info_368_pdest ( io_diffCommits_info_368_pdest ),
    .io_diffCommits_info_369_ldest ( io_diffCommits_info_369_ldest ),
    .io_diffCommits_info_369_pdest ( io_diffCommits_info_369_pdest ),
    .io_diffCommits_info_370_ldest ( io_diffCommits_info_370_ldest ),
    .io_diffCommits_info_370_pdest ( io_diffCommits_info_370_pdest ),
    .io_diffCommits_info_371_ldest ( io_diffCommits_info_371_ldest ),
    .io_diffCommits_info_371_pdest ( io_diffCommits_info_371_pdest ),
    .io_diffCommits_info_372_ldest ( io_diffCommits_info_372_ldest ),
    .io_diffCommits_info_372_pdest ( io_diffCommits_info_372_pdest ),
    .io_diffCommits_info_373_ldest ( io_diffCommits_info_373_ldest ),
    .io_diffCommits_info_373_pdest ( io_diffCommits_info_373_pdest ),
    .io_diffCommits_info_374_ldest ( io_diffCommits_info_374_ldest ),
    .io_diffCommits_info_374_pdest ( io_diffCommits_info_374_pdest ),
    .io_diffCommits_info_375_ldest ( io_diffCommits_info_375_ldest ),
    .io_diffCommits_info_375_pdest ( io_diffCommits_info_375_pdest ),
    .io_diffCommits_info_376_ldest ( io_diffCommits_info_376_ldest ),
    .io_diffCommits_info_376_pdest ( io_diffCommits_info_376_pdest ),
    .io_diffCommits_info_377_ldest ( io_diffCommits_info_377_ldest ),
    .io_diffCommits_info_377_pdest ( io_diffCommits_info_377_pdest ),
    .io_diffCommits_info_378_ldest ( io_diffCommits_info_378_ldest ),
    .io_diffCommits_info_378_pdest ( io_diffCommits_info_378_pdest ),
    .io_diffCommits_info_379_ldest ( io_diffCommits_info_379_ldest ),
    .io_diffCommits_info_379_pdest ( io_diffCommits_info_379_pdest ),
    .io_diffCommits_info_380_ldest ( io_diffCommits_info_380_ldest ),
    .io_diffCommits_info_380_pdest ( io_diffCommits_info_380_pdest ),
    .io_diffCommits_info_381_ldest ( io_diffCommits_info_381_ldest ),
    .io_diffCommits_info_381_pdest ( io_diffCommits_info_381_pdest ),
    .io_diffCommits_info_382_ldest ( io_diffCommits_info_382_ldest ),
    .io_diffCommits_info_382_pdest ( io_diffCommits_info_382_pdest ),
    .io_diffCommits_info_383_ldest ( io_diffCommits_info_383_ldest ),
    .io_diffCommits_info_383_pdest ( io_diffCommits_info_383_pdest ),
    .io_diffCommits_info_384_ldest ( io_diffCommits_info_384_ldest ),
    .io_diffCommits_info_384_pdest ( io_diffCommits_info_384_pdest ),
    .io_diffCommits_info_385_ldest ( io_diffCommits_info_385_ldest ),
    .io_diffCommits_info_385_pdest ( io_diffCommits_info_385_pdest ),
    .io_diffCommits_info_386_ldest ( io_diffCommits_info_386_ldest ),
    .io_diffCommits_info_386_pdest ( io_diffCommits_info_386_pdest ),
    .io_diffCommits_info_387_ldest ( io_diffCommits_info_387_ldest ),
    .io_diffCommits_info_387_pdest ( io_diffCommits_info_387_pdest ),
    .io_diffCommits_info_388_ldest ( io_diffCommits_info_388_ldest ),
    .io_diffCommits_info_388_pdest ( io_diffCommits_info_388_pdest ),
    .io_diffCommits_info_389_ldest ( io_diffCommits_info_389_ldest ),
    .io_diffCommits_info_389_pdest ( io_diffCommits_info_389_pdest ),
    .io_lsq_scommit       ( io_lsq_scommit       ),
    .io_lsq_pendingMMIOld ( io_lsq_pendingMMIOld ),
    .io_lsq_pendingst     ( io_lsq_pendingst     ),
    .io_lsq_pendingPtr_flag ( io_lsq_pendingPtr_flag ),
    .io_lsq_pendingPtr_value ( io_lsq_pendingPtr_value ),
    .io_robDeqPtr_flag    ( io_robDeqPtr_flag    ),
    .io_robDeqPtr_value   ( io_robDeqPtr_value   ),
    .io_csr_fflags_valid  ( io_csr_fflags_valid  ),
    .io_csr_fflags_bits   ( io_csr_fflags_bits   ),
    .io_csr_vxsat_valid   ( io_csr_vxsat_valid   ),
    .io_csr_vxsat_bits    ( io_csr_vxsat_bits    ),
    .io_csr_vstart_valid  ( io_csr_vstart_valid  ),
    .io_csr_vstart_bits   ( io_csr_vstart_bits   ),
    .io_csr_dirty_fs      ( io_csr_dirty_fs      ),
    .io_csr_dirty_vs      ( io_csr_dirty_vs      ),
    .io_csr_perfinfo_retiredInstr ( io_csr_perfinfo_retiredInstr ),
    .io_cpu_halt          ( io_cpu_halt          ),
    .io_wfi_wfiReq        ( io_wfi_wfiReq        ),
    .io_toDecode_isResumeVType ( io_toDecode_isResumeVType ),
    .io_toDecode_walkToArchVType ( io_toDecode_walkToArchVType ),
    .io_toDecode_walkVType_valid ( io_toDecode_walkVType_valid ),
    .io_toDecode_walkVType_bits_illegal ( io_toDecode_walkVType_bits_illegal ),
    .io_toDecode_walkVType_bits_vma ( io_toDecode_walkVType_bits_vma ),
    .io_toDecode_walkVType_bits_vta ( io_toDecode_walkVType_bits_vta ),
    .io_toDecode_walkVType_bits_vsew ( io_toDecode_walkVType_bits_vsew ),
    .io_toDecode_walkVType_bits_vlmul ( io_toDecode_walkVType_bits_vlmul ),
    .io_toDecode_commitVType_vtype_valid ( io_toDecode_commitVType_vtype_valid ),
    .io_toDecode_commitVType_vtype_bits_illegal ( io_toDecode_commitVType_vtype_bits_illegal ),
    .io_toDecode_commitVType_vtype_bits_vma ( io_toDecode_commitVType_vtype_bits_vma ),
    .io_toDecode_commitVType_vtype_bits_vta ( io_toDecode_commitVType_vtype_bits_vta ),
    .io_toDecode_commitVType_vtype_bits_vsew ( io_toDecode_commitVType_vtype_bits_vsew ),
    .io_toDecode_commitVType_vtype_bits_vlmul ( io_toDecode_commitVType_vtype_bits_vlmul ),
    .io_toDecode_commitVType_hasVsetvl ( io_toDecode_commitVType_hasVsetvl ),
    .io_readGPAMemAddr_valid ( io_readGPAMemAddr_valid ),
    .io_readGPAMemAddr_bits_ftqPtr_value ( io_readGPAMemAddr_bits_ftqPtr_value ),
    .io_readGPAMemAddr_bits_ftqOffset ( io_readGPAMemAddr_bits_ftqOffset ),
    .io_toVecExcpMod_logicPhyRegMap_0_valid ( io_toVecExcpMod_logicPhyRegMap_0_valid ),
    .io_toVecExcpMod_logicPhyRegMap_0_bits_lreg ( io_toVecExcpMod_logicPhyRegMap_0_bits_lreg ),
    .io_toVecExcpMod_logicPhyRegMap_0_bits_preg ( io_toVecExcpMod_logicPhyRegMap_0_bits_preg ),
    .io_toVecExcpMod_logicPhyRegMap_1_valid ( io_toVecExcpMod_logicPhyRegMap_1_valid ),
    .io_toVecExcpMod_logicPhyRegMap_1_bits_lreg ( io_toVecExcpMod_logicPhyRegMap_1_bits_lreg ),
    .io_toVecExcpMod_logicPhyRegMap_1_bits_preg ( io_toVecExcpMod_logicPhyRegMap_1_bits_preg ),
    .io_toVecExcpMod_logicPhyRegMap_2_valid ( io_toVecExcpMod_logicPhyRegMap_2_valid ),
    .io_toVecExcpMod_logicPhyRegMap_2_bits_lreg ( io_toVecExcpMod_logicPhyRegMap_2_bits_lreg ),
    .io_toVecExcpMod_logicPhyRegMap_2_bits_preg ( io_toVecExcpMod_logicPhyRegMap_2_bits_preg ),
    .io_toVecExcpMod_logicPhyRegMap_3_valid ( io_toVecExcpMod_logicPhyRegMap_3_valid ),
    .io_toVecExcpMod_logicPhyRegMap_3_bits_lreg ( io_toVecExcpMod_logicPhyRegMap_3_bits_lreg ),
    .io_toVecExcpMod_logicPhyRegMap_3_bits_preg ( io_toVecExcpMod_logicPhyRegMap_3_bits_preg ),
    .io_toVecExcpMod_logicPhyRegMap_4_valid ( io_toVecExcpMod_logicPhyRegMap_4_valid ),
    .io_toVecExcpMod_logicPhyRegMap_4_bits_lreg ( io_toVecExcpMod_logicPhyRegMap_4_bits_lreg ),
    .io_toVecExcpMod_logicPhyRegMap_4_bits_preg ( io_toVecExcpMod_logicPhyRegMap_4_bits_preg ),
    .io_toVecExcpMod_logicPhyRegMap_5_valid ( io_toVecExcpMod_logicPhyRegMap_5_valid ),
    .io_toVecExcpMod_logicPhyRegMap_5_bits_lreg ( io_toVecExcpMod_logicPhyRegMap_5_bits_lreg ),
    .io_toVecExcpMod_logicPhyRegMap_5_bits_preg ( io_toVecExcpMod_logicPhyRegMap_5_bits_preg ),
    .io_toVecExcpMod_excpInfo_valid ( io_toVecExcpMod_excpInfo_valid ),
    .io_toVecExcpMod_excpInfo_bits_vstart ( io_toVecExcpMod_excpInfo_bits_vstart ),
    .io_toVecExcpMod_excpInfo_bits_vsew ( io_toVecExcpMod_excpInfo_bits_vsew ),
    .io_toVecExcpMod_excpInfo_bits_veew ( io_toVecExcpMod_excpInfo_bits_veew ),
    .io_toVecExcpMod_excpInfo_bits_vlmul ( io_toVecExcpMod_excpInfo_bits_vlmul ),
    .io_toVecExcpMod_excpInfo_bits_nf ( io_toVecExcpMod_excpInfo_bits_nf ),
    .io_toVecExcpMod_excpInfo_bits_isStride ( io_toVecExcpMod_excpInfo_bits_isStride ),
    .io_toVecExcpMod_excpInfo_bits_isIndexed ( io_toVecExcpMod_excpInfo_bits_isIndexed ),
    .io_toVecExcpMod_excpInfo_bits_isWhole ( io_toVecExcpMod_excpInfo_bits_isWhole ),
    .io_toVecExcpMod_excpInfo_bits_isVlm ( io_toVecExcpMod_excpInfo_bits_isVlm ),
    .io_storeDebugInfo_1_pc ( io_storeDebugInfo_1_pc ),
    .io_perf_0_value      ( io_perf_0_value      ),
    .io_perf_1_value      ( io_perf_1_value      ),
    .io_perf_2_value      ( io_perf_2_value      ),
    .io_perf_3_value      ( io_perf_3_value      ),
    .io_perf_4_value      ( io_perf_4_value      ),
    .io_perf_5_value      ( io_perf_5_value      ),
    .io_perf_6_value      ( io_perf_6_value      ),
    .io_perf_7_value      ( io_perf_7_value      ),
    .io_perf_8_value      ( io_perf_8_value      ),
    .io_perf_9_value      ( io_perf_9_value      ),
    .io_perf_10_value     ( io_perf_10_value     ),
    .io_perf_11_value     ( io_perf_11_value     ),
    .io_perf_12_value     ( io_perf_12_value     ),
    .io_perf_13_value     ( io_perf_13_value     ),
    .io_perf_14_value     ( io_perf_14_value     ),
    .io_perf_15_value     ( io_perf_15_value     ),
    .io_perf_16_value     ( io_perf_16_value     ),
    .io_perf_17_value     ( io_perf_17_value     ),
    .io_error_0           ( io_error_0           )
);

`endif


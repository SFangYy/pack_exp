//=========================================================
//File name    : WriteBack_in_agent_monitor.sv
//Author       : nanyunhao
//Module name  : WriteBack_in_agent_monitor
//Discribution : WriteBack_in_agent_monitor : monitor
//Date         : 2026-01-22
//=========================================================
`ifndef WRITEBACK_IN_AGENT_MONITOR__SV
`define WRITEBACK_IN_AGENT_MONITOR__SV

class WriteBack_in_agent_monitor  extends tcnt_monitor_base#(virtual WriteBack_in_agent_interface,WriteBack_in_agent_cfg,WriteBack_in_agent_xaction);

    `uvm_component_utils(WriteBack_in_agent_monitor)

    extern function new(string name, uvm_component parent);
    extern virtual function void build_phase(uvm_phase phase);
    extern task run_phase(uvm_phase phase);
    extern task mon_data();
endclass:WriteBack_in_agent_monitor

function WriteBack_in_agent_monitor::new(string name, uvm_component parent);
    super.new(name,parent);
endfunction:new

function void WriteBack_in_agent_monitor::build_phase(uvm_phase phase);
    super.build_phase(phase);
endfunction:build_phase

task WriteBack_in_agent_monitor::run_phase(uvm_phase phase);
    super.run_phase(phase);
    this.mon_data();
endtask:run_phase

task WriteBack_in_agent_monitor::mon_data();

    logic         io_writeback_24_valid;
    logic [127:0] io_writeback_24_bits_data_0;
    logic [6:0]   io_writeback_24_bits_pdest;
    logic         io_writeback_24_bits_robIdx_flag;
    logic [7:0]   io_writeback_24_bits_robIdx_value;
    logic         io_writeback_24_bits_vecWen;
    logic         io_writeback_24_bits_v0Wen;
    logic         io_writeback_24_bits_vlWen;
    logic         io_writeback_24_bits_exceptionVec_0;
    logic         io_writeback_24_bits_exceptionVec_1;
    logic         io_writeback_24_bits_exceptionVec_2;
    logic         io_writeback_24_bits_exceptionVec_3;
    logic         io_writeback_24_bits_exceptionVec_4;
    logic         io_writeback_24_bits_exceptionVec_5;
    logic         io_writeback_24_bits_exceptionVec_6;
    logic         io_writeback_24_bits_exceptionVec_7;
    logic         io_writeback_24_bits_exceptionVec_8;
    logic         io_writeback_24_bits_exceptionVec_9;
    logic         io_writeback_24_bits_exceptionVec_10;
    logic         io_writeback_24_bits_exceptionVec_11;
    logic         io_writeback_24_bits_exceptionVec_12;
    logic         io_writeback_24_bits_exceptionVec_13;
    logic         io_writeback_24_bits_exceptionVec_14;
    logic         io_writeback_24_bits_exceptionVec_15;
    logic         io_writeback_24_bits_exceptionVec_16;
    logic         io_writeback_24_bits_exceptionVec_17;
    logic         io_writeback_24_bits_exceptionVec_18;
    logic         io_writeback_24_bits_exceptionVec_19;
    logic         io_writeback_24_bits_exceptionVec_20;
    logic         io_writeback_24_bits_exceptionVec_21;
    logic         io_writeback_24_bits_exceptionVec_22;
    logic         io_writeback_24_bits_exceptionVec_23;
    logic         io_writeback_24_bits_flushPipe;
    logic         io_writeback_24_bits_replay;
    logic [3:0]   io_writeback_24_bits_trigger;
    logic         io_writeback_24_bits_vls_vpu_vill;
    logic         io_writeback_24_bits_vls_vpu_vma;
    logic         io_writeback_24_bits_vls_vpu_vta;
    logic [1:0]   io_writeback_24_bits_vls_vpu_vsew;
    logic [2:0]   io_writeback_24_bits_vls_vpu_vlmul;
    logic         io_writeback_24_bits_vls_vpu_specVill;
    logic         io_writeback_24_bits_vls_vpu_specVma;
    logic         io_writeback_24_bits_vls_vpu_specVta;
    logic [1:0]   io_writeback_24_bits_vls_vpu_specVsew;
    logic [2:0]   io_writeback_24_bits_vls_vpu_specVlmul;
    logic         io_writeback_24_bits_vls_vpu_vm;
    logic [7:0]   io_writeback_24_bits_vls_vpu_vstart;
    logic [2:0]   io_writeback_24_bits_vls_vpu_frm;
    logic         io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst;
    logic         io_writeback_24_bits_vls_vpu_fpu_isFP32Instr;
    logic         io_writeback_24_bits_vls_vpu_fpu_isFP64Instr;
    logic         io_writeback_24_bits_vls_vpu_fpu_isReduction;
    logic         io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2;
    logic         io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4;
    logic         io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8;
    logic [1:0]   io_writeback_24_bits_vls_vpu_vxrm;
    logic [6:0]   io_writeback_24_bits_vls_vpu_vuopIdx;
    logic         io_writeback_24_bits_vls_vpu_lastUop;
    logic [127:0] io_writeback_24_bits_vls_vpu_vmask;
    logic [7:0]   io_writeback_24_bits_vls_vpu_vl;
    logic [2:0]   io_writeback_24_bits_vls_vpu_nf;
    logic [1:0]   io_writeback_24_bits_vls_vpu_veew;
    logic         io_writeback_24_bits_vls_vpu_isReverse;
    logic         io_writeback_24_bits_vls_vpu_isExt;
    logic         io_writeback_24_bits_vls_vpu_isNarrow;
    logic         io_writeback_24_bits_vls_vpu_isDstMask;
    logic         io_writeback_24_bits_vls_vpu_isOpMask;
    logic         io_writeback_24_bits_vls_vpu_isMove;
    logic         io_writeback_24_bits_vls_vpu_isDependOldVd;
    logic         io_writeback_24_bits_vls_vpu_isWritePartVd;
    logic         io_writeback_24_bits_vls_vpu_isVleff;
    logic [7:0]   io_writeback_24_bits_vls_oldVdPsrc;
    logic [2:0]   io_writeback_24_bits_vls_vdIdx;
    logic [2:0]   io_writeback_24_bits_vls_vdIdxInField;
    logic         io_writeback_24_bits_vls_isIndexed;
    logic         io_writeback_24_bits_vls_isMasked;
    logic         io_writeback_24_bits_vls_isStrided;
    logic         io_writeback_24_bits_vls_isWhole;
    logic         io_writeback_24_bits_vls_isVecLoad;
    logic         io_writeback_24_bits_vls_isVlm;
    logic         io_writeback_24_bits_debug_isMMIO;
    logic         io_writeback_24_bits_debug_isNCIO;
    logic         io_writeback_24_bits_debug_isPerfCnt;
    logic [47:0]  io_writeback_24_bits_debug_paddr;
    logic [49:0]  io_writeback_24_bits_debug_vaddr;
    logic         io_writeback_24_bits_debugInfo_eliminatedMove;
    logic [63:0]  io_writeback_24_bits_debugInfo_renameTime;
    logic [63:0]  io_writeback_24_bits_debugInfo_dispatchTime;
    logic [63:0]  io_writeback_24_bits_debugInfo_enqRsTime;
    logic [63:0]  io_writeback_24_bits_debugInfo_selectTime;
    logic [63:0]  io_writeback_24_bits_debugInfo_issueTime;
    logic [63:0]  io_writeback_24_bits_debugInfo_writebackTime;
    logic [63:0]  io_writeback_24_bits_debugInfo_runahead_checkpoint_id;
    logic [63:0]  io_writeback_24_bits_debugInfo_tlbFirstReqTime;
    logic [63:0]  io_writeback_24_bits_debugInfo_tlbRespTime;
    logic [63:0]  io_writeback_24_bits_debug_seqNum;
    logic         io_writeback_23_valid;
    logic [127:0] io_writeback_23_bits_data_0;
    logic [6:0]   io_writeback_23_bits_pdest;
    logic         io_writeback_23_bits_robIdx_flag;
    logic [7:0]   io_writeback_23_bits_robIdx_value;
    logic         io_writeback_23_bits_vecWen;
    logic         io_writeback_23_bits_v0Wen;
    logic         io_writeback_23_bits_vlWen;
    logic         io_writeback_23_bits_exceptionVec_0;
    logic         io_writeback_23_bits_exceptionVec_1;
    logic         io_writeback_23_bits_exceptionVec_2;
    logic         io_writeback_23_bits_exceptionVec_3;
    logic         io_writeback_23_bits_exceptionVec_4;
    logic         io_writeback_23_bits_exceptionVec_5;
    logic         io_writeback_23_bits_exceptionVec_6;
    logic         io_writeback_23_bits_exceptionVec_7;
    logic         io_writeback_23_bits_exceptionVec_8;
    logic         io_writeback_23_bits_exceptionVec_9;
    logic         io_writeback_23_bits_exceptionVec_10;
    logic         io_writeback_23_bits_exceptionVec_11;
    logic         io_writeback_23_bits_exceptionVec_12;
    logic         io_writeback_23_bits_exceptionVec_13;
    logic         io_writeback_23_bits_exceptionVec_14;
    logic         io_writeback_23_bits_exceptionVec_15;
    logic         io_writeback_23_bits_exceptionVec_16;
    logic         io_writeback_23_bits_exceptionVec_17;
    logic         io_writeback_23_bits_exceptionVec_18;
    logic         io_writeback_23_bits_exceptionVec_19;
    logic         io_writeback_23_bits_exceptionVec_20;
    logic         io_writeback_23_bits_exceptionVec_21;
    logic         io_writeback_23_bits_exceptionVec_22;
    logic         io_writeback_23_bits_exceptionVec_23;
    logic         io_writeback_23_bits_flushPipe;
    logic         io_writeback_23_bits_replay;
    logic [3:0]   io_writeback_23_bits_trigger;
    logic         io_writeback_23_bits_vls_vpu_vill;
    logic         io_writeback_23_bits_vls_vpu_vma;
    logic         io_writeback_23_bits_vls_vpu_vta;
    logic [1:0]   io_writeback_23_bits_vls_vpu_vsew;
    logic [2:0]   io_writeback_23_bits_vls_vpu_vlmul;
    logic         io_writeback_23_bits_vls_vpu_specVill;
    logic         io_writeback_23_bits_vls_vpu_specVma;
    logic         io_writeback_23_bits_vls_vpu_specVta;
    logic [1:0]   io_writeback_23_bits_vls_vpu_specVsew;
    logic [2:0]   io_writeback_23_bits_vls_vpu_specVlmul;
    logic         io_writeback_23_bits_vls_vpu_vm;
    logic [7:0]   io_writeback_23_bits_vls_vpu_vstart;
    logic [2:0]   io_writeback_23_bits_vls_vpu_frm;
    logic         io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst;
    logic         io_writeback_23_bits_vls_vpu_fpu_isFP32Instr;
    logic         io_writeback_23_bits_vls_vpu_fpu_isFP64Instr;
    logic         io_writeback_23_bits_vls_vpu_fpu_isReduction;
    logic         io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2;
    logic         io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4;
    logic         io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8;
    logic [1:0]   io_writeback_23_bits_vls_vpu_vxrm;
    logic [6:0]   io_writeback_23_bits_vls_vpu_vuopIdx;
    logic         io_writeback_23_bits_vls_vpu_lastUop;
    logic [127:0] io_writeback_23_bits_vls_vpu_vmask;
    logic [7:0]   io_writeback_23_bits_vls_vpu_vl;
    logic [2:0]   io_writeback_23_bits_vls_vpu_nf;
    logic [1:0]   io_writeback_23_bits_vls_vpu_veew;
    logic         io_writeback_23_bits_vls_vpu_isReverse;
    logic         io_writeback_23_bits_vls_vpu_isExt;
    logic         io_writeback_23_bits_vls_vpu_isNarrow;
    logic         io_writeback_23_bits_vls_vpu_isDstMask;
    logic         io_writeback_23_bits_vls_vpu_isOpMask;
    logic         io_writeback_23_bits_vls_vpu_isMove;
    logic         io_writeback_23_bits_vls_vpu_isDependOldVd;
    logic         io_writeback_23_bits_vls_vpu_isWritePartVd;
    logic         io_writeback_23_bits_vls_vpu_isVleff;
    logic [7:0]   io_writeback_23_bits_vls_oldVdPsrc;
    logic [2:0]   io_writeback_23_bits_vls_vdIdx;
    logic [2:0]   io_writeback_23_bits_vls_vdIdxInField;
    logic         io_writeback_23_bits_vls_isIndexed;
    logic         io_writeback_23_bits_vls_isMasked;
    logic         io_writeback_23_bits_vls_isStrided;
    logic         io_writeback_23_bits_vls_isWhole;
    logic         io_writeback_23_bits_vls_isVecLoad;
    logic         io_writeback_23_bits_vls_isVlm;
    logic         io_writeback_23_bits_debug_isMMIO;
    logic         io_writeback_23_bits_debug_isNCIO;
    logic         io_writeback_23_bits_debug_isPerfCnt;
    logic [47:0]  io_writeback_23_bits_debug_paddr;
    logic [49:0]  io_writeback_23_bits_debug_vaddr;
    logic         io_writeback_23_bits_debugInfo_eliminatedMove;
    logic [63:0]  io_writeback_23_bits_debugInfo_renameTime;
    logic [63:0]  io_writeback_23_bits_debugInfo_dispatchTime;
    logic [63:0]  io_writeback_23_bits_debugInfo_enqRsTime;
    logic [63:0]  io_writeback_23_bits_debugInfo_selectTime;
    logic [63:0]  io_writeback_23_bits_debugInfo_issueTime;
    logic [63:0]  io_writeback_23_bits_debugInfo_writebackTime;
    logic [63:0]  io_writeback_23_bits_debugInfo_runahead_checkpoint_id;
    logic [63:0]  io_writeback_23_bits_debugInfo_tlbFirstReqTime;
    logic [63:0]  io_writeback_23_bits_debugInfo_tlbRespTime;
    logic [63:0]  io_writeback_23_bits_debug_seqNum;
    logic         io_writeback_22_valid;
    logic [63:0]  io_writeback_22_bits_data_0;
    logic [7:0]   io_writeback_22_bits_pdest;
    logic         io_writeback_22_bits_robIdx_flag;
    logic [7:0]   io_writeback_22_bits_robIdx_value;
    logic         io_writeback_22_bits_intWen;
    logic         io_writeback_22_bits_fpWen;
    logic         io_writeback_22_bits_exceptionVec_0;
    logic         io_writeback_22_bits_exceptionVec_1;
    logic         io_writeback_22_bits_exceptionVec_2;
    logic         io_writeback_22_bits_exceptionVec_3;
    logic         io_writeback_22_bits_exceptionVec_4;
    logic         io_writeback_22_bits_exceptionVec_5;
    logic         io_writeback_22_bits_exceptionVec_6;
    logic         io_writeback_22_bits_exceptionVec_7;
    logic         io_writeback_22_bits_exceptionVec_8;
    logic         io_writeback_22_bits_exceptionVec_9;
    logic         io_writeback_22_bits_exceptionVec_10;
    logic         io_writeback_22_bits_exceptionVec_11;
    logic         io_writeback_22_bits_exceptionVec_12;
    logic         io_writeback_22_bits_exceptionVec_13;
    logic         io_writeback_22_bits_exceptionVec_14;
    logic         io_writeback_22_bits_exceptionVec_15;
    logic         io_writeback_22_bits_exceptionVec_16;
    logic         io_writeback_22_bits_exceptionVec_17;
    logic         io_writeback_22_bits_exceptionVec_18;
    logic         io_writeback_22_bits_exceptionVec_19;
    logic         io_writeback_22_bits_exceptionVec_20;
    logic         io_writeback_22_bits_exceptionVec_21;
    logic         io_writeback_22_bits_exceptionVec_22;
    logic         io_writeback_22_bits_exceptionVec_23;
    logic         io_writeback_22_bits_flushPipe;
    logic         io_writeback_22_bits_replay;
    logic         io_writeback_22_bits_lqIdx_flag;
    logic [6:0]   io_writeback_22_bits_lqIdx_value;
    logic [3:0]   io_writeback_22_bits_trigger;
    logic         io_writeback_22_bits_predecodeInfo_valid;
    logic         io_writeback_22_bits_predecodeInfo_isRVC;
    logic [1:0]   io_writeback_22_bits_predecodeInfo_brType;
    logic         io_writeback_22_bits_predecodeInfo_isCall;
    logic         io_writeback_22_bits_predecodeInfo_isRet;
    logic         io_writeback_22_bits_debug_isMMIO;
    logic         io_writeback_22_bits_debug_isNCIO;
    logic         io_writeback_22_bits_debug_isPerfCnt;
    logic [47:0]  io_writeback_22_bits_debug_paddr;
    logic [49:0]  io_writeback_22_bits_debug_vaddr;
    logic         io_writeback_22_bits_debugInfo_eliminatedMove;
    logic [63:0]  io_writeback_22_bits_debugInfo_renameTime;
    logic [63:0]  io_writeback_22_bits_debugInfo_dispatchTime;
    logic [63:0]  io_writeback_22_bits_debugInfo_enqRsTime;
    logic [63:0]  io_writeback_22_bits_debugInfo_selectTime;
    logic [63:0]  io_writeback_22_bits_debugInfo_issueTime;
    logic [63:0]  io_writeback_22_bits_debugInfo_writebackTime;
    logic [63:0]  io_writeback_22_bits_debugInfo_runahead_checkpoint_id;
    logic [63:0]  io_writeback_22_bits_debugInfo_tlbFirstReqTime;
    logic [63:0]  io_writeback_22_bits_debugInfo_tlbRespTime;
    logic [63:0]  io_writeback_22_bits_debug_seqNum;
    logic         io_writeback_21_valid;
    logic [63:0]  io_writeback_21_bits_data_0;
    logic [7:0]   io_writeback_21_bits_pdest;
    logic         io_writeback_21_bits_robIdx_flag;
    logic [7:0]   io_writeback_21_bits_robIdx_value;
    logic         io_writeback_21_bits_intWen;
    logic         io_writeback_21_bits_fpWen;
    logic         io_writeback_21_bits_exceptionVec_0;
    logic         io_writeback_21_bits_exceptionVec_1;
    logic         io_writeback_21_bits_exceptionVec_2;
    logic         io_writeback_21_bits_exceptionVec_3;
    logic         io_writeback_21_bits_exceptionVec_4;
    logic         io_writeback_21_bits_exceptionVec_5;
    logic         io_writeback_21_bits_exceptionVec_6;
    logic         io_writeback_21_bits_exceptionVec_7;
    logic         io_writeback_21_bits_exceptionVec_8;
    logic         io_writeback_21_bits_exceptionVec_9;
    logic         io_writeback_21_bits_exceptionVec_10;
    logic         io_writeback_21_bits_exceptionVec_11;
    logic         io_writeback_21_bits_exceptionVec_12;
    logic         io_writeback_21_bits_exceptionVec_13;
    logic         io_writeback_21_bits_exceptionVec_14;
    logic         io_writeback_21_bits_exceptionVec_15;
    logic         io_writeback_21_bits_exceptionVec_16;
    logic         io_writeback_21_bits_exceptionVec_17;
    logic         io_writeback_21_bits_exceptionVec_18;
    logic         io_writeback_21_bits_exceptionVec_19;
    logic         io_writeback_21_bits_exceptionVec_20;
    logic         io_writeback_21_bits_exceptionVec_21;
    logic         io_writeback_21_bits_exceptionVec_22;
    logic         io_writeback_21_bits_exceptionVec_23;
    logic         io_writeback_21_bits_flushPipe;
    logic         io_writeback_21_bits_replay;
    logic         io_writeback_21_bits_lqIdx_flag;
    logic [6:0]   io_writeback_21_bits_lqIdx_value;
    logic [3:0]   io_writeback_21_bits_trigger;
    logic         io_writeback_21_bits_predecodeInfo_valid;
    logic         io_writeback_21_bits_predecodeInfo_isRVC;
    logic [1:0]   io_writeback_21_bits_predecodeInfo_brType;
    logic         io_writeback_21_bits_predecodeInfo_isCall;
    logic         io_writeback_21_bits_predecodeInfo_isRet;
    logic         io_writeback_21_bits_debug_isMMIO;
    logic         io_writeback_21_bits_debug_isNCIO;
    logic         io_writeback_21_bits_debug_isPerfCnt;
    logic [47:0]  io_writeback_21_bits_debug_paddr;
    logic [49:0]  io_writeback_21_bits_debug_vaddr;
    logic         io_writeback_21_bits_debugInfo_eliminatedMove;
    logic [63:0]  io_writeback_21_bits_debugInfo_renameTime;
    logic [63:0]  io_writeback_21_bits_debugInfo_dispatchTime;
    logic [63:0]  io_writeback_21_bits_debugInfo_enqRsTime;
    logic [63:0]  io_writeback_21_bits_debugInfo_selectTime;
    logic [63:0]  io_writeback_21_bits_debugInfo_issueTime;
    logic [63:0]  io_writeback_21_bits_debugInfo_writebackTime;
    logic [63:0]  io_writeback_21_bits_debugInfo_runahead_checkpoint_id;
    logic [63:0]  io_writeback_21_bits_debugInfo_tlbFirstReqTime;
    logic [63:0]  io_writeback_21_bits_debugInfo_tlbRespTime;
    logic [63:0]  io_writeback_21_bits_debug_seqNum;
    logic         io_writeback_20_valid;
    logic [63:0]  io_writeback_20_bits_data_0;
    logic [7:0]   io_writeback_20_bits_pdest;
    logic         io_writeback_20_bits_robIdx_flag;
    logic [7:0]   io_writeback_20_bits_robIdx_value;
    logic         io_writeback_20_bits_intWen;
    logic         io_writeback_20_bits_fpWen;
    logic         io_writeback_20_bits_exceptionVec_0;
    logic         io_writeback_20_bits_exceptionVec_1;
    logic         io_writeback_20_bits_exceptionVec_2;
    logic         io_writeback_20_bits_exceptionVec_3;
    logic         io_writeback_20_bits_exceptionVec_4;
    logic         io_writeback_20_bits_exceptionVec_5;
    logic         io_writeback_20_bits_exceptionVec_6;
    logic         io_writeback_20_bits_exceptionVec_7;
    logic         io_writeback_20_bits_exceptionVec_8;
    logic         io_writeback_20_bits_exceptionVec_9;
    logic         io_writeback_20_bits_exceptionVec_10;
    logic         io_writeback_20_bits_exceptionVec_11;
    logic         io_writeback_20_bits_exceptionVec_12;
    logic         io_writeback_20_bits_exceptionVec_13;
    logic         io_writeback_20_bits_exceptionVec_14;
    logic         io_writeback_20_bits_exceptionVec_15;
    logic         io_writeback_20_bits_exceptionVec_16;
    logic         io_writeback_20_bits_exceptionVec_17;
    logic         io_writeback_20_bits_exceptionVec_18;
    logic         io_writeback_20_bits_exceptionVec_19;
    logic         io_writeback_20_bits_exceptionVec_20;
    logic         io_writeback_20_bits_exceptionVec_21;
    logic         io_writeback_20_bits_exceptionVec_22;
    logic         io_writeback_20_bits_exceptionVec_23;
    logic         io_writeback_20_bits_flushPipe;
    logic         io_writeback_20_bits_replay;
    logic         io_writeback_20_bits_lqIdx_flag;
    logic [6:0]   io_writeback_20_bits_lqIdx_value;
    logic [3:0]   io_writeback_20_bits_trigger;
    logic         io_writeback_20_bits_predecodeInfo_valid;
    logic         io_writeback_20_bits_predecodeInfo_isRVC;
    logic [1:0]   io_writeback_20_bits_predecodeInfo_brType;
    logic         io_writeback_20_bits_predecodeInfo_isCall;
    logic         io_writeback_20_bits_predecodeInfo_isRet;
    logic         io_writeback_20_bits_debug_isMMIO;
    logic         io_writeback_20_bits_debug_isNCIO;
    logic         io_writeback_20_bits_debug_isPerfCnt;
    logic [47:0]  io_writeback_20_bits_debug_paddr;
    logic [49:0]  io_writeback_20_bits_debug_vaddr;
    logic         io_writeback_20_bits_debugInfo_eliminatedMove;
    logic [63:0]  io_writeback_20_bits_debugInfo_renameTime;
    logic [63:0]  io_writeback_20_bits_debugInfo_dispatchTime;
    logic [63:0]  io_writeback_20_bits_debugInfo_enqRsTime;
    logic [63:0]  io_writeback_20_bits_debugInfo_selectTime;
    logic [63:0]  io_writeback_20_bits_debugInfo_issueTime;
    logic [63:0]  io_writeback_20_bits_debugInfo_writebackTime;
    logic [63:0]  io_writeback_20_bits_debugInfo_runahead_checkpoint_id;
    logic [63:0]  io_writeback_20_bits_debugInfo_tlbFirstReqTime;
    logic [63:0]  io_writeback_20_bits_debugInfo_tlbRespTime;
    logic [63:0]  io_writeback_20_bits_debug_seqNum;
    logic         io_writeback_19_valid;
    logic [63:0]  io_writeback_19_bits_data_0;
    logic [7:0]   io_writeback_19_bits_pdest;
    logic         io_writeback_19_bits_robIdx_flag;
    logic [7:0]   io_writeback_19_bits_robIdx_value;
    logic         io_writeback_19_bits_intWen;
    logic         io_writeback_19_bits_exceptionVec_0;
    logic         io_writeback_19_bits_exceptionVec_1;
    logic         io_writeback_19_bits_exceptionVec_2;
    logic         io_writeback_19_bits_exceptionVec_3;
    logic         io_writeback_19_bits_exceptionVec_4;
    logic         io_writeback_19_bits_exceptionVec_5;
    logic         io_writeback_19_bits_exceptionVec_6;
    logic         io_writeback_19_bits_exceptionVec_7;
    logic         io_writeback_19_bits_exceptionVec_8;
    logic         io_writeback_19_bits_exceptionVec_9;
    logic         io_writeback_19_bits_exceptionVec_10;
    logic         io_writeback_19_bits_exceptionVec_11;
    logic         io_writeback_19_bits_exceptionVec_12;
    logic         io_writeback_19_bits_exceptionVec_13;
    logic         io_writeback_19_bits_exceptionVec_14;
    logic         io_writeback_19_bits_exceptionVec_15;
    logic         io_writeback_19_bits_exceptionVec_16;
    logic         io_writeback_19_bits_exceptionVec_17;
    logic         io_writeback_19_bits_exceptionVec_18;
    logic         io_writeback_19_bits_exceptionVec_19;
    logic         io_writeback_19_bits_exceptionVec_20;
    logic         io_writeback_19_bits_exceptionVec_21;
    logic         io_writeback_19_bits_exceptionVec_22;
    logic         io_writeback_19_bits_exceptionVec_23;
    logic         io_writeback_19_bits_flushPipe;
    logic         io_writeback_19_bits_sqIdx_flag;
    logic [5:0]   io_writeback_19_bits_sqIdx_value;
    logic [3:0]   io_writeback_19_bits_trigger;
    logic         io_writeback_19_bits_debug_isMMIO;
    logic         io_writeback_19_bits_debug_isNCIO;
    logic         io_writeback_19_bits_debug_isPerfCnt;
    logic [47:0]  io_writeback_19_bits_debug_paddr;
    logic [49:0]  io_writeback_19_bits_debug_vaddr;
    logic         io_writeback_19_bits_debugInfo_eliminatedMove;
    logic [63:0]  io_writeback_19_bits_debugInfo_renameTime;
    logic [63:0]  io_writeback_19_bits_debugInfo_dispatchTime;
    logic [63:0]  io_writeback_19_bits_debugInfo_enqRsTime;
    logic [63:0]  io_writeback_19_bits_debugInfo_selectTime;
    logic [63:0]  io_writeback_19_bits_debugInfo_issueTime;
    logic [63:0]  io_writeback_19_bits_debugInfo_writebackTime;
    logic [63:0]  io_writeback_19_bits_debugInfo_runahead_checkpoint_id;
    logic [63:0]  io_writeback_19_bits_debugInfo_tlbFirstReqTime;
    logic [63:0]  io_writeback_19_bits_debugInfo_tlbRespTime;
    logic [63:0]  io_writeback_19_bits_debug_seqNum;
    logic         io_writeback_18_valid;
    logic [63:0]  io_writeback_18_bits_data_0;
    logic [7:0]   io_writeback_18_bits_pdest;
    logic         io_writeback_18_bits_robIdx_flag;
    logic [7:0]   io_writeback_18_bits_robIdx_value;
    logic         io_writeback_18_bits_intWen;
    logic         io_writeback_18_bits_exceptionVec_0;
    logic         io_writeback_18_bits_exceptionVec_1;
    logic         io_writeback_18_bits_exceptionVec_2;
    logic         io_writeback_18_bits_exceptionVec_3;
    logic         io_writeback_18_bits_exceptionVec_4;
    logic         io_writeback_18_bits_exceptionVec_5;
    logic         io_writeback_18_bits_exceptionVec_6;
    logic         io_writeback_18_bits_exceptionVec_7;
    logic         io_writeback_18_bits_exceptionVec_8;
    logic         io_writeback_18_bits_exceptionVec_9;
    logic         io_writeback_18_bits_exceptionVec_10;
    logic         io_writeback_18_bits_exceptionVec_11;
    logic         io_writeback_18_bits_exceptionVec_12;
    logic         io_writeback_18_bits_exceptionVec_13;
    logic         io_writeback_18_bits_exceptionVec_14;
    logic         io_writeback_18_bits_exceptionVec_15;
    logic         io_writeback_18_bits_exceptionVec_16;
    logic         io_writeback_18_bits_exceptionVec_17;
    logic         io_writeback_18_bits_exceptionVec_18;
    logic         io_writeback_18_bits_exceptionVec_19;
    logic         io_writeback_18_bits_exceptionVec_20;
    logic         io_writeback_18_bits_exceptionVec_21;
    logic         io_writeback_18_bits_exceptionVec_22;
    logic         io_writeback_18_bits_exceptionVec_23;
    logic         io_writeback_18_bits_flushPipe;
    logic         io_writeback_18_bits_sqIdx_flag;
    logic [5:0]   io_writeback_18_bits_sqIdx_value;
    logic [3:0]   io_writeback_18_bits_trigger;
    logic         io_writeback_18_bits_debug_isMMIO;
    logic         io_writeback_18_bits_debug_isNCIO;
    logic         io_writeback_18_bits_debug_isPerfCnt;
    logic [47:0]  io_writeback_18_bits_debug_paddr;
    logic [49:0]  io_writeback_18_bits_debug_vaddr;
    logic         io_writeback_18_bits_debugInfo_eliminatedMove;
    logic [63:0]  io_writeback_18_bits_debugInfo_renameTime;
    logic [63:0]  io_writeback_18_bits_debugInfo_dispatchTime;
    logic [63:0]  io_writeback_18_bits_debugInfo_enqRsTime;
    logic [63:0]  io_writeback_18_bits_debugInfo_selectTime;
    logic [63:0]  io_writeback_18_bits_debugInfo_issueTime;
    logic [63:0]  io_writeback_18_bits_debugInfo_writebackTime;
    logic [63:0]  io_writeback_18_bits_debugInfo_runahead_checkpoint_id;
    logic [63:0]  io_writeback_18_bits_debugInfo_tlbFirstReqTime;
    logic [63:0]  io_writeback_18_bits_debugInfo_tlbRespTime;
    logic [63:0]  io_writeback_18_bits_debug_seqNum;
    logic         io_writeback_17_valid;
    logic [127:0] io_writeback_17_bits_data_0;
    logic [127:0] io_writeback_17_bits_data_1;
    logic [127:0] io_writeback_17_bits_data_2;
    logic [6:0]   io_writeback_17_bits_pdest;
    logic         io_writeback_17_bits_robIdx_flag;
    logic [7:0]   io_writeback_17_bits_robIdx_value;
    logic         io_writeback_17_bits_vecWen;
    logic         io_writeback_17_bits_v0Wen;
    logic [4:0]   io_writeback_17_bits_fflags;
    logic         io_writeback_17_bits_wflags;
    logic         io_writeback_17_bits_debugInfo_eliminatedMove;
    logic [63:0]  io_writeback_17_bits_debugInfo_renameTime;
    logic [63:0]  io_writeback_17_bits_debugInfo_dispatchTime;
    logic [63:0]  io_writeback_17_bits_debugInfo_enqRsTime;
    logic [63:0]  io_writeback_17_bits_debugInfo_selectTime;
    logic [63:0]  io_writeback_17_bits_debugInfo_issueTime;
    logic [63:0]  io_writeback_17_bits_debugInfo_writebackTime;
    logic [63:0]  io_writeback_17_bits_debugInfo_runahead_checkpoint_id;
    logic [63:0]  io_writeback_17_bits_debugInfo_tlbFirstReqTime;
    logic [63:0]  io_writeback_17_bits_debugInfo_tlbRespTime;
    logic [63:0]  io_writeback_17_bits_debug_seqNum;
    logic         io_writeback_16_valid;
    logic [127:0] io_writeback_16_bits_data_0;
    logic [127:0] io_writeback_16_bits_data_1;
    logic [127:0] io_writeback_16_bits_data_2;
    logic [127:0] io_writeback_16_bits_data_3;
    logic [7:0]   io_writeback_16_bits_pdest;
    logic         io_writeback_16_bits_robIdx_flag;
    logic [7:0]   io_writeback_16_bits_robIdx_value;
    logic         io_writeback_16_bits_fpWen;
    logic         io_writeback_16_bits_vecWen;
    logic         io_writeback_16_bits_v0Wen;
    logic [4:0]   io_writeback_16_bits_fflags;
    logic         io_writeback_16_bits_wflags;
    logic         io_writeback_16_bits_debugInfo_eliminatedMove;
    logic [63:0]  io_writeback_16_bits_debugInfo_renameTime;
    logic [63:0]  io_writeback_16_bits_debugInfo_dispatchTime;
    logic [63:0]  io_writeback_16_bits_debugInfo_enqRsTime;
    logic [63:0]  io_writeback_16_bits_debugInfo_selectTime;
    logic [63:0]  io_writeback_16_bits_debugInfo_issueTime;
    logic [63:0]  io_writeback_16_bits_debugInfo_writebackTime;
    logic [63:0]  io_writeback_16_bits_debugInfo_runahead_checkpoint_id;
    logic [63:0]  io_writeback_16_bits_debugInfo_tlbFirstReqTime;
    logic [63:0]  io_writeback_16_bits_debugInfo_tlbRespTime;
    logic [63:0]  io_writeback_16_bits_debug_seqNum;
    logic         io_writeback_15_valid;
    logic [127:0] io_writeback_15_bits_data_0;
    logic [127:0] io_writeback_15_bits_data_1;
    logic [127:0] io_writeback_15_bits_data_2;
    logic [6:0]   io_writeback_15_bits_pdest;
    logic         io_writeback_15_bits_robIdx_flag;
    logic [7:0]   io_writeback_15_bits_robIdx_value;
    logic         io_writeback_15_bits_vecWen;
    logic         io_writeback_15_bits_v0Wen;
    logic [4:0]   io_writeback_15_bits_fflags;
    logic         io_writeback_15_bits_wflags;
    logic         io_writeback_15_bits_vxsat;
    logic         io_writeback_15_bits_debugInfo_eliminatedMove;
    logic [63:0]  io_writeback_15_bits_debugInfo_renameTime;
    logic [63:0]  io_writeback_15_bits_debugInfo_dispatchTime;
    logic [63:0]  io_writeback_15_bits_debugInfo_enqRsTime;
    logic [63:0]  io_writeback_15_bits_debugInfo_selectTime;
    logic [63:0]  io_writeback_15_bits_debugInfo_issueTime;
    logic [63:0]  io_writeback_15_bits_debugInfo_writebackTime;
    logic [63:0]  io_writeback_15_bits_debugInfo_runahead_checkpoint_id;
    logic [63:0]  io_writeback_15_bits_debugInfo_tlbFirstReqTime;
    logic [63:0]  io_writeback_15_bits_debugInfo_tlbRespTime;
    logic [63:0]  io_writeback_15_bits_debug_seqNum;
    logic         io_writeback_14_valid;
    logic [127:0] io_writeback_14_bits_data_0;
    logic [127:0] io_writeback_14_bits_data_1;
    logic [127:0] io_writeback_14_bits_data_2;
    logic [127:0] io_writeback_14_bits_data_3;
    logic [127:0] io_writeback_14_bits_data_4;
    logic [127:0] io_writeback_14_bits_data_5;
    logic [7:0]   io_writeback_14_bits_pdest;
    logic         io_writeback_14_bits_robIdx_flag;
    logic [7:0]   io_writeback_14_bits_robIdx_value;
    logic         io_writeback_14_bits_intWen;
    logic         io_writeback_14_bits_fpWen;
    logic         io_writeback_14_bits_vecWen;
    logic         io_writeback_14_bits_v0Wen;
    logic         io_writeback_14_bits_vlWen;
    logic [4:0]   io_writeback_14_bits_fflags;
    logic         io_writeback_14_bits_wflags;
    logic         io_writeback_14_bits_exceptionVec_2;
    logic         io_writeback_14_bits_debugInfo_eliminatedMove;
    logic [63:0]  io_writeback_14_bits_debugInfo_renameTime;
    logic [63:0]  io_writeback_14_bits_debugInfo_dispatchTime;
    logic [63:0]  io_writeback_14_bits_debugInfo_enqRsTime;
    logic [63:0]  io_writeback_14_bits_debugInfo_selectTime;
    logic [63:0]  io_writeback_14_bits_debugInfo_issueTime;
    logic [63:0]  io_writeback_14_bits_debugInfo_writebackTime;
    logic [63:0]  io_writeback_14_bits_debugInfo_runahead_checkpoint_id;
    logic [63:0]  io_writeback_14_bits_debugInfo_tlbFirstReqTime;
    logic [63:0]  io_writeback_14_bits_debugInfo_tlbRespTime;
    logic [63:0]  io_writeback_14_bits_debug_seqNum;
    logic         io_writeback_13_valid;
    logic [127:0] io_writeback_13_bits_data_0;
    logic [127:0] io_writeback_13_bits_data_1;
    logic [127:0] io_writeback_13_bits_data_2;
    logic [6:0]   io_writeback_13_bits_pdest;
    logic         io_writeback_13_bits_robIdx_flag;
    logic [7:0]   io_writeback_13_bits_robIdx_value;
    logic         io_writeback_13_bits_vecWen;
    logic         io_writeback_13_bits_v0Wen;
    logic [4:0]   io_writeback_13_bits_fflags;
    logic         io_writeback_13_bits_wflags;
    logic         io_writeback_13_bits_vxsat;
    logic         io_writeback_13_bits_exceptionVec_2;
    logic         io_writeback_13_bits_debugInfo_eliminatedMove;
    logic [63:0]  io_writeback_13_bits_debugInfo_renameTime;
    logic [63:0]  io_writeback_13_bits_debugInfo_dispatchTime;
    logic [63:0]  io_writeback_13_bits_debugInfo_enqRsTime;
    logic [63:0]  io_writeback_13_bits_debugInfo_selectTime;
    logic [63:0]  io_writeback_13_bits_debugInfo_issueTime;
    logic [63:0]  io_writeback_13_bits_debugInfo_writebackTime;
    logic [63:0]  io_writeback_13_bits_debugInfo_runahead_checkpoint_id;
    logic [63:0]  io_writeback_13_bits_debugInfo_tlbFirstReqTime;
    logic [63:0]  io_writeback_13_bits_debugInfo_tlbRespTime;
    logic [63:0]  io_writeback_13_bits_debug_seqNum;
    logic         io_writeback_7_valid ;
    logic [63:0]  io_writeback_7_bits_data_0;
    logic [63:0]  io_writeback_7_bits_data_1;
    logic [7:0]   io_writeback_7_bits_pdest;
    logic         io_writeback_7_bits_robIdx_flag;
    logic [7:0]   io_writeback_7_bits_robIdx_value;
    logic         io_writeback_7_bits_intWen;
    logic         io_writeback_7_bits_redirect_valid;
    logic         io_writeback_7_bits_redirect_bits_isRVC;
    logic         io_writeback_7_bits_redirect_bits_robIdx_flag;
    logic [7:0]   io_writeback_7_bits_redirect_bits_robIdx_value;
    logic         io_writeback_7_bits_redirect_bits_ftqIdx_flag;
    logic [5:0]   io_writeback_7_bits_redirect_bits_ftqIdx_value;
    logic [3:0]   io_writeback_7_bits_redirect_bits_ftqOffset;
    logic         io_writeback_7_bits_redirect_bits_level;
    logic         io_writeback_7_bits_redirect_bits_interrupt;
    logic [49:0]  io_writeback_7_bits_redirect_bits_cfiUpdate_pc;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC;
    logic [1:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet;
    logic [3:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_ssp;
    logic [2:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_sctr;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag;
    logic [4:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag;
    logic [4:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag;
    logic [4:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value;
    logic [49:0]  io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr;
    logic [10:0]  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist;
    logic [10:0]  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist;
    logic [6:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist;
    logic [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist;
    logic [8:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist;
    logic [3:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist;
    logic [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist;
    logic [8:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist;
    logic [6:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist;
    logic [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist;
    logic [6:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist;
    logic [8:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist;
    logic [6:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist;
    logic [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist;
    logic [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist;
    logic [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist;
    logic [10:0]  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist;
    logic [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3;
    logic [2:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH;
    logic [3:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_ghr;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag;
    logic [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value;
    logic [9:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0;
    logic [9:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken;
    logic [49:0]  io_writeback_7_bits_redirect_bits_cfiUpdate_target;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_taken;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred;
    logic [1:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_shift;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF;
    logic [63:0]  io_writeback_7_bits_redirect_bits_fullTarget;
    logic         io_writeback_7_bits_redirect_bits_stFtqIdx_flag;
    logic [5:0]   io_writeback_7_bits_redirect_bits_stFtqIdx_value;
    logic [3:0]   io_writeback_7_bits_redirect_bits_stFtqOffset;
    logic [63:0]  io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id;
    logic         io_writeback_7_bits_redirect_bits_debugIsCtrl;
    logic         io_writeback_7_bits_redirect_bits_debugIsMemVio;
    logic         io_writeback_7_bits_exceptionVec_2;
    logic         io_writeback_7_bits_exceptionVec_3;
    logic         io_writeback_7_bits_exceptionVec_8;
    logic         io_writeback_7_bits_exceptionVec_9;
    logic         io_writeback_7_bits_exceptionVec_10;
    logic         io_writeback_7_bits_exceptionVec_11;
    logic         io_writeback_7_bits_exceptionVec_22;
    logic         io_writeback_7_bits_flushPipe;
    logic         io_writeback_7_bits_predecodeInfo_valid;
    logic         io_writeback_7_bits_predecodeInfo_isRVC;
    logic [1:0]   io_writeback_7_bits_predecodeInfo_brType;
    logic         io_writeback_7_bits_predecodeInfo_isCall;
    logic         io_writeback_7_bits_predecodeInfo_isRet;
    logic         io_writeback_7_bits_debug_isPerfCnt;
    logic         io_writeback_7_bits_debugInfo_eliminatedMove;
    logic [63:0]  io_writeback_7_bits_debugInfo_renameTime;
    logic [63:0]  io_writeback_7_bits_debugInfo_dispatchTime;
    logic [63:0]  io_writeback_7_bits_debugInfo_enqRsTime;
    logic [63:0]  io_writeback_7_bits_debugInfo_selectTime;
    logic [63:0]  io_writeback_7_bits_debugInfo_issueTime;
    logic [63:0]  io_writeback_7_bits_debugInfo_writebackTime;
    logic [63:0]  io_writeback_7_bits_debugInfo_runahead_checkpoint_id;
    logic [63:0]  io_writeback_7_bits_debugInfo_tlbFirstReqTime;
    logic [63:0]  io_writeback_7_bits_debugInfo_tlbRespTime;
    logic [63:0]  io_writeback_7_bits_debug_seqNum;
    logic         io_writeback_5_valid ;
    logic         io_writeback_5_bits_redirect_valid;
    logic         io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred;
    logic         io_writeback_3_valid ;
    logic         io_writeback_3_bits_redirect_valid;
    logic         io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred;
    logic         io_writeback_1_valid ;
    logic         io_writeback_1_bits_redirect_valid;
    logic         io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred;
    logic         io_exuWriteback_26_valid;
    logic [7:0]   io_exuWriteback_26_bits_robIdx_value;
    logic         io_exuWriteback_25_valid;
    logic [7:0]   io_exuWriteback_25_bits_robIdx_value;
    logic         io_exuWriteback_24_valid;
    logic [127:0] io_exuWriteback_24_bits_data_0;
    logic [6:0]   io_exuWriteback_24_bits_pdest;
    logic [7:0]   io_exuWriteback_24_bits_robIdx_value;
    logic         io_exuWriteback_24_bits_vecWen;
    logic         io_exuWriteback_24_bits_v0Wen;
    logic [2:0]   io_exuWriteback_24_bits_vls_vdIdx;
    logic         io_exuWriteback_24_bits_debug_isMMIO;
    logic         io_exuWriteback_24_bits_debug_isNCIO;
    logic         io_exuWriteback_24_bits_debug_isPerfCnt;
    logic [47:0]  io_exuWriteback_24_bits_debug_paddr;
    logic         io_exuWriteback_23_valid;
    logic [127:0] io_exuWriteback_23_bits_data_0;
    logic [6:0]   io_exuWriteback_23_bits_pdest;
    logic [7:0]   io_exuWriteback_23_bits_robIdx_value;
    logic         io_exuWriteback_23_bits_vecWen;
    logic         io_exuWriteback_23_bits_v0Wen;
    logic [2:0]   io_exuWriteback_23_bits_vls_vdIdx;
    logic         io_exuWriteback_23_bits_debug_isMMIO;
    logic         io_exuWriteback_23_bits_debug_isNCIO;
    logic         io_exuWriteback_23_bits_debug_isPerfCnt;
    logic [47:0]  io_exuWriteback_23_bits_debug_paddr;
    logic         io_exuWriteback_22_valid;
    logic [63:0]  io_exuWriteback_22_bits_data_0;
    logic [7:0]   io_exuWriteback_22_bits_robIdx_value;
    logic [6:0]   io_exuWriteback_22_bits_lqIdx_value;
    logic         io_exuWriteback_22_bits_debug_isMMIO;
    logic         io_exuWriteback_22_bits_debug_isNCIO;
    logic         io_exuWriteback_22_bits_debug_isPerfCnt;
    logic [47:0]  io_exuWriteback_22_bits_debug_paddr;
    logic         io_exuWriteback_21_valid;
    logic [63:0]  io_exuWriteback_21_bits_data_0;
    logic [7:0]   io_exuWriteback_21_bits_robIdx_value;
    logic [6:0]   io_exuWriteback_21_bits_lqIdx_value;
    logic         io_exuWriteback_21_bits_debug_isMMIO;
    logic         io_exuWriteback_21_bits_debug_isNCIO;
    logic         io_exuWriteback_21_bits_debug_isPerfCnt;
    logic [47:0]  io_exuWriteback_21_bits_debug_paddr;
    logic         io_exuWriteback_20_valid;
    logic [63:0]  io_exuWriteback_20_bits_data_0;
    logic [7:0]   io_exuWriteback_20_bits_robIdx_value;
    logic [6:0]   io_exuWriteback_20_bits_lqIdx_value;
    logic         io_exuWriteback_20_bits_debug_isMMIO;
    logic         io_exuWriteback_20_bits_debug_isNCIO;
    logic         io_exuWriteback_20_bits_debug_isPerfCnt;
    logic [47:0]  io_exuWriteback_20_bits_debug_paddr;
    logic         io_exuWriteback_19_valid;
    logic [63:0]  io_exuWriteback_19_bits_data_0;
    logic [7:0]   io_exuWriteback_19_bits_robIdx_value;
    logic [5:0]   io_exuWriteback_19_bits_sqIdx_value;
    logic         io_exuWriteback_19_bits_debug_isMMIO;
    logic         io_exuWriteback_19_bits_debug_isNCIO;
    logic         io_exuWriteback_19_bits_debug_isPerfCnt;
    logic [47:0]  io_exuWriteback_19_bits_debug_paddr;
    logic         io_exuWriteback_18_valid;
    logic [63:0]  io_exuWriteback_18_bits_data_0;
    logic [7:0]   io_exuWriteback_18_bits_robIdx_value;
    logic [5:0]   io_exuWriteback_18_bits_sqIdx_value;
    logic         io_exuWriteback_18_bits_debug_isMMIO;
    logic         io_exuWriteback_18_bits_debug_isNCIO;
    logic         io_exuWriteback_18_bits_debug_isPerfCnt;
    logic [47:0]  io_exuWriteback_18_bits_debug_paddr;
    logic         io_exuWriteback_17_valid;
    logic [127:0] io_exuWriteback_17_bits_data_0;
    logic [7:0]   io_exuWriteback_17_bits_robIdx_value;
    logic [4:0]   io_exuWriteback_17_bits_fflags;
    logic         io_exuWriteback_17_bits_wflags;
    logic         io_exuWriteback_16_valid;
    logic [127:0] io_exuWriteback_16_bits_data_0;
    logic [7:0]   io_exuWriteback_16_bits_robIdx_value;
    logic [4:0]   io_exuWriteback_16_bits_fflags;
    logic         io_exuWriteback_16_bits_wflags;
    logic         io_exuWriteback_15_valid;
    logic [127:0] io_exuWriteback_15_bits_data_0;
    logic [7:0]   io_exuWriteback_15_bits_robIdx_value;
    logic [4:0]   io_exuWriteback_15_bits_fflags;
    logic         io_exuWriteback_15_bits_wflags;
    logic         io_exuWriteback_15_bits_vxsat;
    logic         io_exuWriteback_14_valid;
    logic [127:0] io_exuWriteback_14_bits_data_0;
    logic [7:0]   io_exuWriteback_14_bits_robIdx_value;
    logic [4:0]   io_exuWriteback_14_bits_fflags;
    logic         io_exuWriteback_14_bits_wflags;
    logic         io_exuWriteback_13_valid;
    logic [127:0] io_exuWriteback_13_bits_data_0;
    logic [7:0]   io_exuWriteback_13_bits_robIdx_value;
    logic [4:0]   io_exuWriteback_13_bits_fflags;
    logic         io_exuWriteback_13_bits_wflags;
    logic         io_exuWriteback_13_bits_vxsat;
    logic         io_exuWriteback_12_valid;
    logic [63:0]  io_exuWriteback_12_bits_data_0;
    logic [7:0]   io_exuWriteback_12_bits_robIdx_value;
    logic [4:0]   io_exuWriteback_12_bits_fflags;
    logic         io_exuWriteback_12_bits_wflags;
    logic         io_exuWriteback_11_valid;
    logic [63:0]  io_exuWriteback_11_bits_data_0;
    logic [7:0]   io_exuWriteback_11_bits_robIdx_value;
    logic [4:0]   io_exuWriteback_11_bits_fflags;
    logic         io_exuWriteback_11_bits_wflags;
    logic         io_exuWriteback_10_valid;
    logic [63:0]  io_exuWriteback_10_bits_data_0;
    logic [7:0]   io_exuWriteback_10_bits_robIdx_value;
    logic [4:0]   io_exuWriteback_10_bits_fflags;
    logic         io_exuWriteback_10_bits_wflags;
    logic         io_exuWriteback_9_valid;
    logic [63:0]  io_exuWriteback_9_bits_data_0;
    logic [7:0]   io_exuWriteback_9_bits_robIdx_value;
    logic [4:0]   io_exuWriteback_9_bits_fflags;
    logic         io_exuWriteback_9_bits_wflags;
    logic         io_exuWriteback_8_valid;
    logic [127:0] io_exuWriteback_8_bits_data_0;
    logic [7:0]   io_exuWriteback_8_bits_robIdx_value;
    logic [4:0]   io_exuWriteback_8_bits_fflags;
    logic         io_exuWriteback_8_bits_wflags;
    logic         io_exuWriteback_7_valid;
    logic [63:0]  io_exuWriteback_7_bits_data_0;
    logic [7:0]   io_exuWriteback_7_bits_robIdx_value;
    logic         io_exuWriteback_7_bits_debug_isPerfCnt;
    logic         io_exuWriteback_6_valid;
    logic [63:0]  io_exuWriteback_6_bits_data_0;
    logic [7:0]   io_exuWriteback_6_bits_robIdx_value;
    logic         io_exuWriteback_5_valid;
    logic [127:0] io_exuWriteback_5_bits_data_0;
    logic [7:0]   io_exuWriteback_5_bits_robIdx_value;
    logic         io_exuWriteback_5_bits_redirect_valid;
    logic         io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken;
    logic [4:0]   io_exuWriteback_5_bits_fflags;
    logic         io_exuWriteback_5_bits_wflags;
    logic         io_exuWriteback_4_valid;
    logic [63:0]  io_exuWriteback_4_bits_data_0;
    logic [7:0]   io_exuWriteback_4_bits_robIdx_value;
    logic         io_exuWriteback_3_valid;
    logic [63:0]  io_exuWriteback_3_bits_data_0;
    logic [7:0]   io_exuWriteback_3_bits_robIdx_value;
    logic         io_exuWriteback_3_bits_redirect_valid;
    logic         io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken;
    logic         io_exuWriteback_2_valid;
    logic [63:0]  io_exuWriteback_2_bits_data_0;
    logic [7:0]   io_exuWriteback_2_bits_robIdx_value;
    logic         io_exuWriteback_1_valid;
    logic [63:0]  io_exuWriteback_1_bits_data_0;
    logic [7:0]   io_exuWriteback_1_bits_robIdx_value;
    logic         io_exuWriteback_1_bits_redirect_valid;
    logic         io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken;
    logic         io_exuWriteback_0_valid;
    logic [63:0]  io_exuWriteback_0_bits_data_0;
    logic [7:0]   io_exuWriteback_0_bits_robIdx_value;
    logic [4:0]   io_writebackNums_0_bits;
    logic [4:0]   io_writebackNums_1_bits;
    logic [4:0]   io_writebackNums_2_bits;
    logic [4:0]   io_writebackNums_3_bits;
    logic [4:0]   io_writebackNums_4_bits;
    logic [4:0]   io_writebackNums_5_bits;
    logic [4:0]   io_writebackNums_6_bits;
    logic [4:0]   io_writebackNums_7_bits;
    logic [4:0]   io_writebackNums_8_bits;
    logic [4:0]   io_writebackNums_9_bits;
    logic [4:0]   io_writebackNums_10_bits;
    logic [4:0]   io_writebackNums_11_bits;
    logic [4:0]   io_writebackNums_12_bits;
    logic [4:0]   io_writebackNums_13_bits;
    logic [4:0]   io_writebackNums_14_bits;
    logic [4:0]   io_writebackNums_15_bits;
    logic [4:0]   io_writebackNums_16_bits;
    logic [4:0]   io_writebackNums_17_bits;
    logic [4:0]   io_writebackNums_18_bits;
    logic [4:0]   io_writebackNums_19_bits;
    logic [4:0]   io_writebackNums_20_bits;
    logic [4:0]   io_writebackNums_21_bits;
    logic [4:0]   io_writebackNums_22_bits;
    logic [4:0]   io_writebackNums_23_bits;
    logic [4:0]   io_writebackNums_24_bits;
    logic         io_writebackNeedFlush_0;
    logic         io_writebackNeedFlush_1;
    logic         io_writebackNeedFlush_2;
    logic         io_writebackNeedFlush_6;
    logic         io_writebackNeedFlush_7;
    logic         io_writebackNeedFlush_8;
    logic         io_writebackNeedFlush_9;
    logic         io_writebackNeedFlush_10;
    logic         io_writebackNeedFlush_11;
    logic         io_writebackNeedFlush_12;

    WriteBack_in_agent_xaction  mon_tr;
    while(1) begin
        @this.vif.mon_mp.mon_cb;
        io_writeback_24_valid = this.vif.mon_mp.mon_cb.io_writeback_24_valid;
        io_writeback_24_bits_data_0 = this.vif.mon_mp.mon_cb.io_writeback_24_bits_data_0;
        io_writeback_24_bits_pdest = this.vif.mon_mp.mon_cb.io_writeback_24_bits_pdest;
        io_writeback_24_bits_robIdx_flag = this.vif.mon_mp.mon_cb.io_writeback_24_bits_robIdx_flag;
        io_writeback_24_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_writeback_24_bits_robIdx_value;
        io_writeback_24_bits_vecWen = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vecWen;
        io_writeback_24_bits_v0Wen = this.vif.mon_mp.mon_cb.io_writeback_24_bits_v0Wen;
        io_writeback_24_bits_vlWen = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vlWen;
        io_writeback_24_bits_exceptionVec_0 = this.vif.mon_mp.mon_cb.io_writeback_24_bits_exceptionVec_0;
        io_writeback_24_bits_exceptionVec_1 = this.vif.mon_mp.mon_cb.io_writeback_24_bits_exceptionVec_1;
        io_writeback_24_bits_exceptionVec_2 = this.vif.mon_mp.mon_cb.io_writeback_24_bits_exceptionVec_2;
        io_writeback_24_bits_exceptionVec_3 = this.vif.mon_mp.mon_cb.io_writeback_24_bits_exceptionVec_3;
        io_writeback_24_bits_exceptionVec_4 = this.vif.mon_mp.mon_cb.io_writeback_24_bits_exceptionVec_4;
        io_writeback_24_bits_exceptionVec_5 = this.vif.mon_mp.mon_cb.io_writeback_24_bits_exceptionVec_5;
        io_writeback_24_bits_exceptionVec_6 = this.vif.mon_mp.mon_cb.io_writeback_24_bits_exceptionVec_6;
        io_writeback_24_bits_exceptionVec_7 = this.vif.mon_mp.mon_cb.io_writeback_24_bits_exceptionVec_7;
        io_writeback_24_bits_exceptionVec_8 = this.vif.mon_mp.mon_cb.io_writeback_24_bits_exceptionVec_8;
        io_writeback_24_bits_exceptionVec_9 = this.vif.mon_mp.mon_cb.io_writeback_24_bits_exceptionVec_9;
        io_writeback_24_bits_exceptionVec_10 = this.vif.mon_mp.mon_cb.io_writeback_24_bits_exceptionVec_10;
        io_writeback_24_bits_exceptionVec_11 = this.vif.mon_mp.mon_cb.io_writeback_24_bits_exceptionVec_11;
        io_writeback_24_bits_exceptionVec_12 = this.vif.mon_mp.mon_cb.io_writeback_24_bits_exceptionVec_12;
        io_writeback_24_bits_exceptionVec_13 = this.vif.mon_mp.mon_cb.io_writeback_24_bits_exceptionVec_13;
        io_writeback_24_bits_exceptionVec_14 = this.vif.mon_mp.mon_cb.io_writeback_24_bits_exceptionVec_14;
        io_writeback_24_bits_exceptionVec_15 = this.vif.mon_mp.mon_cb.io_writeback_24_bits_exceptionVec_15;
        io_writeback_24_bits_exceptionVec_16 = this.vif.mon_mp.mon_cb.io_writeback_24_bits_exceptionVec_16;
        io_writeback_24_bits_exceptionVec_17 = this.vif.mon_mp.mon_cb.io_writeback_24_bits_exceptionVec_17;
        io_writeback_24_bits_exceptionVec_18 = this.vif.mon_mp.mon_cb.io_writeback_24_bits_exceptionVec_18;
        io_writeback_24_bits_exceptionVec_19 = this.vif.mon_mp.mon_cb.io_writeback_24_bits_exceptionVec_19;
        io_writeback_24_bits_exceptionVec_20 = this.vif.mon_mp.mon_cb.io_writeback_24_bits_exceptionVec_20;
        io_writeback_24_bits_exceptionVec_21 = this.vif.mon_mp.mon_cb.io_writeback_24_bits_exceptionVec_21;
        io_writeback_24_bits_exceptionVec_22 = this.vif.mon_mp.mon_cb.io_writeback_24_bits_exceptionVec_22;
        io_writeback_24_bits_exceptionVec_23 = this.vif.mon_mp.mon_cb.io_writeback_24_bits_exceptionVec_23;
        io_writeback_24_bits_flushPipe = this.vif.mon_mp.mon_cb.io_writeback_24_bits_flushPipe;
        io_writeback_24_bits_replay = this.vif.mon_mp.mon_cb.io_writeback_24_bits_replay;
        io_writeback_24_bits_trigger = this.vif.mon_mp.mon_cb.io_writeback_24_bits_trigger;
        io_writeback_24_bits_vls_vpu_vill = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_vill;
        io_writeback_24_bits_vls_vpu_vma = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_vma;
        io_writeback_24_bits_vls_vpu_vta = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_vta;
        io_writeback_24_bits_vls_vpu_vsew = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_vsew;
        io_writeback_24_bits_vls_vpu_vlmul = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_vlmul;
        io_writeback_24_bits_vls_vpu_specVill = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_specVill;
        io_writeback_24_bits_vls_vpu_specVma = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_specVma;
        io_writeback_24_bits_vls_vpu_specVta = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_specVta;
        io_writeback_24_bits_vls_vpu_specVsew = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_specVsew;
        io_writeback_24_bits_vls_vpu_specVlmul = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_specVlmul;
        io_writeback_24_bits_vls_vpu_vm = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_vm;
        io_writeback_24_bits_vls_vpu_vstart = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_vstart;
        io_writeback_24_bits_vls_vpu_frm = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_frm;
        io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst;
        io_writeback_24_bits_vls_vpu_fpu_isFP32Instr = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_fpu_isFP32Instr;
        io_writeback_24_bits_vls_vpu_fpu_isFP64Instr = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_fpu_isFP64Instr;
        io_writeback_24_bits_vls_vpu_fpu_isReduction = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_fpu_isReduction;
        io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2 = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2;
        io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4 = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4;
        io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8 = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8;
        io_writeback_24_bits_vls_vpu_vxrm = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_vxrm;
        io_writeback_24_bits_vls_vpu_vuopIdx = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_vuopIdx;
        io_writeback_24_bits_vls_vpu_lastUop = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_lastUop;
        io_writeback_24_bits_vls_vpu_vmask = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_vmask;
        io_writeback_24_bits_vls_vpu_vl = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_vl;
        io_writeback_24_bits_vls_vpu_nf = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_nf;
        io_writeback_24_bits_vls_vpu_veew = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_veew;
        io_writeback_24_bits_vls_vpu_isReverse = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_isReverse;
        io_writeback_24_bits_vls_vpu_isExt = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_isExt;
        io_writeback_24_bits_vls_vpu_isNarrow = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_isNarrow;
        io_writeback_24_bits_vls_vpu_isDstMask = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_isDstMask;
        io_writeback_24_bits_vls_vpu_isOpMask = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_isOpMask;
        io_writeback_24_bits_vls_vpu_isMove = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_isMove;
        io_writeback_24_bits_vls_vpu_isDependOldVd = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_isDependOldVd;
        io_writeback_24_bits_vls_vpu_isWritePartVd = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_isWritePartVd;
        io_writeback_24_bits_vls_vpu_isVleff = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vpu_isVleff;
        io_writeback_24_bits_vls_oldVdPsrc = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_oldVdPsrc;
        io_writeback_24_bits_vls_vdIdx = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vdIdx;
        io_writeback_24_bits_vls_vdIdxInField = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_vdIdxInField;
        io_writeback_24_bits_vls_isIndexed = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_isIndexed;
        io_writeback_24_bits_vls_isMasked = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_isMasked;
        io_writeback_24_bits_vls_isStrided = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_isStrided;
        io_writeback_24_bits_vls_isWhole = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_isWhole;
        io_writeback_24_bits_vls_isVecLoad = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_isVecLoad;
        io_writeback_24_bits_vls_isVlm = this.vif.mon_mp.mon_cb.io_writeback_24_bits_vls_isVlm;
        io_writeback_24_bits_debug_isMMIO = this.vif.mon_mp.mon_cb.io_writeback_24_bits_debug_isMMIO;
        io_writeback_24_bits_debug_isNCIO = this.vif.mon_mp.mon_cb.io_writeback_24_bits_debug_isNCIO;
        io_writeback_24_bits_debug_isPerfCnt = this.vif.mon_mp.mon_cb.io_writeback_24_bits_debug_isPerfCnt;
        io_writeback_24_bits_debug_paddr = this.vif.mon_mp.mon_cb.io_writeback_24_bits_debug_paddr;
        io_writeback_24_bits_debug_vaddr = this.vif.mon_mp.mon_cb.io_writeback_24_bits_debug_vaddr;
        io_writeback_24_bits_debugInfo_eliminatedMove = this.vif.mon_mp.mon_cb.io_writeback_24_bits_debugInfo_eliminatedMove;
        io_writeback_24_bits_debugInfo_renameTime = this.vif.mon_mp.mon_cb.io_writeback_24_bits_debugInfo_renameTime;
        io_writeback_24_bits_debugInfo_dispatchTime = this.vif.mon_mp.mon_cb.io_writeback_24_bits_debugInfo_dispatchTime;
        io_writeback_24_bits_debugInfo_enqRsTime = this.vif.mon_mp.mon_cb.io_writeback_24_bits_debugInfo_enqRsTime;
        io_writeback_24_bits_debugInfo_selectTime = this.vif.mon_mp.mon_cb.io_writeback_24_bits_debugInfo_selectTime;
        io_writeback_24_bits_debugInfo_issueTime = this.vif.mon_mp.mon_cb.io_writeback_24_bits_debugInfo_issueTime;
        io_writeback_24_bits_debugInfo_writebackTime = this.vif.mon_mp.mon_cb.io_writeback_24_bits_debugInfo_writebackTime;
        io_writeback_24_bits_debugInfo_runahead_checkpoint_id = this.vif.mon_mp.mon_cb.io_writeback_24_bits_debugInfo_runahead_checkpoint_id;
        io_writeback_24_bits_debugInfo_tlbFirstReqTime = this.vif.mon_mp.mon_cb.io_writeback_24_bits_debugInfo_tlbFirstReqTime;
        io_writeback_24_bits_debugInfo_tlbRespTime = this.vif.mon_mp.mon_cb.io_writeback_24_bits_debugInfo_tlbRespTime;
        io_writeback_24_bits_debug_seqNum = this.vif.mon_mp.mon_cb.io_writeback_24_bits_debug_seqNum;
        io_writeback_23_valid = this.vif.mon_mp.mon_cb.io_writeback_23_valid;
        io_writeback_23_bits_data_0 = this.vif.mon_mp.mon_cb.io_writeback_23_bits_data_0;
        io_writeback_23_bits_pdest = this.vif.mon_mp.mon_cb.io_writeback_23_bits_pdest;
        io_writeback_23_bits_robIdx_flag = this.vif.mon_mp.mon_cb.io_writeback_23_bits_robIdx_flag;
        io_writeback_23_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_writeback_23_bits_robIdx_value;
        io_writeback_23_bits_vecWen = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vecWen;
        io_writeback_23_bits_v0Wen = this.vif.mon_mp.mon_cb.io_writeback_23_bits_v0Wen;
        io_writeback_23_bits_vlWen = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vlWen;
        io_writeback_23_bits_exceptionVec_0 = this.vif.mon_mp.mon_cb.io_writeback_23_bits_exceptionVec_0;
        io_writeback_23_bits_exceptionVec_1 = this.vif.mon_mp.mon_cb.io_writeback_23_bits_exceptionVec_1;
        io_writeback_23_bits_exceptionVec_2 = this.vif.mon_mp.mon_cb.io_writeback_23_bits_exceptionVec_2;
        io_writeback_23_bits_exceptionVec_3 = this.vif.mon_mp.mon_cb.io_writeback_23_bits_exceptionVec_3;
        io_writeback_23_bits_exceptionVec_4 = this.vif.mon_mp.mon_cb.io_writeback_23_bits_exceptionVec_4;
        io_writeback_23_bits_exceptionVec_5 = this.vif.mon_mp.mon_cb.io_writeback_23_bits_exceptionVec_5;
        io_writeback_23_bits_exceptionVec_6 = this.vif.mon_mp.mon_cb.io_writeback_23_bits_exceptionVec_6;
        io_writeback_23_bits_exceptionVec_7 = this.vif.mon_mp.mon_cb.io_writeback_23_bits_exceptionVec_7;
        io_writeback_23_bits_exceptionVec_8 = this.vif.mon_mp.mon_cb.io_writeback_23_bits_exceptionVec_8;
        io_writeback_23_bits_exceptionVec_9 = this.vif.mon_mp.mon_cb.io_writeback_23_bits_exceptionVec_9;
        io_writeback_23_bits_exceptionVec_10 = this.vif.mon_mp.mon_cb.io_writeback_23_bits_exceptionVec_10;
        io_writeback_23_bits_exceptionVec_11 = this.vif.mon_mp.mon_cb.io_writeback_23_bits_exceptionVec_11;
        io_writeback_23_bits_exceptionVec_12 = this.vif.mon_mp.mon_cb.io_writeback_23_bits_exceptionVec_12;
        io_writeback_23_bits_exceptionVec_13 = this.vif.mon_mp.mon_cb.io_writeback_23_bits_exceptionVec_13;
        io_writeback_23_bits_exceptionVec_14 = this.vif.mon_mp.mon_cb.io_writeback_23_bits_exceptionVec_14;
        io_writeback_23_bits_exceptionVec_15 = this.vif.mon_mp.mon_cb.io_writeback_23_bits_exceptionVec_15;
        io_writeback_23_bits_exceptionVec_16 = this.vif.mon_mp.mon_cb.io_writeback_23_bits_exceptionVec_16;
        io_writeback_23_bits_exceptionVec_17 = this.vif.mon_mp.mon_cb.io_writeback_23_bits_exceptionVec_17;
        io_writeback_23_bits_exceptionVec_18 = this.vif.mon_mp.mon_cb.io_writeback_23_bits_exceptionVec_18;
        io_writeback_23_bits_exceptionVec_19 = this.vif.mon_mp.mon_cb.io_writeback_23_bits_exceptionVec_19;
        io_writeback_23_bits_exceptionVec_20 = this.vif.mon_mp.mon_cb.io_writeback_23_bits_exceptionVec_20;
        io_writeback_23_bits_exceptionVec_21 = this.vif.mon_mp.mon_cb.io_writeback_23_bits_exceptionVec_21;
        io_writeback_23_bits_exceptionVec_22 = this.vif.mon_mp.mon_cb.io_writeback_23_bits_exceptionVec_22;
        io_writeback_23_bits_exceptionVec_23 = this.vif.mon_mp.mon_cb.io_writeback_23_bits_exceptionVec_23;
        io_writeback_23_bits_flushPipe = this.vif.mon_mp.mon_cb.io_writeback_23_bits_flushPipe;
        io_writeback_23_bits_replay = this.vif.mon_mp.mon_cb.io_writeback_23_bits_replay;
        io_writeback_23_bits_trigger = this.vif.mon_mp.mon_cb.io_writeback_23_bits_trigger;
        io_writeback_23_bits_vls_vpu_vill = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_vill;
        io_writeback_23_bits_vls_vpu_vma = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_vma;
        io_writeback_23_bits_vls_vpu_vta = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_vta;
        io_writeback_23_bits_vls_vpu_vsew = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_vsew;
        io_writeback_23_bits_vls_vpu_vlmul = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_vlmul;
        io_writeback_23_bits_vls_vpu_specVill = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_specVill;
        io_writeback_23_bits_vls_vpu_specVma = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_specVma;
        io_writeback_23_bits_vls_vpu_specVta = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_specVta;
        io_writeback_23_bits_vls_vpu_specVsew = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_specVsew;
        io_writeback_23_bits_vls_vpu_specVlmul = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_specVlmul;
        io_writeback_23_bits_vls_vpu_vm = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_vm;
        io_writeback_23_bits_vls_vpu_vstart = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_vstart;
        io_writeback_23_bits_vls_vpu_frm = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_frm;
        io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst;
        io_writeback_23_bits_vls_vpu_fpu_isFP32Instr = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_fpu_isFP32Instr;
        io_writeback_23_bits_vls_vpu_fpu_isFP64Instr = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_fpu_isFP64Instr;
        io_writeback_23_bits_vls_vpu_fpu_isReduction = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_fpu_isReduction;
        io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2 = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2;
        io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4 = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4;
        io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8 = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8;
        io_writeback_23_bits_vls_vpu_vxrm = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_vxrm;
        io_writeback_23_bits_vls_vpu_vuopIdx = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_vuopIdx;
        io_writeback_23_bits_vls_vpu_lastUop = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_lastUop;
        io_writeback_23_bits_vls_vpu_vmask = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_vmask;
        io_writeback_23_bits_vls_vpu_vl = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_vl;
        io_writeback_23_bits_vls_vpu_nf = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_nf;
        io_writeback_23_bits_vls_vpu_veew = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_veew;
        io_writeback_23_bits_vls_vpu_isReverse = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_isReverse;
        io_writeback_23_bits_vls_vpu_isExt = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_isExt;
        io_writeback_23_bits_vls_vpu_isNarrow = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_isNarrow;
        io_writeback_23_bits_vls_vpu_isDstMask = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_isDstMask;
        io_writeback_23_bits_vls_vpu_isOpMask = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_isOpMask;
        io_writeback_23_bits_vls_vpu_isMove = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_isMove;
        io_writeback_23_bits_vls_vpu_isDependOldVd = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_isDependOldVd;
        io_writeback_23_bits_vls_vpu_isWritePartVd = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_isWritePartVd;
        io_writeback_23_bits_vls_vpu_isVleff = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vpu_isVleff;
        io_writeback_23_bits_vls_oldVdPsrc = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_oldVdPsrc;
        io_writeback_23_bits_vls_vdIdx = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vdIdx;
        io_writeback_23_bits_vls_vdIdxInField = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_vdIdxInField;
        io_writeback_23_bits_vls_isIndexed = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_isIndexed;
        io_writeback_23_bits_vls_isMasked = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_isMasked;
        io_writeback_23_bits_vls_isStrided = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_isStrided;
        io_writeback_23_bits_vls_isWhole = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_isWhole;
        io_writeback_23_bits_vls_isVecLoad = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_isVecLoad;
        io_writeback_23_bits_vls_isVlm = this.vif.mon_mp.mon_cb.io_writeback_23_bits_vls_isVlm;
        io_writeback_23_bits_debug_isMMIO = this.vif.mon_mp.mon_cb.io_writeback_23_bits_debug_isMMIO;
        io_writeback_23_bits_debug_isNCIO = this.vif.mon_mp.mon_cb.io_writeback_23_bits_debug_isNCIO;
        io_writeback_23_bits_debug_isPerfCnt = this.vif.mon_mp.mon_cb.io_writeback_23_bits_debug_isPerfCnt;
        io_writeback_23_bits_debug_paddr = this.vif.mon_mp.mon_cb.io_writeback_23_bits_debug_paddr;
        io_writeback_23_bits_debug_vaddr = this.vif.mon_mp.mon_cb.io_writeback_23_bits_debug_vaddr;
        io_writeback_23_bits_debugInfo_eliminatedMove = this.vif.mon_mp.mon_cb.io_writeback_23_bits_debugInfo_eliminatedMove;
        io_writeback_23_bits_debugInfo_renameTime = this.vif.mon_mp.mon_cb.io_writeback_23_bits_debugInfo_renameTime;
        io_writeback_23_bits_debugInfo_dispatchTime = this.vif.mon_mp.mon_cb.io_writeback_23_bits_debugInfo_dispatchTime;
        io_writeback_23_bits_debugInfo_enqRsTime = this.vif.mon_mp.mon_cb.io_writeback_23_bits_debugInfo_enqRsTime;
        io_writeback_23_bits_debugInfo_selectTime = this.vif.mon_mp.mon_cb.io_writeback_23_bits_debugInfo_selectTime;
        io_writeback_23_bits_debugInfo_issueTime = this.vif.mon_mp.mon_cb.io_writeback_23_bits_debugInfo_issueTime;
        io_writeback_23_bits_debugInfo_writebackTime = this.vif.mon_mp.mon_cb.io_writeback_23_bits_debugInfo_writebackTime;
        io_writeback_23_bits_debugInfo_runahead_checkpoint_id = this.vif.mon_mp.mon_cb.io_writeback_23_bits_debugInfo_runahead_checkpoint_id;
        io_writeback_23_bits_debugInfo_tlbFirstReqTime = this.vif.mon_mp.mon_cb.io_writeback_23_bits_debugInfo_tlbFirstReqTime;
        io_writeback_23_bits_debugInfo_tlbRespTime = this.vif.mon_mp.mon_cb.io_writeback_23_bits_debugInfo_tlbRespTime;
        io_writeback_23_bits_debug_seqNum = this.vif.mon_mp.mon_cb.io_writeback_23_bits_debug_seqNum;
        io_writeback_22_valid = this.vif.mon_mp.mon_cb.io_writeback_22_valid;
        io_writeback_22_bits_data_0 = this.vif.mon_mp.mon_cb.io_writeback_22_bits_data_0;
        io_writeback_22_bits_pdest = this.vif.mon_mp.mon_cb.io_writeback_22_bits_pdest;
        io_writeback_22_bits_robIdx_flag = this.vif.mon_mp.mon_cb.io_writeback_22_bits_robIdx_flag;
        io_writeback_22_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_writeback_22_bits_robIdx_value;
        io_writeback_22_bits_intWen = this.vif.mon_mp.mon_cb.io_writeback_22_bits_intWen;
        io_writeback_22_bits_fpWen = this.vif.mon_mp.mon_cb.io_writeback_22_bits_fpWen;
        io_writeback_22_bits_exceptionVec_0 = this.vif.mon_mp.mon_cb.io_writeback_22_bits_exceptionVec_0;
        io_writeback_22_bits_exceptionVec_1 = this.vif.mon_mp.mon_cb.io_writeback_22_bits_exceptionVec_1;
        io_writeback_22_bits_exceptionVec_2 = this.vif.mon_mp.mon_cb.io_writeback_22_bits_exceptionVec_2;
        io_writeback_22_bits_exceptionVec_3 = this.vif.mon_mp.mon_cb.io_writeback_22_bits_exceptionVec_3;
        io_writeback_22_bits_exceptionVec_4 = this.vif.mon_mp.mon_cb.io_writeback_22_bits_exceptionVec_4;
        io_writeback_22_bits_exceptionVec_5 = this.vif.mon_mp.mon_cb.io_writeback_22_bits_exceptionVec_5;
        io_writeback_22_bits_exceptionVec_6 = this.vif.mon_mp.mon_cb.io_writeback_22_bits_exceptionVec_6;
        io_writeback_22_bits_exceptionVec_7 = this.vif.mon_mp.mon_cb.io_writeback_22_bits_exceptionVec_7;
        io_writeback_22_bits_exceptionVec_8 = this.vif.mon_mp.mon_cb.io_writeback_22_bits_exceptionVec_8;
        io_writeback_22_bits_exceptionVec_9 = this.vif.mon_mp.mon_cb.io_writeback_22_bits_exceptionVec_9;
        io_writeback_22_bits_exceptionVec_10 = this.vif.mon_mp.mon_cb.io_writeback_22_bits_exceptionVec_10;
        io_writeback_22_bits_exceptionVec_11 = this.vif.mon_mp.mon_cb.io_writeback_22_bits_exceptionVec_11;
        io_writeback_22_bits_exceptionVec_12 = this.vif.mon_mp.mon_cb.io_writeback_22_bits_exceptionVec_12;
        io_writeback_22_bits_exceptionVec_13 = this.vif.mon_mp.mon_cb.io_writeback_22_bits_exceptionVec_13;
        io_writeback_22_bits_exceptionVec_14 = this.vif.mon_mp.mon_cb.io_writeback_22_bits_exceptionVec_14;
        io_writeback_22_bits_exceptionVec_15 = this.vif.mon_mp.mon_cb.io_writeback_22_bits_exceptionVec_15;
        io_writeback_22_bits_exceptionVec_16 = this.vif.mon_mp.mon_cb.io_writeback_22_bits_exceptionVec_16;
        io_writeback_22_bits_exceptionVec_17 = this.vif.mon_mp.mon_cb.io_writeback_22_bits_exceptionVec_17;
        io_writeback_22_bits_exceptionVec_18 = this.vif.mon_mp.mon_cb.io_writeback_22_bits_exceptionVec_18;
        io_writeback_22_bits_exceptionVec_19 = this.vif.mon_mp.mon_cb.io_writeback_22_bits_exceptionVec_19;
        io_writeback_22_bits_exceptionVec_20 = this.vif.mon_mp.mon_cb.io_writeback_22_bits_exceptionVec_20;
        io_writeback_22_bits_exceptionVec_21 = this.vif.mon_mp.mon_cb.io_writeback_22_bits_exceptionVec_21;
        io_writeback_22_bits_exceptionVec_22 = this.vif.mon_mp.mon_cb.io_writeback_22_bits_exceptionVec_22;
        io_writeback_22_bits_exceptionVec_23 = this.vif.mon_mp.mon_cb.io_writeback_22_bits_exceptionVec_23;
        io_writeback_22_bits_flushPipe = this.vif.mon_mp.mon_cb.io_writeback_22_bits_flushPipe;
        io_writeback_22_bits_replay = this.vif.mon_mp.mon_cb.io_writeback_22_bits_replay;
        io_writeback_22_bits_lqIdx_flag = this.vif.mon_mp.mon_cb.io_writeback_22_bits_lqIdx_flag;
        io_writeback_22_bits_lqIdx_value = this.vif.mon_mp.mon_cb.io_writeback_22_bits_lqIdx_value;
        io_writeback_22_bits_trigger = this.vif.mon_mp.mon_cb.io_writeback_22_bits_trigger;
        io_writeback_22_bits_predecodeInfo_valid = this.vif.mon_mp.mon_cb.io_writeback_22_bits_predecodeInfo_valid;
        io_writeback_22_bits_predecodeInfo_isRVC = this.vif.mon_mp.mon_cb.io_writeback_22_bits_predecodeInfo_isRVC;
        io_writeback_22_bits_predecodeInfo_brType = this.vif.mon_mp.mon_cb.io_writeback_22_bits_predecodeInfo_brType;
        io_writeback_22_bits_predecodeInfo_isCall = this.vif.mon_mp.mon_cb.io_writeback_22_bits_predecodeInfo_isCall;
        io_writeback_22_bits_predecodeInfo_isRet = this.vif.mon_mp.mon_cb.io_writeback_22_bits_predecodeInfo_isRet;
        io_writeback_22_bits_debug_isMMIO = this.vif.mon_mp.mon_cb.io_writeback_22_bits_debug_isMMIO;
        io_writeback_22_bits_debug_isNCIO = this.vif.mon_mp.mon_cb.io_writeback_22_bits_debug_isNCIO;
        io_writeback_22_bits_debug_isPerfCnt = this.vif.mon_mp.mon_cb.io_writeback_22_bits_debug_isPerfCnt;
        io_writeback_22_bits_debug_paddr = this.vif.mon_mp.mon_cb.io_writeback_22_bits_debug_paddr;
        io_writeback_22_bits_debug_vaddr = this.vif.mon_mp.mon_cb.io_writeback_22_bits_debug_vaddr;
        io_writeback_22_bits_debugInfo_eliminatedMove = this.vif.mon_mp.mon_cb.io_writeback_22_bits_debugInfo_eliminatedMove;
        io_writeback_22_bits_debugInfo_renameTime = this.vif.mon_mp.mon_cb.io_writeback_22_bits_debugInfo_renameTime;
        io_writeback_22_bits_debugInfo_dispatchTime = this.vif.mon_mp.mon_cb.io_writeback_22_bits_debugInfo_dispatchTime;
        io_writeback_22_bits_debugInfo_enqRsTime = this.vif.mon_mp.mon_cb.io_writeback_22_bits_debugInfo_enqRsTime;
        io_writeback_22_bits_debugInfo_selectTime = this.vif.mon_mp.mon_cb.io_writeback_22_bits_debugInfo_selectTime;
        io_writeback_22_bits_debugInfo_issueTime = this.vif.mon_mp.mon_cb.io_writeback_22_bits_debugInfo_issueTime;
        io_writeback_22_bits_debugInfo_writebackTime = this.vif.mon_mp.mon_cb.io_writeback_22_bits_debugInfo_writebackTime;
        io_writeback_22_bits_debugInfo_runahead_checkpoint_id = this.vif.mon_mp.mon_cb.io_writeback_22_bits_debugInfo_runahead_checkpoint_id;
        io_writeback_22_bits_debugInfo_tlbFirstReqTime = this.vif.mon_mp.mon_cb.io_writeback_22_bits_debugInfo_tlbFirstReqTime;
        io_writeback_22_bits_debugInfo_tlbRespTime = this.vif.mon_mp.mon_cb.io_writeback_22_bits_debugInfo_tlbRespTime;
        io_writeback_22_bits_debug_seqNum = this.vif.mon_mp.mon_cb.io_writeback_22_bits_debug_seqNum;
        io_writeback_21_valid = this.vif.mon_mp.mon_cb.io_writeback_21_valid;
        io_writeback_21_bits_data_0 = this.vif.mon_mp.mon_cb.io_writeback_21_bits_data_0;
        io_writeback_21_bits_pdest = this.vif.mon_mp.mon_cb.io_writeback_21_bits_pdest;
        io_writeback_21_bits_robIdx_flag = this.vif.mon_mp.mon_cb.io_writeback_21_bits_robIdx_flag;
        io_writeback_21_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_writeback_21_bits_robIdx_value;
        io_writeback_21_bits_intWen = this.vif.mon_mp.mon_cb.io_writeback_21_bits_intWen;
        io_writeback_21_bits_fpWen = this.vif.mon_mp.mon_cb.io_writeback_21_bits_fpWen;
        io_writeback_21_bits_exceptionVec_0 = this.vif.mon_mp.mon_cb.io_writeback_21_bits_exceptionVec_0;
        io_writeback_21_bits_exceptionVec_1 = this.vif.mon_mp.mon_cb.io_writeback_21_bits_exceptionVec_1;
        io_writeback_21_bits_exceptionVec_2 = this.vif.mon_mp.mon_cb.io_writeback_21_bits_exceptionVec_2;
        io_writeback_21_bits_exceptionVec_3 = this.vif.mon_mp.mon_cb.io_writeback_21_bits_exceptionVec_3;
        io_writeback_21_bits_exceptionVec_4 = this.vif.mon_mp.mon_cb.io_writeback_21_bits_exceptionVec_4;
        io_writeback_21_bits_exceptionVec_5 = this.vif.mon_mp.mon_cb.io_writeback_21_bits_exceptionVec_5;
        io_writeback_21_bits_exceptionVec_6 = this.vif.mon_mp.mon_cb.io_writeback_21_bits_exceptionVec_6;
        io_writeback_21_bits_exceptionVec_7 = this.vif.mon_mp.mon_cb.io_writeback_21_bits_exceptionVec_7;
        io_writeback_21_bits_exceptionVec_8 = this.vif.mon_mp.mon_cb.io_writeback_21_bits_exceptionVec_8;
        io_writeback_21_bits_exceptionVec_9 = this.vif.mon_mp.mon_cb.io_writeback_21_bits_exceptionVec_9;
        io_writeback_21_bits_exceptionVec_10 = this.vif.mon_mp.mon_cb.io_writeback_21_bits_exceptionVec_10;
        io_writeback_21_bits_exceptionVec_11 = this.vif.mon_mp.mon_cb.io_writeback_21_bits_exceptionVec_11;
        io_writeback_21_bits_exceptionVec_12 = this.vif.mon_mp.mon_cb.io_writeback_21_bits_exceptionVec_12;
        io_writeback_21_bits_exceptionVec_13 = this.vif.mon_mp.mon_cb.io_writeback_21_bits_exceptionVec_13;
        io_writeback_21_bits_exceptionVec_14 = this.vif.mon_mp.mon_cb.io_writeback_21_bits_exceptionVec_14;
        io_writeback_21_bits_exceptionVec_15 = this.vif.mon_mp.mon_cb.io_writeback_21_bits_exceptionVec_15;
        io_writeback_21_bits_exceptionVec_16 = this.vif.mon_mp.mon_cb.io_writeback_21_bits_exceptionVec_16;
        io_writeback_21_bits_exceptionVec_17 = this.vif.mon_mp.mon_cb.io_writeback_21_bits_exceptionVec_17;
        io_writeback_21_bits_exceptionVec_18 = this.vif.mon_mp.mon_cb.io_writeback_21_bits_exceptionVec_18;
        io_writeback_21_bits_exceptionVec_19 = this.vif.mon_mp.mon_cb.io_writeback_21_bits_exceptionVec_19;
        io_writeback_21_bits_exceptionVec_20 = this.vif.mon_mp.mon_cb.io_writeback_21_bits_exceptionVec_20;
        io_writeback_21_bits_exceptionVec_21 = this.vif.mon_mp.mon_cb.io_writeback_21_bits_exceptionVec_21;
        io_writeback_21_bits_exceptionVec_22 = this.vif.mon_mp.mon_cb.io_writeback_21_bits_exceptionVec_22;
        io_writeback_21_bits_exceptionVec_23 = this.vif.mon_mp.mon_cb.io_writeback_21_bits_exceptionVec_23;
        io_writeback_21_bits_flushPipe = this.vif.mon_mp.mon_cb.io_writeback_21_bits_flushPipe;
        io_writeback_21_bits_replay = this.vif.mon_mp.mon_cb.io_writeback_21_bits_replay;
        io_writeback_21_bits_lqIdx_flag = this.vif.mon_mp.mon_cb.io_writeback_21_bits_lqIdx_flag;
        io_writeback_21_bits_lqIdx_value = this.vif.mon_mp.mon_cb.io_writeback_21_bits_lqIdx_value;
        io_writeback_21_bits_trigger = this.vif.mon_mp.mon_cb.io_writeback_21_bits_trigger;
        io_writeback_21_bits_predecodeInfo_valid = this.vif.mon_mp.mon_cb.io_writeback_21_bits_predecodeInfo_valid;
        io_writeback_21_bits_predecodeInfo_isRVC = this.vif.mon_mp.mon_cb.io_writeback_21_bits_predecodeInfo_isRVC;
        io_writeback_21_bits_predecodeInfo_brType = this.vif.mon_mp.mon_cb.io_writeback_21_bits_predecodeInfo_brType;
        io_writeback_21_bits_predecodeInfo_isCall = this.vif.mon_mp.mon_cb.io_writeback_21_bits_predecodeInfo_isCall;
        io_writeback_21_bits_predecodeInfo_isRet = this.vif.mon_mp.mon_cb.io_writeback_21_bits_predecodeInfo_isRet;
        io_writeback_21_bits_debug_isMMIO = this.vif.mon_mp.mon_cb.io_writeback_21_bits_debug_isMMIO;
        io_writeback_21_bits_debug_isNCIO = this.vif.mon_mp.mon_cb.io_writeback_21_bits_debug_isNCIO;
        io_writeback_21_bits_debug_isPerfCnt = this.vif.mon_mp.mon_cb.io_writeback_21_bits_debug_isPerfCnt;
        io_writeback_21_bits_debug_paddr = this.vif.mon_mp.mon_cb.io_writeback_21_bits_debug_paddr;
        io_writeback_21_bits_debug_vaddr = this.vif.mon_mp.mon_cb.io_writeback_21_bits_debug_vaddr;
        io_writeback_21_bits_debugInfo_eliminatedMove = this.vif.mon_mp.mon_cb.io_writeback_21_bits_debugInfo_eliminatedMove;
        io_writeback_21_bits_debugInfo_renameTime = this.vif.mon_mp.mon_cb.io_writeback_21_bits_debugInfo_renameTime;
        io_writeback_21_bits_debugInfo_dispatchTime = this.vif.mon_mp.mon_cb.io_writeback_21_bits_debugInfo_dispatchTime;
        io_writeback_21_bits_debugInfo_enqRsTime = this.vif.mon_mp.mon_cb.io_writeback_21_bits_debugInfo_enqRsTime;
        io_writeback_21_bits_debugInfo_selectTime = this.vif.mon_mp.mon_cb.io_writeback_21_bits_debugInfo_selectTime;
        io_writeback_21_bits_debugInfo_issueTime = this.vif.mon_mp.mon_cb.io_writeback_21_bits_debugInfo_issueTime;
        io_writeback_21_bits_debugInfo_writebackTime = this.vif.mon_mp.mon_cb.io_writeback_21_bits_debugInfo_writebackTime;
        io_writeback_21_bits_debugInfo_runahead_checkpoint_id = this.vif.mon_mp.mon_cb.io_writeback_21_bits_debugInfo_runahead_checkpoint_id;
        io_writeback_21_bits_debugInfo_tlbFirstReqTime = this.vif.mon_mp.mon_cb.io_writeback_21_bits_debugInfo_tlbFirstReqTime;
        io_writeback_21_bits_debugInfo_tlbRespTime = this.vif.mon_mp.mon_cb.io_writeback_21_bits_debugInfo_tlbRespTime;
        io_writeback_21_bits_debug_seqNum = this.vif.mon_mp.mon_cb.io_writeback_21_bits_debug_seqNum;
        io_writeback_20_valid = this.vif.mon_mp.mon_cb.io_writeback_20_valid;
        io_writeback_20_bits_data_0 = this.vif.mon_mp.mon_cb.io_writeback_20_bits_data_0;
        io_writeback_20_bits_pdest = this.vif.mon_mp.mon_cb.io_writeback_20_bits_pdest;
        io_writeback_20_bits_robIdx_flag = this.vif.mon_mp.mon_cb.io_writeback_20_bits_robIdx_flag;
        io_writeback_20_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_writeback_20_bits_robIdx_value;
        io_writeback_20_bits_intWen = this.vif.mon_mp.mon_cb.io_writeback_20_bits_intWen;
        io_writeback_20_bits_fpWen = this.vif.mon_mp.mon_cb.io_writeback_20_bits_fpWen;
        io_writeback_20_bits_exceptionVec_0 = this.vif.mon_mp.mon_cb.io_writeback_20_bits_exceptionVec_0;
        io_writeback_20_bits_exceptionVec_1 = this.vif.mon_mp.mon_cb.io_writeback_20_bits_exceptionVec_1;
        io_writeback_20_bits_exceptionVec_2 = this.vif.mon_mp.mon_cb.io_writeback_20_bits_exceptionVec_2;
        io_writeback_20_bits_exceptionVec_3 = this.vif.mon_mp.mon_cb.io_writeback_20_bits_exceptionVec_3;
        io_writeback_20_bits_exceptionVec_4 = this.vif.mon_mp.mon_cb.io_writeback_20_bits_exceptionVec_4;
        io_writeback_20_bits_exceptionVec_5 = this.vif.mon_mp.mon_cb.io_writeback_20_bits_exceptionVec_5;
        io_writeback_20_bits_exceptionVec_6 = this.vif.mon_mp.mon_cb.io_writeback_20_bits_exceptionVec_6;
        io_writeback_20_bits_exceptionVec_7 = this.vif.mon_mp.mon_cb.io_writeback_20_bits_exceptionVec_7;
        io_writeback_20_bits_exceptionVec_8 = this.vif.mon_mp.mon_cb.io_writeback_20_bits_exceptionVec_8;
        io_writeback_20_bits_exceptionVec_9 = this.vif.mon_mp.mon_cb.io_writeback_20_bits_exceptionVec_9;
        io_writeback_20_bits_exceptionVec_10 = this.vif.mon_mp.mon_cb.io_writeback_20_bits_exceptionVec_10;
        io_writeback_20_bits_exceptionVec_11 = this.vif.mon_mp.mon_cb.io_writeback_20_bits_exceptionVec_11;
        io_writeback_20_bits_exceptionVec_12 = this.vif.mon_mp.mon_cb.io_writeback_20_bits_exceptionVec_12;
        io_writeback_20_bits_exceptionVec_13 = this.vif.mon_mp.mon_cb.io_writeback_20_bits_exceptionVec_13;
        io_writeback_20_bits_exceptionVec_14 = this.vif.mon_mp.mon_cb.io_writeback_20_bits_exceptionVec_14;
        io_writeback_20_bits_exceptionVec_15 = this.vif.mon_mp.mon_cb.io_writeback_20_bits_exceptionVec_15;
        io_writeback_20_bits_exceptionVec_16 = this.vif.mon_mp.mon_cb.io_writeback_20_bits_exceptionVec_16;
        io_writeback_20_bits_exceptionVec_17 = this.vif.mon_mp.mon_cb.io_writeback_20_bits_exceptionVec_17;
        io_writeback_20_bits_exceptionVec_18 = this.vif.mon_mp.mon_cb.io_writeback_20_bits_exceptionVec_18;
        io_writeback_20_bits_exceptionVec_19 = this.vif.mon_mp.mon_cb.io_writeback_20_bits_exceptionVec_19;
        io_writeback_20_bits_exceptionVec_20 = this.vif.mon_mp.mon_cb.io_writeback_20_bits_exceptionVec_20;
        io_writeback_20_bits_exceptionVec_21 = this.vif.mon_mp.mon_cb.io_writeback_20_bits_exceptionVec_21;
        io_writeback_20_bits_exceptionVec_22 = this.vif.mon_mp.mon_cb.io_writeback_20_bits_exceptionVec_22;
        io_writeback_20_bits_exceptionVec_23 = this.vif.mon_mp.mon_cb.io_writeback_20_bits_exceptionVec_23;
        io_writeback_20_bits_flushPipe = this.vif.mon_mp.mon_cb.io_writeback_20_bits_flushPipe;
        io_writeback_20_bits_replay = this.vif.mon_mp.mon_cb.io_writeback_20_bits_replay;
        io_writeback_20_bits_lqIdx_flag = this.vif.mon_mp.mon_cb.io_writeback_20_bits_lqIdx_flag;
        io_writeback_20_bits_lqIdx_value = this.vif.mon_mp.mon_cb.io_writeback_20_bits_lqIdx_value;
        io_writeback_20_bits_trigger = this.vif.mon_mp.mon_cb.io_writeback_20_bits_trigger;
        io_writeback_20_bits_predecodeInfo_valid = this.vif.mon_mp.mon_cb.io_writeback_20_bits_predecodeInfo_valid;
        io_writeback_20_bits_predecodeInfo_isRVC = this.vif.mon_mp.mon_cb.io_writeback_20_bits_predecodeInfo_isRVC;
        io_writeback_20_bits_predecodeInfo_brType = this.vif.mon_mp.mon_cb.io_writeback_20_bits_predecodeInfo_brType;
        io_writeback_20_bits_predecodeInfo_isCall = this.vif.mon_mp.mon_cb.io_writeback_20_bits_predecodeInfo_isCall;
        io_writeback_20_bits_predecodeInfo_isRet = this.vif.mon_mp.mon_cb.io_writeback_20_bits_predecodeInfo_isRet;
        io_writeback_20_bits_debug_isMMIO = this.vif.mon_mp.mon_cb.io_writeback_20_bits_debug_isMMIO;
        io_writeback_20_bits_debug_isNCIO = this.vif.mon_mp.mon_cb.io_writeback_20_bits_debug_isNCIO;
        io_writeback_20_bits_debug_isPerfCnt = this.vif.mon_mp.mon_cb.io_writeback_20_bits_debug_isPerfCnt;
        io_writeback_20_bits_debug_paddr = this.vif.mon_mp.mon_cb.io_writeback_20_bits_debug_paddr;
        io_writeback_20_bits_debug_vaddr = this.vif.mon_mp.mon_cb.io_writeback_20_bits_debug_vaddr;
        io_writeback_20_bits_debugInfo_eliminatedMove = this.vif.mon_mp.mon_cb.io_writeback_20_bits_debugInfo_eliminatedMove;
        io_writeback_20_bits_debugInfo_renameTime = this.vif.mon_mp.mon_cb.io_writeback_20_bits_debugInfo_renameTime;
        io_writeback_20_bits_debugInfo_dispatchTime = this.vif.mon_mp.mon_cb.io_writeback_20_bits_debugInfo_dispatchTime;
        io_writeback_20_bits_debugInfo_enqRsTime = this.vif.mon_mp.mon_cb.io_writeback_20_bits_debugInfo_enqRsTime;
        io_writeback_20_bits_debugInfo_selectTime = this.vif.mon_mp.mon_cb.io_writeback_20_bits_debugInfo_selectTime;
        io_writeback_20_bits_debugInfo_issueTime = this.vif.mon_mp.mon_cb.io_writeback_20_bits_debugInfo_issueTime;
        io_writeback_20_bits_debugInfo_writebackTime = this.vif.mon_mp.mon_cb.io_writeback_20_bits_debugInfo_writebackTime;
        io_writeback_20_bits_debugInfo_runahead_checkpoint_id = this.vif.mon_mp.mon_cb.io_writeback_20_bits_debugInfo_runahead_checkpoint_id;
        io_writeback_20_bits_debugInfo_tlbFirstReqTime = this.vif.mon_mp.mon_cb.io_writeback_20_bits_debugInfo_tlbFirstReqTime;
        io_writeback_20_bits_debugInfo_tlbRespTime = this.vif.mon_mp.mon_cb.io_writeback_20_bits_debugInfo_tlbRespTime;
        io_writeback_20_bits_debug_seqNum = this.vif.mon_mp.mon_cb.io_writeback_20_bits_debug_seqNum;
        io_writeback_19_valid = this.vif.mon_mp.mon_cb.io_writeback_19_valid;
        io_writeback_19_bits_data_0 = this.vif.mon_mp.mon_cb.io_writeback_19_bits_data_0;
        io_writeback_19_bits_pdest = this.vif.mon_mp.mon_cb.io_writeback_19_bits_pdest;
        io_writeback_19_bits_robIdx_flag = this.vif.mon_mp.mon_cb.io_writeback_19_bits_robIdx_flag;
        io_writeback_19_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_writeback_19_bits_robIdx_value;
        io_writeback_19_bits_intWen = this.vif.mon_mp.mon_cb.io_writeback_19_bits_intWen;
        io_writeback_19_bits_exceptionVec_0 = this.vif.mon_mp.mon_cb.io_writeback_19_bits_exceptionVec_0;
        io_writeback_19_bits_exceptionVec_1 = this.vif.mon_mp.mon_cb.io_writeback_19_bits_exceptionVec_1;
        io_writeback_19_bits_exceptionVec_2 = this.vif.mon_mp.mon_cb.io_writeback_19_bits_exceptionVec_2;
        io_writeback_19_bits_exceptionVec_3 = this.vif.mon_mp.mon_cb.io_writeback_19_bits_exceptionVec_3;
        io_writeback_19_bits_exceptionVec_4 = this.vif.mon_mp.mon_cb.io_writeback_19_bits_exceptionVec_4;
        io_writeback_19_bits_exceptionVec_5 = this.vif.mon_mp.mon_cb.io_writeback_19_bits_exceptionVec_5;
        io_writeback_19_bits_exceptionVec_6 = this.vif.mon_mp.mon_cb.io_writeback_19_bits_exceptionVec_6;
        io_writeback_19_bits_exceptionVec_7 = this.vif.mon_mp.mon_cb.io_writeback_19_bits_exceptionVec_7;
        io_writeback_19_bits_exceptionVec_8 = this.vif.mon_mp.mon_cb.io_writeback_19_bits_exceptionVec_8;
        io_writeback_19_bits_exceptionVec_9 = this.vif.mon_mp.mon_cb.io_writeback_19_bits_exceptionVec_9;
        io_writeback_19_bits_exceptionVec_10 = this.vif.mon_mp.mon_cb.io_writeback_19_bits_exceptionVec_10;
        io_writeback_19_bits_exceptionVec_11 = this.vif.mon_mp.mon_cb.io_writeback_19_bits_exceptionVec_11;
        io_writeback_19_bits_exceptionVec_12 = this.vif.mon_mp.mon_cb.io_writeback_19_bits_exceptionVec_12;
        io_writeback_19_bits_exceptionVec_13 = this.vif.mon_mp.mon_cb.io_writeback_19_bits_exceptionVec_13;
        io_writeback_19_bits_exceptionVec_14 = this.vif.mon_mp.mon_cb.io_writeback_19_bits_exceptionVec_14;
        io_writeback_19_bits_exceptionVec_15 = this.vif.mon_mp.mon_cb.io_writeback_19_bits_exceptionVec_15;
        io_writeback_19_bits_exceptionVec_16 = this.vif.mon_mp.mon_cb.io_writeback_19_bits_exceptionVec_16;
        io_writeback_19_bits_exceptionVec_17 = this.vif.mon_mp.mon_cb.io_writeback_19_bits_exceptionVec_17;
        io_writeback_19_bits_exceptionVec_18 = this.vif.mon_mp.mon_cb.io_writeback_19_bits_exceptionVec_18;
        io_writeback_19_bits_exceptionVec_19 = this.vif.mon_mp.mon_cb.io_writeback_19_bits_exceptionVec_19;
        io_writeback_19_bits_exceptionVec_20 = this.vif.mon_mp.mon_cb.io_writeback_19_bits_exceptionVec_20;
        io_writeback_19_bits_exceptionVec_21 = this.vif.mon_mp.mon_cb.io_writeback_19_bits_exceptionVec_21;
        io_writeback_19_bits_exceptionVec_22 = this.vif.mon_mp.mon_cb.io_writeback_19_bits_exceptionVec_22;
        io_writeback_19_bits_exceptionVec_23 = this.vif.mon_mp.mon_cb.io_writeback_19_bits_exceptionVec_23;
        io_writeback_19_bits_flushPipe = this.vif.mon_mp.mon_cb.io_writeback_19_bits_flushPipe;
        io_writeback_19_bits_sqIdx_flag = this.vif.mon_mp.mon_cb.io_writeback_19_bits_sqIdx_flag;
        io_writeback_19_bits_sqIdx_value = this.vif.mon_mp.mon_cb.io_writeback_19_bits_sqIdx_value;
        io_writeback_19_bits_trigger = this.vif.mon_mp.mon_cb.io_writeback_19_bits_trigger;
        io_writeback_19_bits_debug_isMMIO = this.vif.mon_mp.mon_cb.io_writeback_19_bits_debug_isMMIO;
        io_writeback_19_bits_debug_isNCIO = this.vif.mon_mp.mon_cb.io_writeback_19_bits_debug_isNCIO;
        io_writeback_19_bits_debug_isPerfCnt = this.vif.mon_mp.mon_cb.io_writeback_19_bits_debug_isPerfCnt;
        io_writeback_19_bits_debug_paddr = this.vif.mon_mp.mon_cb.io_writeback_19_bits_debug_paddr;
        io_writeback_19_bits_debug_vaddr = this.vif.mon_mp.mon_cb.io_writeback_19_bits_debug_vaddr;
        io_writeback_19_bits_debugInfo_eliminatedMove = this.vif.mon_mp.mon_cb.io_writeback_19_bits_debugInfo_eliminatedMove;
        io_writeback_19_bits_debugInfo_renameTime = this.vif.mon_mp.mon_cb.io_writeback_19_bits_debugInfo_renameTime;
        io_writeback_19_bits_debugInfo_dispatchTime = this.vif.mon_mp.mon_cb.io_writeback_19_bits_debugInfo_dispatchTime;
        io_writeback_19_bits_debugInfo_enqRsTime = this.vif.mon_mp.mon_cb.io_writeback_19_bits_debugInfo_enqRsTime;
        io_writeback_19_bits_debugInfo_selectTime = this.vif.mon_mp.mon_cb.io_writeback_19_bits_debugInfo_selectTime;
        io_writeback_19_bits_debugInfo_issueTime = this.vif.mon_mp.mon_cb.io_writeback_19_bits_debugInfo_issueTime;
        io_writeback_19_bits_debugInfo_writebackTime = this.vif.mon_mp.mon_cb.io_writeback_19_bits_debugInfo_writebackTime;
        io_writeback_19_bits_debugInfo_runahead_checkpoint_id = this.vif.mon_mp.mon_cb.io_writeback_19_bits_debugInfo_runahead_checkpoint_id;
        io_writeback_19_bits_debugInfo_tlbFirstReqTime = this.vif.mon_mp.mon_cb.io_writeback_19_bits_debugInfo_tlbFirstReqTime;
        io_writeback_19_bits_debugInfo_tlbRespTime = this.vif.mon_mp.mon_cb.io_writeback_19_bits_debugInfo_tlbRespTime;
        io_writeback_19_bits_debug_seqNum = this.vif.mon_mp.mon_cb.io_writeback_19_bits_debug_seqNum;
        io_writeback_18_valid = this.vif.mon_mp.mon_cb.io_writeback_18_valid;
        io_writeback_18_bits_data_0 = this.vif.mon_mp.mon_cb.io_writeback_18_bits_data_0;
        io_writeback_18_bits_pdest = this.vif.mon_mp.mon_cb.io_writeback_18_bits_pdest;
        io_writeback_18_bits_robIdx_flag = this.vif.mon_mp.mon_cb.io_writeback_18_bits_robIdx_flag;
        io_writeback_18_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_writeback_18_bits_robIdx_value;
        io_writeback_18_bits_intWen = this.vif.mon_mp.mon_cb.io_writeback_18_bits_intWen;
        io_writeback_18_bits_exceptionVec_0 = this.vif.mon_mp.mon_cb.io_writeback_18_bits_exceptionVec_0;
        io_writeback_18_bits_exceptionVec_1 = this.vif.mon_mp.mon_cb.io_writeback_18_bits_exceptionVec_1;
        io_writeback_18_bits_exceptionVec_2 = this.vif.mon_mp.mon_cb.io_writeback_18_bits_exceptionVec_2;
        io_writeback_18_bits_exceptionVec_3 = this.vif.mon_mp.mon_cb.io_writeback_18_bits_exceptionVec_3;
        io_writeback_18_bits_exceptionVec_4 = this.vif.mon_mp.mon_cb.io_writeback_18_bits_exceptionVec_4;
        io_writeback_18_bits_exceptionVec_5 = this.vif.mon_mp.mon_cb.io_writeback_18_bits_exceptionVec_5;
        io_writeback_18_bits_exceptionVec_6 = this.vif.mon_mp.mon_cb.io_writeback_18_bits_exceptionVec_6;
        io_writeback_18_bits_exceptionVec_7 = this.vif.mon_mp.mon_cb.io_writeback_18_bits_exceptionVec_7;
        io_writeback_18_bits_exceptionVec_8 = this.vif.mon_mp.mon_cb.io_writeback_18_bits_exceptionVec_8;
        io_writeback_18_bits_exceptionVec_9 = this.vif.mon_mp.mon_cb.io_writeback_18_bits_exceptionVec_9;
        io_writeback_18_bits_exceptionVec_10 = this.vif.mon_mp.mon_cb.io_writeback_18_bits_exceptionVec_10;
        io_writeback_18_bits_exceptionVec_11 = this.vif.mon_mp.mon_cb.io_writeback_18_bits_exceptionVec_11;
        io_writeback_18_bits_exceptionVec_12 = this.vif.mon_mp.mon_cb.io_writeback_18_bits_exceptionVec_12;
        io_writeback_18_bits_exceptionVec_13 = this.vif.mon_mp.mon_cb.io_writeback_18_bits_exceptionVec_13;
        io_writeback_18_bits_exceptionVec_14 = this.vif.mon_mp.mon_cb.io_writeback_18_bits_exceptionVec_14;
        io_writeback_18_bits_exceptionVec_15 = this.vif.mon_mp.mon_cb.io_writeback_18_bits_exceptionVec_15;
        io_writeback_18_bits_exceptionVec_16 = this.vif.mon_mp.mon_cb.io_writeback_18_bits_exceptionVec_16;
        io_writeback_18_bits_exceptionVec_17 = this.vif.mon_mp.mon_cb.io_writeback_18_bits_exceptionVec_17;
        io_writeback_18_bits_exceptionVec_18 = this.vif.mon_mp.mon_cb.io_writeback_18_bits_exceptionVec_18;
        io_writeback_18_bits_exceptionVec_19 = this.vif.mon_mp.mon_cb.io_writeback_18_bits_exceptionVec_19;
        io_writeback_18_bits_exceptionVec_20 = this.vif.mon_mp.mon_cb.io_writeback_18_bits_exceptionVec_20;
        io_writeback_18_bits_exceptionVec_21 = this.vif.mon_mp.mon_cb.io_writeback_18_bits_exceptionVec_21;
        io_writeback_18_bits_exceptionVec_22 = this.vif.mon_mp.mon_cb.io_writeback_18_bits_exceptionVec_22;
        io_writeback_18_bits_exceptionVec_23 = this.vif.mon_mp.mon_cb.io_writeback_18_bits_exceptionVec_23;
        io_writeback_18_bits_flushPipe = this.vif.mon_mp.mon_cb.io_writeback_18_bits_flushPipe;
        io_writeback_18_bits_sqIdx_flag = this.vif.mon_mp.mon_cb.io_writeback_18_bits_sqIdx_flag;
        io_writeback_18_bits_sqIdx_value = this.vif.mon_mp.mon_cb.io_writeback_18_bits_sqIdx_value;
        io_writeback_18_bits_trigger = this.vif.mon_mp.mon_cb.io_writeback_18_bits_trigger;
        io_writeback_18_bits_debug_isMMIO = this.vif.mon_mp.mon_cb.io_writeback_18_bits_debug_isMMIO;
        io_writeback_18_bits_debug_isNCIO = this.vif.mon_mp.mon_cb.io_writeback_18_bits_debug_isNCIO;
        io_writeback_18_bits_debug_isPerfCnt = this.vif.mon_mp.mon_cb.io_writeback_18_bits_debug_isPerfCnt;
        io_writeback_18_bits_debug_paddr = this.vif.mon_mp.mon_cb.io_writeback_18_bits_debug_paddr;
        io_writeback_18_bits_debug_vaddr = this.vif.mon_mp.mon_cb.io_writeback_18_bits_debug_vaddr;
        io_writeback_18_bits_debugInfo_eliminatedMove = this.vif.mon_mp.mon_cb.io_writeback_18_bits_debugInfo_eliminatedMove;
        io_writeback_18_bits_debugInfo_renameTime = this.vif.mon_mp.mon_cb.io_writeback_18_bits_debugInfo_renameTime;
        io_writeback_18_bits_debugInfo_dispatchTime = this.vif.mon_mp.mon_cb.io_writeback_18_bits_debugInfo_dispatchTime;
        io_writeback_18_bits_debugInfo_enqRsTime = this.vif.mon_mp.mon_cb.io_writeback_18_bits_debugInfo_enqRsTime;
        io_writeback_18_bits_debugInfo_selectTime = this.vif.mon_mp.mon_cb.io_writeback_18_bits_debugInfo_selectTime;
        io_writeback_18_bits_debugInfo_issueTime = this.vif.mon_mp.mon_cb.io_writeback_18_bits_debugInfo_issueTime;
        io_writeback_18_bits_debugInfo_writebackTime = this.vif.mon_mp.mon_cb.io_writeback_18_bits_debugInfo_writebackTime;
        io_writeback_18_bits_debugInfo_runahead_checkpoint_id = this.vif.mon_mp.mon_cb.io_writeback_18_bits_debugInfo_runahead_checkpoint_id;
        io_writeback_18_bits_debugInfo_tlbFirstReqTime = this.vif.mon_mp.mon_cb.io_writeback_18_bits_debugInfo_tlbFirstReqTime;
        io_writeback_18_bits_debugInfo_tlbRespTime = this.vif.mon_mp.mon_cb.io_writeback_18_bits_debugInfo_tlbRespTime;
        io_writeback_18_bits_debug_seqNum = this.vif.mon_mp.mon_cb.io_writeback_18_bits_debug_seqNum;
        io_writeback_17_valid = this.vif.mon_mp.mon_cb.io_writeback_17_valid;
        io_writeback_17_bits_data_0 = this.vif.mon_mp.mon_cb.io_writeback_17_bits_data_0;
        io_writeback_17_bits_data_1 = this.vif.mon_mp.mon_cb.io_writeback_17_bits_data_1;
        io_writeback_17_bits_data_2 = this.vif.mon_mp.mon_cb.io_writeback_17_bits_data_2;
        io_writeback_17_bits_pdest = this.vif.mon_mp.mon_cb.io_writeback_17_bits_pdest;
        io_writeback_17_bits_robIdx_flag = this.vif.mon_mp.mon_cb.io_writeback_17_bits_robIdx_flag;
        io_writeback_17_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_writeback_17_bits_robIdx_value;
        io_writeback_17_bits_vecWen = this.vif.mon_mp.mon_cb.io_writeback_17_bits_vecWen;
        io_writeback_17_bits_v0Wen = this.vif.mon_mp.mon_cb.io_writeback_17_bits_v0Wen;
        io_writeback_17_bits_fflags = this.vif.mon_mp.mon_cb.io_writeback_17_bits_fflags;
        io_writeback_17_bits_wflags = this.vif.mon_mp.mon_cb.io_writeback_17_bits_wflags;
        io_writeback_17_bits_debugInfo_eliminatedMove = this.vif.mon_mp.mon_cb.io_writeback_17_bits_debugInfo_eliminatedMove;
        io_writeback_17_bits_debugInfo_renameTime = this.vif.mon_mp.mon_cb.io_writeback_17_bits_debugInfo_renameTime;
        io_writeback_17_bits_debugInfo_dispatchTime = this.vif.mon_mp.mon_cb.io_writeback_17_bits_debugInfo_dispatchTime;
        io_writeback_17_bits_debugInfo_enqRsTime = this.vif.mon_mp.mon_cb.io_writeback_17_bits_debugInfo_enqRsTime;
        io_writeback_17_bits_debugInfo_selectTime = this.vif.mon_mp.mon_cb.io_writeback_17_bits_debugInfo_selectTime;
        io_writeback_17_bits_debugInfo_issueTime = this.vif.mon_mp.mon_cb.io_writeback_17_bits_debugInfo_issueTime;
        io_writeback_17_bits_debugInfo_writebackTime = this.vif.mon_mp.mon_cb.io_writeback_17_bits_debugInfo_writebackTime;
        io_writeback_17_bits_debugInfo_runahead_checkpoint_id = this.vif.mon_mp.mon_cb.io_writeback_17_bits_debugInfo_runahead_checkpoint_id;
        io_writeback_17_bits_debugInfo_tlbFirstReqTime = this.vif.mon_mp.mon_cb.io_writeback_17_bits_debugInfo_tlbFirstReqTime;
        io_writeback_17_bits_debugInfo_tlbRespTime = this.vif.mon_mp.mon_cb.io_writeback_17_bits_debugInfo_tlbRespTime;
        io_writeback_17_bits_debug_seqNum = this.vif.mon_mp.mon_cb.io_writeback_17_bits_debug_seqNum;
        io_writeback_16_valid = this.vif.mon_mp.mon_cb.io_writeback_16_valid;
        io_writeback_16_bits_data_0 = this.vif.mon_mp.mon_cb.io_writeback_16_bits_data_0;
        io_writeback_16_bits_data_1 = this.vif.mon_mp.mon_cb.io_writeback_16_bits_data_1;
        io_writeback_16_bits_data_2 = this.vif.mon_mp.mon_cb.io_writeback_16_bits_data_2;
        io_writeback_16_bits_data_3 = this.vif.mon_mp.mon_cb.io_writeback_16_bits_data_3;
        io_writeback_16_bits_pdest = this.vif.mon_mp.mon_cb.io_writeback_16_bits_pdest;
        io_writeback_16_bits_robIdx_flag = this.vif.mon_mp.mon_cb.io_writeback_16_bits_robIdx_flag;
        io_writeback_16_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_writeback_16_bits_robIdx_value;
        io_writeback_16_bits_fpWen = this.vif.mon_mp.mon_cb.io_writeback_16_bits_fpWen;
        io_writeback_16_bits_vecWen = this.vif.mon_mp.mon_cb.io_writeback_16_bits_vecWen;
        io_writeback_16_bits_v0Wen = this.vif.mon_mp.mon_cb.io_writeback_16_bits_v0Wen;
        io_writeback_16_bits_fflags = this.vif.mon_mp.mon_cb.io_writeback_16_bits_fflags;
        io_writeback_16_bits_wflags = this.vif.mon_mp.mon_cb.io_writeback_16_bits_wflags;
        io_writeback_16_bits_debugInfo_eliminatedMove = this.vif.mon_mp.mon_cb.io_writeback_16_bits_debugInfo_eliminatedMove;
        io_writeback_16_bits_debugInfo_renameTime = this.vif.mon_mp.mon_cb.io_writeback_16_bits_debugInfo_renameTime;
        io_writeback_16_bits_debugInfo_dispatchTime = this.vif.mon_mp.mon_cb.io_writeback_16_bits_debugInfo_dispatchTime;
        io_writeback_16_bits_debugInfo_enqRsTime = this.vif.mon_mp.mon_cb.io_writeback_16_bits_debugInfo_enqRsTime;
        io_writeback_16_bits_debugInfo_selectTime = this.vif.mon_mp.mon_cb.io_writeback_16_bits_debugInfo_selectTime;
        io_writeback_16_bits_debugInfo_issueTime = this.vif.mon_mp.mon_cb.io_writeback_16_bits_debugInfo_issueTime;
        io_writeback_16_bits_debugInfo_writebackTime = this.vif.mon_mp.mon_cb.io_writeback_16_bits_debugInfo_writebackTime;
        io_writeback_16_bits_debugInfo_runahead_checkpoint_id = this.vif.mon_mp.mon_cb.io_writeback_16_bits_debugInfo_runahead_checkpoint_id;
        io_writeback_16_bits_debugInfo_tlbFirstReqTime = this.vif.mon_mp.mon_cb.io_writeback_16_bits_debugInfo_tlbFirstReqTime;
        io_writeback_16_bits_debugInfo_tlbRespTime = this.vif.mon_mp.mon_cb.io_writeback_16_bits_debugInfo_tlbRespTime;
        io_writeback_16_bits_debug_seqNum = this.vif.mon_mp.mon_cb.io_writeback_16_bits_debug_seqNum;
        io_writeback_15_valid = this.vif.mon_mp.mon_cb.io_writeback_15_valid;
        io_writeback_15_bits_data_0 = this.vif.mon_mp.mon_cb.io_writeback_15_bits_data_0;
        io_writeback_15_bits_data_1 = this.vif.mon_mp.mon_cb.io_writeback_15_bits_data_1;
        io_writeback_15_bits_data_2 = this.vif.mon_mp.mon_cb.io_writeback_15_bits_data_2;
        io_writeback_15_bits_pdest = this.vif.mon_mp.mon_cb.io_writeback_15_bits_pdest;
        io_writeback_15_bits_robIdx_flag = this.vif.mon_mp.mon_cb.io_writeback_15_bits_robIdx_flag;
        io_writeback_15_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_writeback_15_bits_robIdx_value;
        io_writeback_15_bits_vecWen = this.vif.mon_mp.mon_cb.io_writeback_15_bits_vecWen;
        io_writeback_15_bits_v0Wen = this.vif.mon_mp.mon_cb.io_writeback_15_bits_v0Wen;
        io_writeback_15_bits_fflags = this.vif.mon_mp.mon_cb.io_writeback_15_bits_fflags;
        io_writeback_15_bits_wflags = this.vif.mon_mp.mon_cb.io_writeback_15_bits_wflags;
        io_writeback_15_bits_vxsat = this.vif.mon_mp.mon_cb.io_writeback_15_bits_vxsat;
        io_writeback_15_bits_debugInfo_eliminatedMove = this.vif.mon_mp.mon_cb.io_writeback_15_bits_debugInfo_eliminatedMove;
        io_writeback_15_bits_debugInfo_renameTime = this.vif.mon_mp.mon_cb.io_writeback_15_bits_debugInfo_renameTime;
        io_writeback_15_bits_debugInfo_dispatchTime = this.vif.mon_mp.mon_cb.io_writeback_15_bits_debugInfo_dispatchTime;
        io_writeback_15_bits_debugInfo_enqRsTime = this.vif.mon_mp.mon_cb.io_writeback_15_bits_debugInfo_enqRsTime;
        io_writeback_15_bits_debugInfo_selectTime = this.vif.mon_mp.mon_cb.io_writeback_15_bits_debugInfo_selectTime;
        io_writeback_15_bits_debugInfo_issueTime = this.vif.mon_mp.mon_cb.io_writeback_15_bits_debugInfo_issueTime;
        io_writeback_15_bits_debugInfo_writebackTime = this.vif.mon_mp.mon_cb.io_writeback_15_bits_debugInfo_writebackTime;
        io_writeback_15_bits_debugInfo_runahead_checkpoint_id = this.vif.mon_mp.mon_cb.io_writeback_15_bits_debugInfo_runahead_checkpoint_id;
        io_writeback_15_bits_debugInfo_tlbFirstReqTime = this.vif.mon_mp.mon_cb.io_writeback_15_bits_debugInfo_tlbFirstReqTime;
        io_writeback_15_bits_debugInfo_tlbRespTime = this.vif.mon_mp.mon_cb.io_writeback_15_bits_debugInfo_tlbRespTime;
        io_writeback_15_bits_debug_seqNum = this.vif.mon_mp.mon_cb.io_writeback_15_bits_debug_seqNum;
        io_writeback_14_valid = this.vif.mon_mp.mon_cb.io_writeback_14_valid;
        io_writeback_14_bits_data_0 = this.vif.mon_mp.mon_cb.io_writeback_14_bits_data_0;
        io_writeback_14_bits_data_1 = this.vif.mon_mp.mon_cb.io_writeback_14_bits_data_1;
        io_writeback_14_bits_data_2 = this.vif.mon_mp.mon_cb.io_writeback_14_bits_data_2;
        io_writeback_14_bits_data_3 = this.vif.mon_mp.mon_cb.io_writeback_14_bits_data_3;
        io_writeback_14_bits_data_4 = this.vif.mon_mp.mon_cb.io_writeback_14_bits_data_4;
        io_writeback_14_bits_data_5 = this.vif.mon_mp.mon_cb.io_writeback_14_bits_data_5;
        io_writeback_14_bits_pdest = this.vif.mon_mp.mon_cb.io_writeback_14_bits_pdest;
        io_writeback_14_bits_robIdx_flag = this.vif.mon_mp.mon_cb.io_writeback_14_bits_robIdx_flag;
        io_writeback_14_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_writeback_14_bits_robIdx_value;
        io_writeback_14_bits_intWen = this.vif.mon_mp.mon_cb.io_writeback_14_bits_intWen;
        io_writeback_14_bits_fpWen = this.vif.mon_mp.mon_cb.io_writeback_14_bits_fpWen;
        io_writeback_14_bits_vecWen = this.vif.mon_mp.mon_cb.io_writeback_14_bits_vecWen;
        io_writeback_14_bits_v0Wen = this.vif.mon_mp.mon_cb.io_writeback_14_bits_v0Wen;
        io_writeback_14_bits_vlWen = this.vif.mon_mp.mon_cb.io_writeback_14_bits_vlWen;
        io_writeback_14_bits_fflags = this.vif.mon_mp.mon_cb.io_writeback_14_bits_fflags;
        io_writeback_14_bits_wflags = this.vif.mon_mp.mon_cb.io_writeback_14_bits_wflags;
        io_writeback_14_bits_exceptionVec_2 = this.vif.mon_mp.mon_cb.io_writeback_14_bits_exceptionVec_2;
        io_writeback_14_bits_debugInfo_eliminatedMove = this.vif.mon_mp.mon_cb.io_writeback_14_bits_debugInfo_eliminatedMove;
        io_writeback_14_bits_debugInfo_renameTime = this.vif.mon_mp.mon_cb.io_writeback_14_bits_debugInfo_renameTime;
        io_writeback_14_bits_debugInfo_dispatchTime = this.vif.mon_mp.mon_cb.io_writeback_14_bits_debugInfo_dispatchTime;
        io_writeback_14_bits_debugInfo_enqRsTime = this.vif.mon_mp.mon_cb.io_writeback_14_bits_debugInfo_enqRsTime;
        io_writeback_14_bits_debugInfo_selectTime = this.vif.mon_mp.mon_cb.io_writeback_14_bits_debugInfo_selectTime;
        io_writeback_14_bits_debugInfo_issueTime = this.vif.mon_mp.mon_cb.io_writeback_14_bits_debugInfo_issueTime;
        io_writeback_14_bits_debugInfo_writebackTime = this.vif.mon_mp.mon_cb.io_writeback_14_bits_debugInfo_writebackTime;
        io_writeback_14_bits_debugInfo_runahead_checkpoint_id = this.vif.mon_mp.mon_cb.io_writeback_14_bits_debugInfo_runahead_checkpoint_id;
        io_writeback_14_bits_debugInfo_tlbFirstReqTime = this.vif.mon_mp.mon_cb.io_writeback_14_bits_debugInfo_tlbFirstReqTime;
        io_writeback_14_bits_debugInfo_tlbRespTime = this.vif.mon_mp.mon_cb.io_writeback_14_bits_debugInfo_tlbRespTime;
        io_writeback_14_bits_debug_seqNum = this.vif.mon_mp.mon_cb.io_writeback_14_bits_debug_seqNum;
        io_writeback_13_valid = this.vif.mon_mp.mon_cb.io_writeback_13_valid;
        io_writeback_13_bits_data_0 = this.vif.mon_mp.mon_cb.io_writeback_13_bits_data_0;
        io_writeback_13_bits_data_1 = this.vif.mon_mp.mon_cb.io_writeback_13_bits_data_1;
        io_writeback_13_bits_data_2 = this.vif.mon_mp.mon_cb.io_writeback_13_bits_data_2;
        io_writeback_13_bits_pdest = this.vif.mon_mp.mon_cb.io_writeback_13_bits_pdest;
        io_writeback_13_bits_robIdx_flag = this.vif.mon_mp.mon_cb.io_writeback_13_bits_robIdx_flag;
        io_writeback_13_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_writeback_13_bits_robIdx_value;
        io_writeback_13_bits_vecWen = this.vif.mon_mp.mon_cb.io_writeback_13_bits_vecWen;
        io_writeback_13_bits_v0Wen = this.vif.mon_mp.mon_cb.io_writeback_13_bits_v0Wen;
        io_writeback_13_bits_fflags = this.vif.mon_mp.mon_cb.io_writeback_13_bits_fflags;
        io_writeback_13_bits_wflags = this.vif.mon_mp.mon_cb.io_writeback_13_bits_wflags;
        io_writeback_13_bits_vxsat = this.vif.mon_mp.mon_cb.io_writeback_13_bits_vxsat;
        io_writeback_13_bits_exceptionVec_2 = this.vif.mon_mp.mon_cb.io_writeback_13_bits_exceptionVec_2;
        io_writeback_13_bits_debugInfo_eliminatedMove = this.vif.mon_mp.mon_cb.io_writeback_13_bits_debugInfo_eliminatedMove;
        io_writeback_13_bits_debugInfo_renameTime = this.vif.mon_mp.mon_cb.io_writeback_13_bits_debugInfo_renameTime;
        io_writeback_13_bits_debugInfo_dispatchTime = this.vif.mon_mp.mon_cb.io_writeback_13_bits_debugInfo_dispatchTime;
        io_writeback_13_bits_debugInfo_enqRsTime = this.vif.mon_mp.mon_cb.io_writeback_13_bits_debugInfo_enqRsTime;
        io_writeback_13_bits_debugInfo_selectTime = this.vif.mon_mp.mon_cb.io_writeback_13_bits_debugInfo_selectTime;
        io_writeback_13_bits_debugInfo_issueTime = this.vif.mon_mp.mon_cb.io_writeback_13_bits_debugInfo_issueTime;
        io_writeback_13_bits_debugInfo_writebackTime = this.vif.mon_mp.mon_cb.io_writeback_13_bits_debugInfo_writebackTime;
        io_writeback_13_bits_debugInfo_runahead_checkpoint_id = this.vif.mon_mp.mon_cb.io_writeback_13_bits_debugInfo_runahead_checkpoint_id;
        io_writeback_13_bits_debugInfo_tlbFirstReqTime = this.vif.mon_mp.mon_cb.io_writeback_13_bits_debugInfo_tlbFirstReqTime;
        io_writeback_13_bits_debugInfo_tlbRespTime = this.vif.mon_mp.mon_cb.io_writeback_13_bits_debugInfo_tlbRespTime;
        io_writeback_13_bits_debug_seqNum = this.vif.mon_mp.mon_cb.io_writeback_13_bits_debug_seqNum;
        io_writeback_7_valid = this.vif.mon_mp.mon_cb.io_writeback_7_valid;
        io_writeback_7_bits_data_0 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_data_0;
        io_writeback_7_bits_data_1 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_data_1;
        io_writeback_7_bits_pdest = this.vif.mon_mp.mon_cb.io_writeback_7_bits_pdest;
        io_writeback_7_bits_robIdx_flag = this.vif.mon_mp.mon_cb.io_writeback_7_bits_robIdx_flag;
        io_writeback_7_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_writeback_7_bits_robIdx_value;
        io_writeback_7_bits_intWen = this.vif.mon_mp.mon_cb.io_writeback_7_bits_intWen;
        io_writeback_7_bits_redirect_valid = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_valid;
        io_writeback_7_bits_redirect_bits_isRVC = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_isRVC;
        io_writeback_7_bits_redirect_bits_robIdx_flag = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_robIdx_flag;
        io_writeback_7_bits_redirect_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_robIdx_value;
        io_writeback_7_bits_redirect_bits_ftqIdx_flag = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_ftqIdx_flag;
        io_writeback_7_bits_redirect_bits_ftqIdx_value = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_ftqIdx_value;
        io_writeback_7_bits_redirect_bits_ftqOffset = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_ftqOffset;
        io_writeback_7_bits_redirect_bits_level = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_level;
        io_writeback_7_bits_redirect_bits_interrupt = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_interrupt;
        io_writeback_7_bits_redirect_bits_cfiUpdate_pc = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pc;
        io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid;
        io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC;
        io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType;
        io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall;
        io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet;
        io_writeback_7_bits_redirect_bits_cfiUpdate_ssp = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_ssp;
        io_writeback_7_bits_redirect_bits_cfiUpdate_sctr = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_sctr;
        io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag;
        io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value;
        io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag;
        io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value;
        io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag;
        io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value;
        io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr;
        io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist;
        io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist;
        io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist;
        io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist;
        io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist;
        io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist;
        io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist;
        io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist;
        io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist;
        io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist;
        io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist;
        io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist;
        io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist;
        io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist;
        io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist;
        io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist;
        io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist;
        io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist;
        io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0;
        io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1;
        io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2;
        io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3;
        io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0;
        io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1;
        io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2;
        io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3;
        io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0;
        io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1;
        io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2;
        io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3;
        io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0;
        io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1;
        io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2;
        io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3;
        io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0;
        io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1;
        io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2;
        io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3;
        io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0;
        io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1;
        io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2;
        io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3;
        io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH;
        io_writeback_7_bits_redirect_bits_cfiUpdate_ghr = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_ghr;
        io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag;
        io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value;
        io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0;
        io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1;
        io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit;
        io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit;
        io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit;
        io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken;
        io_writeback_7_bits_redirect_bits_cfiUpdate_target = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_target;
        io_writeback_7_bits_redirect_bits_cfiUpdate_taken = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_taken;
        io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred;
        io_writeback_7_bits_redirect_bits_cfiUpdate_shift = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_shift;
        io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist;
        io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF;
        io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF;
        io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF;
        io_writeback_7_bits_redirect_bits_fullTarget = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_fullTarget;
        io_writeback_7_bits_redirect_bits_stFtqIdx_flag = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_stFtqIdx_flag;
        io_writeback_7_bits_redirect_bits_stFtqIdx_value = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_stFtqIdx_value;
        io_writeback_7_bits_redirect_bits_stFtqOffset = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_stFtqOffset;
        io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id;
        io_writeback_7_bits_redirect_bits_debugIsCtrl = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_debugIsCtrl;
        io_writeback_7_bits_redirect_bits_debugIsMemVio = this.vif.mon_mp.mon_cb.io_writeback_7_bits_redirect_bits_debugIsMemVio;
        io_writeback_7_bits_exceptionVec_2 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_exceptionVec_2;
        io_writeback_7_bits_exceptionVec_3 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_exceptionVec_3;
        io_writeback_7_bits_exceptionVec_8 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_exceptionVec_8;
        io_writeback_7_bits_exceptionVec_9 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_exceptionVec_9;
        io_writeback_7_bits_exceptionVec_10 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_exceptionVec_10;
        io_writeback_7_bits_exceptionVec_11 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_exceptionVec_11;
        io_writeback_7_bits_exceptionVec_22 = this.vif.mon_mp.mon_cb.io_writeback_7_bits_exceptionVec_22;
        io_writeback_7_bits_flushPipe = this.vif.mon_mp.mon_cb.io_writeback_7_bits_flushPipe;
        io_writeback_7_bits_predecodeInfo_valid = this.vif.mon_mp.mon_cb.io_writeback_7_bits_predecodeInfo_valid;
        io_writeback_7_bits_predecodeInfo_isRVC = this.vif.mon_mp.mon_cb.io_writeback_7_bits_predecodeInfo_isRVC;
        io_writeback_7_bits_predecodeInfo_brType = this.vif.mon_mp.mon_cb.io_writeback_7_bits_predecodeInfo_brType;
        io_writeback_7_bits_predecodeInfo_isCall = this.vif.mon_mp.mon_cb.io_writeback_7_bits_predecodeInfo_isCall;
        io_writeback_7_bits_predecodeInfo_isRet = this.vif.mon_mp.mon_cb.io_writeback_7_bits_predecodeInfo_isRet;
        io_writeback_7_bits_debug_isPerfCnt = this.vif.mon_mp.mon_cb.io_writeback_7_bits_debug_isPerfCnt;
        io_writeback_7_bits_debugInfo_eliminatedMove = this.vif.mon_mp.mon_cb.io_writeback_7_bits_debugInfo_eliminatedMove;
        io_writeback_7_bits_debugInfo_renameTime = this.vif.mon_mp.mon_cb.io_writeback_7_bits_debugInfo_renameTime;
        io_writeback_7_bits_debugInfo_dispatchTime = this.vif.mon_mp.mon_cb.io_writeback_7_bits_debugInfo_dispatchTime;
        io_writeback_7_bits_debugInfo_enqRsTime = this.vif.mon_mp.mon_cb.io_writeback_7_bits_debugInfo_enqRsTime;
        io_writeback_7_bits_debugInfo_selectTime = this.vif.mon_mp.mon_cb.io_writeback_7_bits_debugInfo_selectTime;
        io_writeback_7_bits_debugInfo_issueTime = this.vif.mon_mp.mon_cb.io_writeback_7_bits_debugInfo_issueTime;
        io_writeback_7_bits_debugInfo_writebackTime = this.vif.mon_mp.mon_cb.io_writeback_7_bits_debugInfo_writebackTime;
        io_writeback_7_bits_debugInfo_runahead_checkpoint_id = this.vif.mon_mp.mon_cb.io_writeback_7_bits_debugInfo_runahead_checkpoint_id;
        io_writeback_7_bits_debugInfo_tlbFirstReqTime = this.vif.mon_mp.mon_cb.io_writeback_7_bits_debugInfo_tlbFirstReqTime;
        io_writeback_7_bits_debugInfo_tlbRespTime = this.vif.mon_mp.mon_cb.io_writeback_7_bits_debugInfo_tlbRespTime;
        io_writeback_7_bits_debug_seqNum = this.vif.mon_mp.mon_cb.io_writeback_7_bits_debug_seqNum;
        io_writeback_5_valid = this.vif.mon_mp.mon_cb.io_writeback_5_valid;
        io_writeback_5_bits_redirect_valid = this.vif.mon_mp.mon_cb.io_writeback_5_bits_redirect_valid;
        io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred = this.vif.mon_mp.mon_cb.io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred;
        io_writeback_3_valid = this.vif.mon_mp.mon_cb.io_writeback_3_valid;
        io_writeback_3_bits_redirect_valid = this.vif.mon_mp.mon_cb.io_writeback_3_bits_redirect_valid;
        io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred = this.vif.mon_mp.mon_cb.io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred;
        io_writeback_1_valid = this.vif.mon_mp.mon_cb.io_writeback_1_valid;
        io_writeback_1_bits_redirect_valid = this.vif.mon_mp.mon_cb.io_writeback_1_bits_redirect_valid;
        io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred = this.vif.mon_mp.mon_cb.io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred;
        io_exuWriteback_26_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_26_valid;
        io_exuWriteback_26_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_26_bits_robIdx_value;
        io_exuWriteback_25_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_25_valid;
        io_exuWriteback_25_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_25_bits_robIdx_value;
        io_exuWriteback_24_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_24_valid;
        io_exuWriteback_24_bits_data_0 = this.vif.mon_mp.mon_cb.io_exuWriteback_24_bits_data_0;
        io_exuWriteback_24_bits_pdest = this.vif.mon_mp.mon_cb.io_exuWriteback_24_bits_pdest;
        io_exuWriteback_24_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_24_bits_robIdx_value;
        io_exuWriteback_24_bits_vecWen = this.vif.mon_mp.mon_cb.io_exuWriteback_24_bits_vecWen;
        io_exuWriteback_24_bits_v0Wen = this.vif.mon_mp.mon_cb.io_exuWriteback_24_bits_v0Wen;
        io_exuWriteback_24_bits_vls_vdIdx = this.vif.mon_mp.mon_cb.io_exuWriteback_24_bits_vls_vdIdx;
        io_exuWriteback_24_bits_debug_isMMIO = this.vif.mon_mp.mon_cb.io_exuWriteback_24_bits_debug_isMMIO;
        io_exuWriteback_24_bits_debug_isNCIO = this.vif.mon_mp.mon_cb.io_exuWriteback_24_bits_debug_isNCIO;
        io_exuWriteback_24_bits_debug_isPerfCnt = this.vif.mon_mp.mon_cb.io_exuWriteback_24_bits_debug_isPerfCnt;
        io_exuWriteback_24_bits_debug_paddr = this.vif.mon_mp.mon_cb.io_exuWriteback_24_bits_debug_paddr;
        io_exuWriteback_23_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_23_valid;
        io_exuWriteback_23_bits_data_0 = this.vif.mon_mp.mon_cb.io_exuWriteback_23_bits_data_0;
        io_exuWriteback_23_bits_pdest = this.vif.mon_mp.mon_cb.io_exuWriteback_23_bits_pdest;
        io_exuWriteback_23_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_23_bits_robIdx_value;
        io_exuWriteback_23_bits_vecWen = this.vif.mon_mp.mon_cb.io_exuWriteback_23_bits_vecWen;
        io_exuWriteback_23_bits_v0Wen = this.vif.mon_mp.mon_cb.io_exuWriteback_23_bits_v0Wen;
        io_exuWriteback_23_bits_vls_vdIdx = this.vif.mon_mp.mon_cb.io_exuWriteback_23_bits_vls_vdIdx;
        io_exuWriteback_23_bits_debug_isMMIO = this.vif.mon_mp.mon_cb.io_exuWriteback_23_bits_debug_isMMIO;
        io_exuWriteback_23_bits_debug_isNCIO = this.vif.mon_mp.mon_cb.io_exuWriteback_23_bits_debug_isNCIO;
        io_exuWriteback_23_bits_debug_isPerfCnt = this.vif.mon_mp.mon_cb.io_exuWriteback_23_bits_debug_isPerfCnt;
        io_exuWriteback_23_bits_debug_paddr = this.vif.mon_mp.mon_cb.io_exuWriteback_23_bits_debug_paddr;
        io_exuWriteback_22_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_22_valid;
        io_exuWriteback_22_bits_data_0 = this.vif.mon_mp.mon_cb.io_exuWriteback_22_bits_data_0;
        io_exuWriteback_22_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_22_bits_robIdx_value;
        io_exuWriteback_22_bits_lqIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_22_bits_lqIdx_value;
        io_exuWriteback_22_bits_debug_isMMIO = this.vif.mon_mp.mon_cb.io_exuWriteback_22_bits_debug_isMMIO;
        io_exuWriteback_22_bits_debug_isNCIO = this.vif.mon_mp.mon_cb.io_exuWriteback_22_bits_debug_isNCIO;
        io_exuWriteback_22_bits_debug_isPerfCnt = this.vif.mon_mp.mon_cb.io_exuWriteback_22_bits_debug_isPerfCnt;
        io_exuWriteback_22_bits_debug_paddr = this.vif.mon_mp.mon_cb.io_exuWriteback_22_bits_debug_paddr;
        io_exuWriteback_21_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_21_valid;
        io_exuWriteback_21_bits_data_0 = this.vif.mon_mp.mon_cb.io_exuWriteback_21_bits_data_0;
        io_exuWriteback_21_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_21_bits_robIdx_value;
        io_exuWriteback_21_bits_lqIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_21_bits_lqIdx_value;
        io_exuWriteback_21_bits_debug_isMMIO = this.vif.mon_mp.mon_cb.io_exuWriteback_21_bits_debug_isMMIO;
        io_exuWriteback_21_bits_debug_isNCIO = this.vif.mon_mp.mon_cb.io_exuWriteback_21_bits_debug_isNCIO;
        io_exuWriteback_21_bits_debug_isPerfCnt = this.vif.mon_mp.mon_cb.io_exuWriteback_21_bits_debug_isPerfCnt;
        io_exuWriteback_21_bits_debug_paddr = this.vif.mon_mp.mon_cb.io_exuWriteback_21_bits_debug_paddr;
        io_exuWriteback_20_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_20_valid;
        io_exuWriteback_20_bits_data_0 = this.vif.mon_mp.mon_cb.io_exuWriteback_20_bits_data_0;
        io_exuWriteback_20_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_20_bits_robIdx_value;
        io_exuWriteback_20_bits_lqIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_20_bits_lqIdx_value;
        io_exuWriteback_20_bits_debug_isMMIO = this.vif.mon_mp.mon_cb.io_exuWriteback_20_bits_debug_isMMIO;
        io_exuWriteback_20_bits_debug_isNCIO = this.vif.mon_mp.mon_cb.io_exuWriteback_20_bits_debug_isNCIO;
        io_exuWriteback_20_bits_debug_isPerfCnt = this.vif.mon_mp.mon_cb.io_exuWriteback_20_bits_debug_isPerfCnt;
        io_exuWriteback_20_bits_debug_paddr = this.vif.mon_mp.mon_cb.io_exuWriteback_20_bits_debug_paddr;
        io_exuWriteback_19_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_19_valid;
        io_exuWriteback_19_bits_data_0 = this.vif.mon_mp.mon_cb.io_exuWriteback_19_bits_data_0;
        io_exuWriteback_19_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_19_bits_robIdx_value;
        io_exuWriteback_19_bits_sqIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_19_bits_sqIdx_value;
        io_exuWriteback_19_bits_debug_isMMIO = this.vif.mon_mp.mon_cb.io_exuWriteback_19_bits_debug_isMMIO;
        io_exuWriteback_19_bits_debug_isNCIO = this.vif.mon_mp.mon_cb.io_exuWriteback_19_bits_debug_isNCIO;
        io_exuWriteback_19_bits_debug_isPerfCnt = this.vif.mon_mp.mon_cb.io_exuWriteback_19_bits_debug_isPerfCnt;
        io_exuWriteback_19_bits_debug_paddr = this.vif.mon_mp.mon_cb.io_exuWriteback_19_bits_debug_paddr;
        io_exuWriteback_18_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_18_valid;
        io_exuWriteback_18_bits_data_0 = this.vif.mon_mp.mon_cb.io_exuWriteback_18_bits_data_0;
        io_exuWriteback_18_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_18_bits_robIdx_value;
        io_exuWriteback_18_bits_sqIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_18_bits_sqIdx_value;
        io_exuWriteback_18_bits_debug_isMMIO = this.vif.mon_mp.mon_cb.io_exuWriteback_18_bits_debug_isMMIO;
        io_exuWriteback_18_bits_debug_isNCIO = this.vif.mon_mp.mon_cb.io_exuWriteback_18_bits_debug_isNCIO;
        io_exuWriteback_18_bits_debug_isPerfCnt = this.vif.mon_mp.mon_cb.io_exuWriteback_18_bits_debug_isPerfCnt;
        io_exuWriteback_18_bits_debug_paddr = this.vif.mon_mp.mon_cb.io_exuWriteback_18_bits_debug_paddr;
        io_exuWriteback_17_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_17_valid;
        io_exuWriteback_17_bits_data_0 = this.vif.mon_mp.mon_cb.io_exuWriteback_17_bits_data_0;
        io_exuWriteback_17_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_17_bits_robIdx_value;
        io_exuWriteback_17_bits_fflags = this.vif.mon_mp.mon_cb.io_exuWriteback_17_bits_fflags;
        io_exuWriteback_17_bits_wflags = this.vif.mon_mp.mon_cb.io_exuWriteback_17_bits_wflags;
        io_exuWriteback_16_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_16_valid;
        io_exuWriteback_16_bits_data_0 = this.vif.mon_mp.mon_cb.io_exuWriteback_16_bits_data_0;
        io_exuWriteback_16_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_16_bits_robIdx_value;
        io_exuWriteback_16_bits_fflags = this.vif.mon_mp.mon_cb.io_exuWriteback_16_bits_fflags;
        io_exuWriteback_16_bits_wflags = this.vif.mon_mp.mon_cb.io_exuWriteback_16_bits_wflags;
        io_exuWriteback_15_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_15_valid;
        io_exuWriteback_15_bits_data_0 = this.vif.mon_mp.mon_cb.io_exuWriteback_15_bits_data_0;
        io_exuWriteback_15_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_15_bits_robIdx_value;
        io_exuWriteback_15_bits_fflags = this.vif.mon_mp.mon_cb.io_exuWriteback_15_bits_fflags;
        io_exuWriteback_15_bits_wflags = this.vif.mon_mp.mon_cb.io_exuWriteback_15_bits_wflags;
        io_exuWriteback_15_bits_vxsat = this.vif.mon_mp.mon_cb.io_exuWriteback_15_bits_vxsat;
        io_exuWriteback_14_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_14_valid;
        io_exuWriteback_14_bits_data_0 = this.vif.mon_mp.mon_cb.io_exuWriteback_14_bits_data_0;
        io_exuWriteback_14_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_14_bits_robIdx_value;
        io_exuWriteback_14_bits_fflags = this.vif.mon_mp.mon_cb.io_exuWriteback_14_bits_fflags;
        io_exuWriteback_14_bits_wflags = this.vif.mon_mp.mon_cb.io_exuWriteback_14_bits_wflags;
        io_exuWriteback_13_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_13_valid;
        io_exuWriteback_13_bits_data_0 = this.vif.mon_mp.mon_cb.io_exuWriteback_13_bits_data_0;
        io_exuWriteback_13_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_13_bits_robIdx_value;
        io_exuWriteback_13_bits_fflags = this.vif.mon_mp.mon_cb.io_exuWriteback_13_bits_fflags;
        io_exuWriteback_13_bits_wflags = this.vif.mon_mp.mon_cb.io_exuWriteback_13_bits_wflags;
        io_exuWriteback_13_bits_vxsat = this.vif.mon_mp.mon_cb.io_exuWriteback_13_bits_vxsat;
        io_exuWriteback_12_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_12_valid;
        io_exuWriteback_12_bits_data_0 = this.vif.mon_mp.mon_cb.io_exuWriteback_12_bits_data_0;
        io_exuWriteback_12_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_12_bits_robIdx_value;
        io_exuWriteback_12_bits_fflags = this.vif.mon_mp.mon_cb.io_exuWriteback_12_bits_fflags;
        io_exuWriteback_12_bits_wflags = this.vif.mon_mp.mon_cb.io_exuWriteback_12_bits_wflags;
        io_exuWriteback_11_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_11_valid;
        io_exuWriteback_11_bits_data_0 = this.vif.mon_mp.mon_cb.io_exuWriteback_11_bits_data_0;
        io_exuWriteback_11_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_11_bits_robIdx_value;
        io_exuWriteback_11_bits_fflags = this.vif.mon_mp.mon_cb.io_exuWriteback_11_bits_fflags;
        io_exuWriteback_11_bits_wflags = this.vif.mon_mp.mon_cb.io_exuWriteback_11_bits_wflags;
        io_exuWriteback_10_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_10_valid;
        io_exuWriteback_10_bits_data_0 = this.vif.mon_mp.mon_cb.io_exuWriteback_10_bits_data_0;
        io_exuWriteback_10_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_10_bits_robIdx_value;
        io_exuWriteback_10_bits_fflags = this.vif.mon_mp.mon_cb.io_exuWriteback_10_bits_fflags;
        io_exuWriteback_10_bits_wflags = this.vif.mon_mp.mon_cb.io_exuWriteback_10_bits_wflags;
        io_exuWriteback_9_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_9_valid;
        io_exuWriteback_9_bits_data_0 = this.vif.mon_mp.mon_cb.io_exuWriteback_9_bits_data_0;
        io_exuWriteback_9_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_9_bits_robIdx_value;
        io_exuWriteback_9_bits_fflags = this.vif.mon_mp.mon_cb.io_exuWriteback_9_bits_fflags;
        io_exuWriteback_9_bits_wflags = this.vif.mon_mp.mon_cb.io_exuWriteback_9_bits_wflags;
        io_exuWriteback_8_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_8_valid;
        io_exuWriteback_8_bits_data_0 = this.vif.mon_mp.mon_cb.io_exuWriteback_8_bits_data_0;
        io_exuWriteback_8_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_8_bits_robIdx_value;
        io_exuWriteback_8_bits_fflags = this.vif.mon_mp.mon_cb.io_exuWriteback_8_bits_fflags;
        io_exuWriteback_8_bits_wflags = this.vif.mon_mp.mon_cb.io_exuWriteback_8_bits_wflags;
        io_exuWriteback_7_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_7_valid;
        io_exuWriteback_7_bits_data_0 = this.vif.mon_mp.mon_cb.io_exuWriteback_7_bits_data_0;
        io_exuWriteback_7_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_7_bits_robIdx_value;
        io_exuWriteback_7_bits_debug_isPerfCnt = this.vif.mon_mp.mon_cb.io_exuWriteback_7_bits_debug_isPerfCnt;
        io_exuWriteback_6_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_6_valid;
        io_exuWriteback_6_bits_data_0 = this.vif.mon_mp.mon_cb.io_exuWriteback_6_bits_data_0;
        io_exuWriteback_6_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_6_bits_robIdx_value;
        io_exuWriteback_5_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_5_valid;
        io_exuWriteback_5_bits_data_0 = this.vif.mon_mp.mon_cb.io_exuWriteback_5_bits_data_0;
        io_exuWriteback_5_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_5_bits_robIdx_value;
        io_exuWriteback_5_bits_redirect_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_5_bits_redirect_valid;
        io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken = this.vif.mon_mp.mon_cb.io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken;
        io_exuWriteback_5_bits_fflags = this.vif.mon_mp.mon_cb.io_exuWriteback_5_bits_fflags;
        io_exuWriteback_5_bits_wflags = this.vif.mon_mp.mon_cb.io_exuWriteback_5_bits_wflags;
        io_exuWriteback_4_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_4_valid;
        io_exuWriteback_4_bits_data_0 = this.vif.mon_mp.mon_cb.io_exuWriteback_4_bits_data_0;
        io_exuWriteback_4_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_4_bits_robIdx_value;
        io_exuWriteback_3_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_3_valid;
        io_exuWriteback_3_bits_data_0 = this.vif.mon_mp.mon_cb.io_exuWriteback_3_bits_data_0;
        io_exuWriteback_3_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_3_bits_robIdx_value;
        io_exuWriteback_3_bits_redirect_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_3_bits_redirect_valid;
        io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken = this.vif.mon_mp.mon_cb.io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken;
        io_exuWriteback_2_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_2_valid;
        io_exuWriteback_2_bits_data_0 = this.vif.mon_mp.mon_cb.io_exuWriteback_2_bits_data_0;
        io_exuWriteback_2_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_2_bits_robIdx_value;
        io_exuWriteback_1_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_1_valid;
        io_exuWriteback_1_bits_data_0 = this.vif.mon_mp.mon_cb.io_exuWriteback_1_bits_data_0;
        io_exuWriteback_1_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_1_bits_robIdx_value;
        io_exuWriteback_1_bits_redirect_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_1_bits_redirect_valid;
        io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken = this.vif.mon_mp.mon_cb.io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken;
        io_exuWriteback_0_valid = this.vif.mon_mp.mon_cb.io_exuWriteback_0_valid;
        io_exuWriteback_0_bits_data_0 = this.vif.mon_mp.mon_cb.io_exuWriteback_0_bits_data_0;
        io_exuWriteback_0_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_exuWriteback_0_bits_robIdx_value;
        io_writebackNums_0_bits = this.vif.mon_mp.mon_cb.io_writebackNums_0_bits;
        io_writebackNums_1_bits = this.vif.mon_mp.mon_cb.io_writebackNums_1_bits;
        io_writebackNums_2_bits = this.vif.mon_mp.mon_cb.io_writebackNums_2_bits;
        io_writebackNums_3_bits = this.vif.mon_mp.mon_cb.io_writebackNums_3_bits;
        io_writebackNums_4_bits = this.vif.mon_mp.mon_cb.io_writebackNums_4_bits;
        io_writebackNums_5_bits = this.vif.mon_mp.mon_cb.io_writebackNums_5_bits;
        io_writebackNums_6_bits = this.vif.mon_mp.mon_cb.io_writebackNums_6_bits;
        io_writebackNums_7_bits = this.vif.mon_mp.mon_cb.io_writebackNums_7_bits;
        io_writebackNums_8_bits = this.vif.mon_mp.mon_cb.io_writebackNums_8_bits;
        io_writebackNums_9_bits = this.vif.mon_mp.mon_cb.io_writebackNums_9_bits;
        io_writebackNums_10_bits = this.vif.mon_mp.mon_cb.io_writebackNums_10_bits;
        io_writebackNums_11_bits = this.vif.mon_mp.mon_cb.io_writebackNums_11_bits;
        io_writebackNums_12_bits = this.vif.mon_mp.mon_cb.io_writebackNums_12_bits;
        io_writebackNums_13_bits = this.vif.mon_mp.mon_cb.io_writebackNums_13_bits;
        io_writebackNums_14_bits = this.vif.mon_mp.mon_cb.io_writebackNums_14_bits;
        io_writebackNums_15_bits = this.vif.mon_mp.mon_cb.io_writebackNums_15_bits;
        io_writebackNums_16_bits = this.vif.mon_mp.mon_cb.io_writebackNums_16_bits;
        io_writebackNums_17_bits = this.vif.mon_mp.mon_cb.io_writebackNums_17_bits;
        io_writebackNums_18_bits = this.vif.mon_mp.mon_cb.io_writebackNums_18_bits;
        io_writebackNums_19_bits = this.vif.mon_mp.mon_cb.io_writebackNums_19_bits;
        io_writebackNums_20_bits = this.vif.mon_mp.mon_cb.io_writebackNums_20_bits;
        io_writebackNums_21_bits = this.vif.mon_mp.mon_cb.io_writebackNums_21_bits;
        io_writebackNums_22_bits = this.vif.mon_mp.mon_cb.io_writebackNums_22_bits;
        io_writebackNums_23_bits = this.vif.mon_mp.mon_cb.io_writebackNums_23_bits;
        io_writebackNums_24_bits = this.vif.mon_mp.mon_cb.io_writebackNums_24_bits;
        io_writebackNeedFlush_0 = this.vif.mon_mp.mon_cb.io_writebackNeedFlush_0;
        io_writebackNeedFlush_1 = this.vif.mon_mp.mon_cb.io_writebackNeedFlush_1;
        io_writebackNeedFlush_2 = this.vif.mon_mp.mon_cb.io_writebackNeedFlush_2;
        io_writebackNeedFlush_6 = this.vif.mon_mp.mon_cb.io_writebackNeedFlush_6;
        io_writebackNeedFlush_7 = this.vif.mon_mp.mon_cb.io_writebackNeedFlush_7;
        io_writebackNeedFlush_8 = this.vif.mon_mp.mon_cb.io_writebackNeedFlush_8;
        io_writebackNeedFlush_9 = this.vif.mon_mp.mon_cb.io_writebackNeedFlush_9;
        io_writebackNeedFlush_10 = this.vif.mon_mp.mon_cb.io_writebackNeedFlush_10;
        io_writebackNeedFlush_11 = this.vif.mon_mp.mon_cb.io_writebackNeedFlush_11;
        io_writebackNeedFlush_12 = this.vif.mon_mp.mon_cb.io_writebackNeedFlush_12;

        if(this.cfg.xz_sw==tcnt_dec_base::ON & this.vif.rst_n==1'b1) begin
            `TCNT_CHECK_SIG_XZ(io_writeback_24_valid,io_writeback_24_valid,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_data_0,io_writeback_24_bits_data_0,128);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_pdest,io_writeback_24_bits_pdest,7);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_robIdx_flag,io_writeback_24_bits_robIdx_flag,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_robIdx_value,io_writeback_24_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vecWen,io_writeback_24_bits_vecWen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_v0Wen,io_writeback_24_bits_v0Wen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vlWen,io_writeback_24_bits_vlWen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_exceptionVec_0,io_writeback_24_bits_exceptionVec_0,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_exceptionVec_1,io_writeback_24_bits_exceptionVec_1,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_exceptionVec_2,io_writeback_24_bits_exceptionVec_2,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_exceptionVec_3,io_writeback_24_bits_exceptionVec_3,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_exceptionVec_4,io_writeback_24_bits_exceptionVec_4,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_exceptionVec_5,io_writeback_24_bits_exceptionVec_5,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_exceptionVec_6,io_writeback_24_bits_exceptionVec_6,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_exceptionVec_7,io_writeback_24_bits_exceptionVec_7,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_exceptionVec_8,io_writeback_24_bits_exceptionVec_8,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_exceptionVec_9,io_writeback_24_bits_exceptionVec_9,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_exceptionVec_10,io_writeback_24_bits_exceptionVec_10,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_exceptionVec_11,io_writeback_24_bits_exceptionVec_11,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_exceptionVec_12,io_writeback_24_bits_exceptionVec_12,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_exceptionVec_13,io_writeback_24_bits_exceptionVec_13,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_exceptionVec_14,io_writeback_24_bits_exceptionVec_14,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_exceptionVec_15,io_writeback_24_bits_exceptionVec_15,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_exceptionVec_16,io_writeback_24_bits_exceptionVec_16,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_exceptionVec_17,io_writeback_24_bits_exceptionVec_17,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_exceptionVec_18,io_writeback_24_bits_exceptionVec_18,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_exceptionVec_19,io_writeback_24_bits_exceptionVec_19,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_exceptionVec_20,io_writeback_24_bits_exceptionVec_20,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_exceptionVec_21,io_writeback_24_bits_exceptionVec_21,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_exceptionVec_22,io_writeback_24_bits_exceptionVec_22,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_exceptionVec_23,io_writeback_24_bits_exceptionVec_23,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_flushPipe,io_writeback_24_bits_flushPipe,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_replay,io_writeback_24_bits_replay,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_trigger,io_writeback_24_bits_trigger,4);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_vill,io_writeback_24_bits_vls_vpu_vill,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_vma,io_writeback_24_bits_vls_vpu_vma,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_vta,io_writeback_24_bits_vls_vpu_vta,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_vsew,io_writeback_24_bits_vls_vpu_vsew,2);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_vlmul,io_writeback_24_bits_vls_vpu_vlmul,3);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_specVill,io_writeback_24_bits_vls_vpu_specVill,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_specVma,io_writeback_24_bits_vls_vpu_specVma,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_specVta,io_writeback_24_bits_vls_vpu_specVta,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_specVsew,io_writeback_24_bits_vls_vpu_specVsew,2);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_specVlmul,io_writeback_24_bits_vls_vpu_specVlmul,3);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_vm,io_writeback_24_bits_vls_vpu_vm,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_vstart,io_writeback_24_bits_vls_vpu_vstart,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_frm,io_writeback_24_bits_vls_vpu_frm,3);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst,io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_fpu_isFP32Instr,io_writeback_24_bits_vls_vpu_fpu_isFP32Instr,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_fpu_isFP64Instr,io_writeback_24_bits_vls_vpu_fpu_isFP64Instr,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_fpu_isReduction,io_writeback_24_bits_vls_vpu_fpu_isReduction,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2,io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4,io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8,io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_vxrm,io_writeback_24_bits_vls_vpu_vxrm,2);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_vuopIdx,io_writeback_24_bits_vls_vpu_vuopIdx,7);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_lastUop,io_writeback_24_bits_vls_vpu_lastUop,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_vmask,io_writeback_24_bits_vls_vpu_vmask,128);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_vl,io_writeback_24_bits_vls_vpu_vl,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_nf,io_writeback_24_bits_vls_vpu_nf,3);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_veew,io_writeback_24_bits_vls_vpu_veew,2);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_isReverse,io_writeback_24_bits_vls_vpu_isReverse,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_isExt,io_writeback_24_bits_vls_vpu_isExt,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_isNarrow,io_writeback_24_bits_vls_vpu_isNarrow,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_isDstMask,io_writeback_24_bits_vls_vpu_isDstMask,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_isOpMask,io_writeback_24_bits_vls_vpu_isOpMask,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_isMove,io_writeback_24_bits_vls_vpu_isMove,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_isDependOldVd,io_writeback_24_bits_vls_vpu_isDependOldVd,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_isWritePartVd,io_writeback_24_bits_vls_vpu_isWritePartVd,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vpu_isVleff,io_writeback_24_bits_vls_vpu_isVleff,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_oldVdPsrc,io_writeback_24_bits_vls_oldVdPsrc,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vdIdx,io_writeback_24_bits_vls_vdIdx,3);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_vdIdxInField,io_writeback_24_bits_vls_vdIdxInField,3);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_isIndexed,io_writeback_24_bits_vls_isIndexed,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_isMasked,io_writeback_24_bits_vls_isMasked,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_isStrided,io_writeback_24_bits_vls_isStrided,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_isWhole,io_writeback_24_bits_vls_isWhole,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_isVecLoad,io_writeback_24_bits_vls_isVecLoad,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_vls_isVlm,io_writeback_24_bits_vls_isVlm,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_debug_isMMIO,io_writeback_24_bits_debug_isMMIO,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_debug_isNCIO,io_writeback_24_bits_debug_isNCIO,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_debug_isPerfCnt,io_writeback_24_bits_debug_isPerfCnt,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_debug_paddr,io_writeback_24_bits_debug_paddr,48);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_debug_vaddr,io_writeback_24_bits_debug_vaddr,50);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_debugInfo_eliminatedMove,io_writeback_24_bits_debugInfo_eliminatedMove,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_debugInfo_renameTime,io_writeback_24_bits_debugInfo_renameTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_debugInfo_dispatchTime,io_writeback_24_bits_debugInfo_dispatchTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_debugInfo_enqRsTime,io_writeback_24_bits_debugInfo_enqRsTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_debugInfo_selectTime,io_writeback_24_bits_debugInfo_selectTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_debugInfo_issueTime,io_writeback_24_bits_debugInfo_issueTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_debugInfo_writebackTime,io_writeback_24_bits_debugInfo_writebackTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_debugInfo_runahead_checkpoint_id,io_writeback_24_bits_debugInfo_runahead_checkpoint_id,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_debugInfo_tlbFirstReqTime,io_writeback_24_bits_debugInfo_tlbFirstReqTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_debugInfo_tlbRespTime,io_writeback_24_bits_debugInfo_tlbRespTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_24_bits_debug_seqNum,io_writeback_24_bits_debug_seqNum,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_valid,io_writeback_23_valid,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_data_0,io_writeback_23_bits_data_0,128);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_pdest,io_writeback_23_bits_pdest,7);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_robIdx_flag,io_writeback_23_bits_robIdx_flag,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_robIdx_value,io_writeback_23_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vecWen,io_writeback_23_bits_vecWen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_v0Wen,io_writeback_23_bits_v0Wen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vlWen,io_writeback_23_bits_vlWen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_exceptionVec_0,io_writeback_23_bits_exceptionVec_0,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_exceptionVec_1,io_writeback_23_bits_exceptionVec_1,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_exceptionVec_2,io_writeback_23_bits_exceptionVec_2,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_exceptionVec_3,io_writeback_23_bits_exceptionVec_3,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_exceptionVec_4,io_writeback_23_bits_exceptionVec_4,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_exceptionVec_5,io_writeback_23_bits_exceptionVec_5,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_exceptionVec_6,io_writeback_23_bits_exceptionVec_6,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_exceptionVec_7,io_writeback_23_bits_exceptionVec_7,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_exceptionVec_8,io_writeback_23_bits_exceptionVec_8,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_exceptionVec_9,io_writeback_23_bits_exceptionVec_9,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_exceptionVec_10,io_writeback_23_bits_exceptionVec_10,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_exceptionVec_11,io_writeback_23_bits_exceptionVec_11,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_exceptionVec_12,io_writeback_23_bits_exceptionVec_12,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_exceptionVec_13,io_writeback_23_bits_exceptionVec_13,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_exceptionVec_14,io_writeback_23_bits_exceptionVec_14,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_exceptionVec_15,io_writeback_23_bits_exceptionVec_15,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_exceptionVec_16,io_writeback_23_bits_exceptionVec_16,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_exceptionVec_17,io_writeback_23_bits_exceptionVec_17,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_exceptionVec_18,io_writeback_23_bits_exceptionVec_18,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_exceptionVec_19,io_writeback_23_bits_exceptionVec_19,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_exceptionVec_20,io_writeback_23_bits_exceptionVec_20,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_exceptionVec_21,io_writeback_23_bits_exceptionVec_21,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_exceptionVec_22,io_writeback_23_bits_exceptionVec_22,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_exceptionVec_23,io_writeback_23_bits_exceptionVec_23,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_flushPipe,io_writeback_23_bits_flushPipe,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_replay,io_writeback_23_bits_replay,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_trigger,io_writeback_23_bits_trigger,4);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_vill,io_writeback_23_bits_vls_vpu_vill,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_vma,io_writeback_23_bits_vls_vpu_vma,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_vta,io_writeback_23_bits_vls_vpu_vta,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_vsew,io_writeback_23_bits_vls_vpu_vsew,2);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_vlmul,io_writeback_23_bits_vls_vpu_vlmul,3);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_specVill,io_writeback_23_bits_vls_vpu_specVill,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_specVma,io_writeback_23_bits_vls_vpu_specVma,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_specVta,io_writeback_23_bits_vls_vpu_specVta,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_specVsew,io_writeback_23_bits_vls_vpu_specVsew,2);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_specVlmul,io_writeback_23_bits_vls_vpu_specVlmul,3);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_vm,io_writeback_23_bits_vls_vpu_vm,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_vstart,io_writeback_23_bits_vls_vpu_vstart,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_frm,io_writeback_23_bits_vls_vpu_frm,3);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst,io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_fpu_isFP32Instr,io_writeback_23_bits_vls_vpu_fpu_isFP32Instr,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_fpu_isFP64Instr,io_writeback_23_bits_vls_vpu_fpu_isFP64Instr,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_fpu_isReduction,io_writeback_23_bits_vls_vpu_fpu_isReduction,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2,io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4,io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8,io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_vxrm,io_writeback_23_bits_vls_vpu_vxrm,2);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_vuopIdx,io_writeback_23_bits_vls_vpu_vuopIdx,7);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_lastUop,io_writeback_23_bits_vls_vpu_lastUop,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_vmask,io_writeback_23_bits_vls_vpu_vmask,128);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_vl,io_writeback_23_bits_vls_vpu_vl,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_nf,io_writeback_23_bits_vls_vpu_nf,3);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_veew,io_writeback_23_bits_vls_vpu_veew,2);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_isReverse,io_writeback_23_bits_vls_vpu_isReverse,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_isExt,io_writeback_23_bits_vls_vpu_isExt,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_isNarrow,io_writeback_23_bits_vls_vpu_isNarrow,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_isDstMask,io_writeback_23_bits_vls_vpu_isDstMask,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_isOpMask,io_writeback_23_bits_vls_vpu_isOpMask,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_isMove,io_writeback_23_bits_vls_vpu_isMove,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_isDependOldVd,io_writeback_23_bits_vls_vpu_isDependOldVd,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_isWritePartVd,io_writeback_23_bits_vls_vpu_isWritePartVd,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vpu_isVleff,io_writeback_23_bits_vls_vpu_isVleff,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_oldVdPsrc,io_writeback_23_bits_vls_oldVdPsrc,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vdIdx,io_writeback_23_bits_vls_vdIdx,3);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_vdIdxInField,io_writeback_23_bits_vls_vdIdxInField,3);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_isIndexed,io_writeback_23_bits_vls_isIndexed,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_isMasked,io_writeback_23_bits_vls_isMasked,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_isStrided,io_writeback_23_bits_vls_isStrided,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_isWhole,io_writeback_23_bits_vls_isWhole,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_isVecLoad,io_writeback_23_bits_vls_isVecLoad,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_vls_isVlm,io_writeback_23_bits_vls_isVlm,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_debug_isMMIO,io_writeback_23_bits_debug_isMMIO,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_debug_isNCIO,io_writeback_23_bits_debug_isNCIO,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_debug_isPerfCnt,io_writeback_23_bits_debug_isPerfCnt,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_debug_paddr,io_writeback_23_bits_debug_paddr,48);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_debug_vaddr,io_writeback_23_bits_debug_vaddr,50);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_debugInfo_eliminatedMove,io_writeback_23_bits_debugInfo_eliminatedMove,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_debugInfo_renameTime,io_writeback_23_bits_debugInfo_renameTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_debugInfo_dispatchTime,io_writeback_23_bits_debugInfo_dispatchTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_debugInfo_enqRsTime,io_writeback_23_bits_debugInfo_enqRsTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_debugInfo_selectTime,io_writeback_23_bits_debugInfo_selectTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_debugInfo_issueTime,io_writeback_23_bits_debugInfo_issueTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_debugInfo_writebackTime,io_writeback_23_bits_debugInfo_writebackTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_debugInfo_runahead_checkpoint_id,io_writeback_23_bits_debugInfo_runahead_checkpoint_id,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_debugInfo_tlbFirstReqTime,io_writeback_23_bits_debugInfo_tlbFirstReqTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_debugInfo_tlbRespTime,io_writeback_23_bits_debugInfo_tlbRespTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_23_bits_debug_seqNum,io_writeback_23_bits_debug_seqNum,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_valid,io_writeback_22_valid,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_data_0,io_writeback_22_bits_data_0,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_pdest,io_writeback_22_bits_pdest,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_robIdx_flag,io_writeback_22_bits_robIdx_flag,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_robIdx_value,io_writeback_22_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_intWen,io_writeback_22_bits_intWen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_fpWen,io_writeback_22_bits_fpWen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_exceptionVec_0,io_writeback_22_bits_exceptionVec_0,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_exceptionVec_1,io_writeback_22_bits_exceptionVec_1,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_exceptionVec_2,io_writeback_22_bits_exceptionVec_2,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_exceptionVec_3,io_writeback_22_bits_exceptionVec_3,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_exceptionVec_4,io_writeback_22_bits_exceptionVec_4,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_exceptionVec_5,io_writeback_22_bits_exceptionVec_5,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_exceptionVec_6,io_writeback_22_bits_exceptionVec_6,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_exceptionVec_7,io_writeback_22_bits_exceptionVec_7,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_exceptionVec_8,io_writeback_22_bits_exceptionVec_8,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_exceptionVec_9,io_writeback_22_bits_exceptionVec_9,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_exceptionVec_10,io_writeback_22_bits_exceptionVec_10,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_exceptionVec_11,io_writeback_22_bits_exceptionVec_11,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_exceptionVec_12,io_writeback_22_bits_exceptionVec_12,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_exceptionVec_13,io_writeback_22_bits_exceptionVec_13,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_exceptionVec_14,io_writeback_22_bits_exceptionVec_14,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_exceptionVec_15,io_writeback_22_bits_exceptionVec_15,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_exceptionVec_16,io_writeback_22_bits_exceptionVec_16,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_exceptionVec_17,io_writeback_22_bits_exceptionVec_17,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_exceptionVec_18,io_writeback_22_bits_exceptionVec_18,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_exceptionVec_19,io_writeback_22_bits_exceptionVec_19,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_exceptionVec_20,io_writeback_22_bits_exceptionVec_20,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_exceptionVec_21,io_writeback_22_bits_exceptionVec_21,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_exceptionVec_22,io_writeback_22_bits_exceptionVec_22,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_exceptionVec_23,io_writeback_22_bits_exceptionVec_23,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_flushPipe,io_writeback_22_bits_flushPipe,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_replay,io_writeback_22_bits_replay,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_lqIdx_flag,io_writeback_22_bits_lqIdx_flag,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_lqIdx_value,io_writeback_22_bits_lqIdx_value,7);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_trigger,io_writeback_22_bits_trigger,4);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_predecodeInfo_valid,io_writeback_22_bits_predecodeInfo_valid,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_predecodeInfo_isRVC,io_writeback_22_bits_predecodeInfo_isRVC,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_predecodeInfo_brType,io_writeback_22_bits_predecodeInfo_brType,2);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_predecodeInfo_isCall,io_writeback_22_bits_predecodeInfo_isCall,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_predecodeInfo_isRet,io_writeback_22_bits_predecodeInfo_isRet,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_debug_isMMIO,io_writeback_22_bits_debug_isMMIO,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_debug_isNCIO,io_writeback_22_bits_debug_isNCIO,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_debug_isPerfCnt,io_writeback_22_bits_debug_isPerfCnt,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_debug_paddr,io_writeback_22_bits_debug_paddr,48);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_debug_vaddr,io_writeback_22_bits_debug_vaddr,50);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_debugInfo_eliminatedMove,io_writeback_22_bits_debugInfo_eliminatedMove,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_debugInfo_renameTime,io_writeback_22_bits_debugInfo_renameTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_debugInfo_dispatchTime,io_writeback_22_bits_debugInfo_dispatchTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_debugInfo_enqRsTime,io_writeback_22_bits_debugInfo_enqRsTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_debugInfo_selectTime,io_writeback_22_bits_debugInfo_selectTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_debugInfo_issueTime,io_writeback_22_bits_debugInfo_issueTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_debugInfo_writebackTime,io_writeback_22_bits_debugInfo_writebackTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_debugInfo_runahead_checkpoint_id,io_writeback_22_bits_debugInfo_runahead_checkpoint_id,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_debugInfo_tlbFirstReqTime,io_writeback_22_bits_debugInfo_tlbFirstReqTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_debugInfo_tlbRespTime,io_writeback_22_bits_debugInfo_tlbRespTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_22_bits_debug_seqNum,io_writeback_22_bits_debug_seqNum,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_valid,io_writeback_21_valid,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_data_0,io_writeback_21_bits_data_0,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_pdest,io_writeback_21_bits_pdest,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_robIdx_flag,io_writeback_21_bits_robIdx_flag,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_robIdx_value,io_writeback_21_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_intWen,io_writeback_21_bits_intWen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_fpWen,io_writeback_21_bits_fpWen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_exceptionVec_0,io_writeback_21_bits_exceptionVec_0,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_exceptionVec_1,io_writeback_21_bits_exceptionVec_1,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_exceptionVec_2,io_writeback_21_bits_exceptionVec_2,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_exceptionVec_3,io_writeback_21_bits_exceptionVec_3,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_exceptionVec_4,io_writeback_21_bits_exceptionVec_4,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_exceptionVec_5,io_writeback_21_bits_exceptionVec_5,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_exceptionVec_6,io_writeback_21_bits_exceptionVec_6,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_exceptionVec_7,io_writeback_21_bits_exceptionVec_7,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_exceptionVec_8,io_writeback_21_bits_exceptionVec_8,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_exceptionVec_9,io_writeback_21_bits_exceptionVec_9,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_exceptionVec_10,io_writeback_21_bits_exceptionVec_10,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_exceptionVec_11,io_writeback_21_bits_exceptionVec_11,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_exceptionVec_12,io_writeback_21_bits_exceptionVec_12,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_exceptionVec_13,io_writeback_21_bits_exceptionVec_13,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_exceptionVec_14,io_writeback_21_bits_exceptionVec_14,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_exceptionVec_15,io_writeback_21_bits_exceptionVec_15,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_exceptionVec_16,io_writeback_21_bits_exceptionVec_16,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_exceptionVec_17,io_writeback_21_bits_exceptionVec_17,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_exceptionVec_18,io_writeback_21_bits_exceptionVec_18,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_exceptionVec_19,io_writeback_21_bits_exceptionVec_19,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_exceptionVec_20,io_writeback_21_bits_exceptionVec_20,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_exceptionVec_21,io_writeback_21_bits_exceptionVec_21,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_exceptionVec_22,io_writeback_21_bits_exceptionVec_22,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_exceptionVec_23,io_writeback_21_bits_exceptionVec_23,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_flushPipe,io_writeback_21_bits_flushPipe,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_replay,io_writeback_21_bits_replay,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_lqIdx_flag,io_writeback_21_bits_lqIdx_flag,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_lqIdx_value,io_writeback_21_bits_lqIdx_value,7);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_trigger,io_writeback_21_bits_trigger,4);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_predecodeInfo_valid,io_writeback_21_bits_predecodeInfo_valid,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_predecodeInfo_isRVC,io_writeback_21_bits_predecodeInfo_isRVC,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_predecodeInfo_brType,io_writeback_21_bits_predecodeInfo_brType,2);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_predecodeInfo_isCall,io_writeback_21_bits_predecodeInfo_isCall,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_predecodeInfo_isRet,io_writeback_21_bits_predecodeInfo_isRet,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_debug_isMMIO,io_writeback_21_bits_debug_isMMIO,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_debug_isNCIO,io_writeback_21_bits_debug_isNCIO,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_debug_isPerfCnt,io_writeback_21_bits_debug_isPerfCnt,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_debug_paddr,io_writeback_21_bits_debug_paddr,48);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_debug_vaddr,io_writeback_21_bits_debug_vaddr,50);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_debugInfo_eliminatedMove,io_writeback_21_bits_debugInfo_eliminatedMove,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_debugInfo_renameTime,io_writeback_21_bits_debugInfo_renameTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_debugInfo_dispatchTime,io_writeback_21_bits_debugInfo_dispatchTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_debugInfo_enqRsTime,io_writeback_21_bits_debugInfo_enqRsTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_debugInfo_selectTime,io_writeback_21_bits_debugInfo_selectTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_debugInfo_issueTime,io_writeback_21_bits_debugInfo_issueTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_debugInfo_writebackTime,io_writeback_21_bits_debugInfo_writebackTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_debugInfo_runahead_checkpoint_id,io_writeback_21_bits_debugInfo_runahead_checkpoint_id,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_debugInfo_tlbFirstReqTime,io_writeback_21_bits_debugInfo_tlbFirstReqTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_debugInfo_tlbRespTime,io_writeback_21_bits_debugInfo_tlbRespTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_21_bits_debug_seqNum,io_writeback_21_bits_debug_seqNum,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_valid,io_writeback_20_valid,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_data_0,io_writeback_20_bits_data_0,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_pdest,io_writeback_20_bits_pdest,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_robIdx_flag,io_writeback_20_bits_robIdx_flag,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_robIdx_value,io_writeback_20_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_intWen,io_writeback_20_bits_intWen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_fpWen,io_writeback_20_bits_fpWen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_exceptionVec_0,io_writeback_20_bits_exceptionVec_0,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_exceptionVec_1,io_writeback_20_bits_exceptionVec_1,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_exceptionVec_2,io_writeback_20_bits_exceptionVec_2,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_exceptionVec_3,io_writeback_20_bits_exceptionVec_3,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_exceptionVec_4,io_writeback_20_bits_exceptionVec_4,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_exceptionVec_5,io_writeback_20_bits_exceptionVec_5,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_exceptionVec_6,io_writeback_20_bits_exceptionVec_6,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_exceptionVec_7,io_writeback_20_bits_exceptionVec_7,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_exceptionVec_8,io_writeback_20_bits_exceptionVec_8,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_exceptionVec_9,io_writeback_20_bits_exceptionVec_9,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_exceptionVec_10,io_writeback_20_bits_exceptionVec_10,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_exceptionVec_11,io_writeback_20_bits_exceptionVec_11,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_exceptionVec_12,io_writeback_20_bits_exceptionVec_12,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_exceptionVec_13,io_writeback_20_bits_exceptionVec_13,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_exceptionVec_14,io_writeback_20_bits_exceptionVec_14,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_exceptionVec_15,io_writeback_20_bits_exceptionVec_15,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_exceptionVec_16,io_writeback_20_bits_exceptionVec_16,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_exceptionVec_17,io_writeback_20_bits_exceptionVec_17,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_exceptionVec_18,io_writeback_20_bits_exceptionVec_18,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_exceptionVec_19,io_writeback_20_bits_exceptionVec_19,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_exceptionVec_20,io_writeback_20_bits_exceptionVec_20,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_exceptionVec_21,io_writeback_20_bits_exceptionVec_21,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_exceptionVec_22,io_writeback_20_bits_exceptionVec_22,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_exceptionVec_23,io_writeback_20_bits_exceptionVec_23,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_flushPipe,io_writeback_20_bits_flushPipe,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_replay,io_writeback_20_bits_replay,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_lqIdx_flag,io_writeback_20_bits_lqIdx_flag,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_lqIdx_value,io_writeback_20_bits_lqIdx_value,7);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_trigger,io_writeback_20_bits_trigger,4);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_predecodeInfo_valid,io_writeback_20_bits_predecodeInfo_valid,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_predecodeInfo_isRVC,io_writeback_20_bits_predecodeInfo_isRVC,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_predecodeInfo_brType,io_writeback_20_bits_predecodeInfo_brType,2);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_predecodeInfo_isCall,io_writeback_20_bits_predecodeInfo_isCall,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_predecodeInfo_isRet,io_writeback_20_bits_predecodeInfo_isRet,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_debug_isMMIO,io_writeback_20_bits_debug_isMMIO,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_debug_isNCIO,io_writeback_20_bits_debug_isNCIO,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_debug_isPerfCnt,io_writeback_20_bits_debug_isPerfCnt,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_debug_paddr,io_writeback_20_bits_debug_paddr,48);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_debug_vaddr,io_writeback_20_bits_debug_vaddr,50);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_debugInfo_eliminatedMove,io_writeback_20_bits_debugInfo_eliminatedMove,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_debugInfo_renameTime,io_writeback_20_bits_debugInfo_renameTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_debugInfo_dispatchTime,io_writeback_20_bits_debugInfo_dispatchTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_debugInfo_enqRsTime,io_writeback_20_bits_debugInfo_enqRsTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_debugInfo_selectTime,io_writeback_20_bits_debugInfo_selectTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_debugInfo_issueTime,io_writeback_20_bits_debugInfo_issueTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_debugInfo_writebackTime,io_writeback_20_bits_debugInfo_writebackTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_debugInfo_runahead_checkpoint_id,io_writeback_20_bits_debugInfo_runahead_checkpoint_id,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_debugInfo_tlbFirstReqTime,io_writeback_20_bits_debugInfo_tlbFirstReqTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_debugInfo_tlbRespTime,io_writeback_20_bits_debugInfo_tlbRespTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_20_bits_debug_seqNum,io_writeback_20_bits_debug_seqNum,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_valid,io_writeback_19_valid,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_data_0,io_writeback_19_bits_data_0,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_pdest,io_writeback_19_bits_pdest,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_robIdx_flag,io_writeback_19_bits_robIdx_flag,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_robIdx_value,io_writeback_19_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_intWen,io_writeback_19_bits_intWen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_exceptionVec_0,io_writeback_19_bits_exceptionVec_0,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_exceptionVec_1,io_writeback_19_bits_exceptionVec_1,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_exceptionVec_2,io_writeback_19_bits_exceptionVec_2,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_exceptionVec_3,io_writeback_19_bits_exceptionVec_3,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_exceptionVec_4,io_writeback_19_bits_exceptionVec_4,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_exceptionVec_5,io_writeback_19_bits_exceptionVec_5,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_exceptionVec_6,io_writeback_19_bits_exceptionVec_6,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_exceptionVec_7,io_writeback_19_bits_exceptionVec_7,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_exceptionVec_8,io_writeback_19_bits_exceptionVec_8,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_exceptionVec_9,io_writeback_19_bits_exceptionVec_9,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_exceptionVec_10,io_writeback_19_bits_exceptionVec_10,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_exceptionVec_11,io_writeback_19_bits_exceptionVec_11,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_exceptionVec_12,io_writeback_19_bits_exceptionVec_12,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_exceptionVec_13,io_writeback_19_bits_exceptionVec_13,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_exceptionVec_14,io_writeback_19_bits_exceptionVec_14,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_exceptionVec_15,io_writeback_19_bits_exceptionVec_15,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_exceptionVec_16,io_writeback_19_bits_exceptionVec_16,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_exceptionVec_17,io_writeback_19_bits_exceptionVec_17,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_exceptionVec_18,io_writeback_19_bits_exceptionVec_18,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_exceptionVec_19,io_writeback_19_bits_exceptionVec_19,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_exceptionVec_20,io_writeback_19_bits_exceptionVec_20,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_exceptionVec_21,io_writeback_19_bits_exceptionVec_21,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_exceptionVec_22,io_writeback_19_bits_exceptionVec_22,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_exceptionVec_23,io_writeback_19_bits_exceptionVec_23,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_flushPipe,io_writeback_19_bits_flushPipe,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_sqIdx_flag,io_writeback_19_bits_sqIdx_flag,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_sqIdx_value,io_writeback_19_bits_sqIdx_value,6);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_trigger,io_writeback_19_bits_trigger,4);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_debug_isMMIO,io_writeback_19_bits_debug_isMMIO,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_debug_isNCIO,io_writeback_19_bits_debug_isNCIO,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_debug_isPerfCnt,io_writeback_19_bits_debug_isPerfCnt,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_debug_paddr,io_writeback_19_bits_debug_paddr,48);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_debug_vaddr,io_writeback_19_bits_debug_vaddr,50);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_debugInfo_eliminatedMove,io_writeback_19_bits_debugInfo_eliminatedMove,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_debugInfo_renameTime,io_writeback_19_bits_debugInfo_renameTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_debugInfo_dispatchTime,io_writeback_19_bits_debugInfo_dispatchTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_debugInfo_enqRsTime,io_writeback_19_bits_debugInfo_enqRsTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_debugInfo_selectTime,io_writeback_19_bits_debugInfo_selectTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_debugInfo_issueTime,io_writeback_19_bits_debugInfo_issueTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_debugInfo_writebackTime,io_writeback_19_bits_debugInfo_writebackTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_debugInfo_runahead_checkpoint_id,io_writeback_19_bits_debugInfo_runahead_checkpoint_id,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_debugInfo_tlbFirstReqTime,io_writeback_19_bits_debugInfo_tlbFirstReqTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_debugInfo_tlbRespTime,io_writeback_19_bits_debugInfo_tlbRespTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_19_bits_debug_seqNum,io_writeback_19_bits_debug_seqNum,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_valid,io_writeback_18_valid,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_data_0,io_writeback_18_bits_data_0,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_pdest,io_writeback_18_bits_pdest,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_robIdx_flag,io_writeback_18_bits_robIdx_flag,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_robIdx_value,io_writeback_18_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_intWen,io_writeback_18_bits_intWen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_exceptionVec_0,io_writeback_18_bits_exceptionVec_0,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_exceptionVec_1,io_writeback_18_bits_exceptionVec_1,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_exceptionVec_2,io_writeback_18_bits_exceptionVec_2,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_exceptionVec_3,io_writeback_18_bits_exceptionVec_3,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_exceptionVec_4,io_writeback_18_bits_exceptionVec_4,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_exceptionVec_5,io_writeback_18_bits_exceptionVec_5,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_exceptionVec_6,io_writeback_18_bits_exceptionVec_6,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_exceptionVec_7,io_writeback_18_bits_exceptionVec_7,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_exceptionVec_8,io_writeback_18_bits_exceptionVec_8,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_exceptionVec_9,io_writeback_18_bits_exceptionVec_9,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_exceptionVec_10,io_writeback_18_bits_exceptionVec_10,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_exceptionVec_11,io_writeback_18_bits_exceptionVec_11,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_exceptionVec_12,io_writeback_18_bits_exceptionVec_12,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_exceptionVec_13,io_writeback_18_bits_exceptionVec_13,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_exceptionVec_14,io_writeback_18_bits_exceptionVec_14,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_exceptionVec_15,io_writeback_18_bits_exceptionVec_15,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_exceptionVec_16,io_writeback_18_bits_exceptionVec_16,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_exceptionVec_17,io_writeback_18_bits_exceptionVec_17,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_exceptionVec_18,io_writeback_18_bits_exceptionVec_18,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_exceptionVec_19,io_writeback_18_bits_exceptionVec_19,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_exceptionVec_20,io_writeback_18_bits_exceptionVec_20,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_exceptionVec_21,io_writeback_18_bits_exceptionVec_21,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_exceptionVec_22,io_writeback_18_bits_exceptionVec_22,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_exceptionVec_23,io_writeback_18_bits_exceptionVec_23,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_flushPipe,io_writeback_18_bits_flushPipe,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_sqIdx_flag,io_writeback_18_bits_sqIdx_flag,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_sqIdx_value,io_writeback_18_bits_sqIdx_value,6);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_trigger,io_writeback_18_bits_trigger,4);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_debug_isMMIO,io_writeback_18_bits_debug_isMMIO,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_debug_isNCIO,io_writeback_18_bits_debug_isNCIO,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_debug_isPerfCnt,io_writeback_18_bits_debug_isPerfCnt,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_debug_paddr,io_writeback_18_bits_debug_paddr,48);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_debug_vaddr,io_writeback_18_bits_debug_vaddr,50);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_debugInfo_eliminatedMove,io_writeback_18_bits_debugInfo_eliminatedMove,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_debugInfo_renameTime,io_writeback_18_bits_debugInfo_renameTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_debugInfo_dispatchTime,io_writeback_18_bits_debugInfo_dispatchTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_debugInfo_enqRsTime,io_writeback_18_bits_debugInfo_enqRsTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_debugInfo_selectTime,io_writeback_18_bits_debugInfo_selectTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_debugInfo_issueTime,io_writeback_18_bits_debugInfo_issueTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_debugInfo_writebackTime,io_writeback_18_bits_debugInfo_writebackTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_debugInfo_runahead_checkpoint_id,io_writeback_18_bits_debugInfo_runahead_checkpoint_id,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_debugInfo_tlbFirstReqTime,io_writeback_18_bits_debugInfo_tlbFirstReqTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_debugInfo_tlbRespTime,io_writeback_18_bits_debugInfo_tlbRespTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_18_bits_debug_seqNum,io_writeback_18_bits_debug_seqNum,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_17_valid,io_writeback_17_valid,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_17_bits_data_0,io_writeback_17_bits_data_0,128);
            `TCNT_CHECK_SIG_XZ(io_writeback_17_bits_data_1,io_writeback_17_bits_data_1,128);
            `TCNT_CHECK_SIG_XZ(io_writeback_17_bits_data_2,io_writeback_17_bits_data_2,128);
            `TCNT_CHECK_SIG_XZ(io_writeback_17_bits_pdest,io_writeback_17_bits_pdest,7);
            `TCNT_CHECK_SIG_XZ(io_writeback_17_bits_robIdx_flag,io_writeback_17_bits_robIdx_flag,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_17_bits_robIdx_value,io_writeback_17_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_17_bits_vecWen,io_writeback_17_bits_vecWen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_17_bits_v0Wen,io_writeback_17_bits_v0Wen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_17_bits_fflags,io_writeback_17_bits_fflags,5);
            `TCNT_CHECK_SIG_XZ(io_writeback_17_bits_wflags,io_writeback_17_bits_wflags,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_17_bits_debugInfo_eliminatedMove,io_writeback_17_bits_debugInfo_eliminatedMove,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_17_bits_debugInfo_renameTime,io_writeback_17_bits_debugInfo_renameTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_17_bits_debugInfo_dispatchTime,io_writeback_17_bits_debugInfo_dispatchTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_17_bits_debugInfo_enqRsTime,io_writeback_17_bits_debugInfo_enqRsTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_17_bits_debugInfo_selectTime,io_writeback_17_bits_debugInfo_selectTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_17_bits_debugInfo_issueTime,io_writeback_17_bits_debugInfo_issueTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_17_bits_debugInfo_writebackTime,io_writeback_17_bits_debugInfo_writebackTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_17_bits_debugInfo_runahead_checkpoint_id,io_writeback_17_bits_debugInfo_runahead_checkpoint_id,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_17_bits_debugInfo_tlbFirstReqTime,io_writeback_17_bits_debugInfo_tlbFirstReqTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_17_bits_debugInfo_tlbRespTime,io_writeback_17_bits_debugInfo_tlbRespTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_17_bits_debug_seqNum,io_writeback_17_bits_debug_seqNum,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_16_valid,io_writeback_16_valid,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_16_bits_data_0,io_writeback_16_bits_data_0,128);
            `TCNT_CHECK_SIG_XZ(io_writeback_16_bits_data_1,io_writeback_16_bits_data_1,128);
            `TCNT_CHECK_SIG_XZ(io_writeback_16_bits_data_2,io_writeback_16_bits_data_2,128);
            `TCNT_CHECK_SIG_XZ(io_writeback_16_bits_data_3,io_writeback_16_bits_data_3,128);
            `TCNT_CHECK_SIG_XZ(io_writeback_16_bits_pdest,io_writeback_16_bits_pdest,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_16_bits_robIdx_flag,io_writeback_16_bits_robIdx_flag,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_16_bits_robIdx_value,io_writeback_16_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_16_bits_fpWen,io_writeback_16_bits_fpWen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_16_bits_vecWen,io_writeback_16_bits_vecWen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_16_bits_v0Wen,io_writeback_16_bits_v0Wen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_16_bits_fflags,io_writeback_16_bits_fflags,5);
            `TCNT_CHECK_SIG_XZ(io_writeback_16_bits_wflags,io_writeback_16_bits_wflags,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_16_bits_debugInfo_eliminatedMove,io_writeback_16_bits_debugInfo_eliminatedMove,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_16_bits_debugInfo_renameTime,io_writeback_16_bits_debugInfo_renameTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_16_bits_debugInfo_dispatchTime,io_writeback_16_bits_debugInfo_dispatchTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_16_bits_debugInfo_enqRsTime,io_writeback_16_bits_debugInfo_enqRsTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_16_bits_debugInfo_selectTime,io_writeback_16_bits_debugInfo_selectTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_16_bits_debugInfo_issueTime,io_writeback_16_bits_debugInfo_issueTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_16_bits_debugInfo_writebackTime,io_writeback_16_bits_debugInfo_writebackTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_16_bits_debugInfo_runahead_checkpoint_id,io_writeback_16_bits_debugInfo_runahead_checkpoint_id,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_16_bits_debugInfo_tlbFirstReqTime,io_writeback_16_bits_debugInfo_tlbFirstReqTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_16_bits_debugInfo_tlbRespTime,io_writeback_16_bits_debugInfo_tlbRespTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_16_bits_debug_seqNum,io_writeback_16_bits_debug_seqNum,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_15_valid,io_writeback_15_valid,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_15_bits_data_0,io_writeback_15_bits_data_0,128);
            `TCNT_CHECK_SIG_XZ(io_writeback_15_bits_data_1,io_writeback_15_bits_data_1,128);
            `TCNT_CHECK_SIG_XZ(io_writeback_15_bits_data_2,io_writeback_15_bits_data_2,128);
            `TCNT_CHECK_SIG_XZ(io_writeback_15_bits_pdest,io_writeback_15_bits_pdest,7);
            `TCNT_CHECK_SIG_XZ(io_writeback_15_bits_robIdx_flag,io_writeback_15_bits_robIdx_flag,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_15_bits_robIdx_value,io_writeback_15_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_15_bits_vecWen,io_writeback_15_bits_vecWen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_15_bits_v0Wen,io_writeback_15_bits_v0Wen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_15_bits_fflags,io_writeback_15_bits_fflags,5);
            `TCNT_CHECK_SIG_XZ(io_writeback_15_bits_wflags,io_writeback_15_bits_wflags,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_15_bits_vxsat,io_writeback_15_bits_vxsat,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_15_bits_debugInfo_eliminatedMove,io_writeback_15_bits_debugInfo_eliminatedMove,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_15_bits_debugInfo_renameTime,io_writeback_15_bits_debugInfo_renameTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_15_bits_debugInfo_dispatchTime,io_writeback_15_bits_debugInfo_dispatchTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_15_bits_debugInfo_enqRsTime,io_writeback_15_bits_debugInfo_enqRsTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_15_bits_debugInfo_selectTime,io_writeback_15_bits_debugInfo_selectTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_15_bits_debugInfo_issueTime,io_writeback_15_bits_debugInfo_issueTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_15_bits_debugInfo_writebackTime,io_writeback_15_bits_debugInfo_writebackTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_15_bits_debugInfo_runahead_checkpoint_id,io_writeback_15_bits_debugInfo_runahead_checkpoint_id,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_15_bits_debugInfo_tlbFirstReqTime,io_writeback_15_bits_debugInfo_tlbFirstReqTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_15_bits_debugInfo_tlbRespTime,io_writeback_15_bits_debugInfo_tlbRespTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_15_bits_debug_seqNum,io_writeback_15_bits_debug_seqNum,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_valid,io_writeback_14_valid,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_bits_data_0,io_writeback_14_bits_data_0,128);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_bits_data_1,io_writeback_14_bits_data_1,128);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_bits_data_2,io_writeback_14_bits_data_2,128);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_bits_data_3,io_writeback_14_bits_data_3,128);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_bits_data_4,io_writeback_14_bits_data_4,128);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_bits_data_5,io_writeback_14_bits_data_5,128);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_bits_pdest,io_writeback_14_bits_pdest,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_bits_robIdx_flag,io_writeback_14_bits_robIdx_flag,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_bits_robIdx_value,io_writeback_14_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_bits_intWen,io_writeback_14_bits_intWen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_bits_fpWen,io_writeback_14_bits_fpWen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_bits_vecWen,io_writeback_14_bits_vecWen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_bits_v0Wen,io_writeback_14_bits_v0Wen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_bits_vlWen,io_writeback_14_bits_vlWen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_bits_fflags,io_writeback_14_bits_fflags,5);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_bits_wflags,io_writeback_14_bits_wflags,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_bits_exceptionVec_2,io_writeback_14_bits_exceptionVec_2,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_bits_debugInfo_eliminatedMove,io_writeback_14_bits_debugInfo_eliminatedMove,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_bits_debugInfo_renameTime,io_writeback_14_bits_debugInfo_renameTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_bits_debugInfo_dispatchTime,io_writeback_14_bits_debugInfo_dispatchTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_bits_debugInfo_enqRsTime,io_writeback_14_bits_debugInfo_enqRsTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_bits_debugInfo_selectTime,io_writeback_14_bits_debugInfo_selectTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_bits_debugInfo_issueTime,io_writeback_14_bits_debugInfo_issueTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_bits_debugInfo_writebackTime,io_writeback_14_bits_debugInfo_writebackTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_bits_debugInfo_runahead_checkpoint_id,io_writeback_14_bits_debugInfo_runahead_checkpoint_id,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_bits_debugInfo_tlbFirstReqTime,io_writeback_14_bits_debugInfo_tlbFirstReqTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_bits_debugInfo_tlbRespTime,io_writeback_14_bits_debugInfo_tlbRespTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_14_bits_debug_seqNum,io_writeback_14_bits_debug_seqNum,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_13_valid,io_writeback_13_valid,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_13_bits_data_0,io_writeback_13_bits_data_0,128);
            `TCNT_CHECK_SIG_XZ(io_writeback_13_bits_data_1,io_writeback_13_bits_data_1,128);
            `TCNT_CHECK_SIG_XZ(io_writeback_13_bits_data_2,io_writeback_13_bits_data_2,128);
            `TCNT_CHECK_SIG_XZ(io_writeback_13_bits_pdest,io_writeback_13_bits_pdest,7);
            `TCNT_CHECK_SIG_XZ(io_writeback_13_bits_robIdx_flag,io_writeback_13_bits_robIdx_flag,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_13_bits_robIdx_value,io_writeback_13_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_13_bits_vecWen,io_writeback_13_bits_vecWen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_13_bits_v0Wen,io_writeback_13_bits_v0Wen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_13_bits_fflags,io_writeback_13_bits_fflags,5);
            `TCNT_CHECK_SIG_XZ(io_writeback_13_bits_wflags,io_writeback_13_bits_wflags,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_13_bits_vxsat,io_writeback_13_bits_vxsat,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_13_bits_exceptionVec_2,io_writeback_13_bits_exceptionVec_2,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_13_bits_debugInfo_eliminatedMove,io_writeback_13_bits_debugInfo_eliminatedMove,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_13_bits_debugInfo_renameTime,io_writeback_13_bits_debugInfo_renameTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_13_bits_debugInfo_dispatchTime,io_writeback_13_bits_debugInfo_dispatchTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_13_bits_debugInfo_enqRsTime,io_writeback_13_bits_debugInfo_enqRsTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_13_bits_debugInfo_selectTime,io_writeback_13_bits_debugInfo_selectTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_13_bits_debugInfo_issueTime,io_writeback_13_bits_debugInfo_issueTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_13_bits_debugInfo_writebackTime,io_writeback_13_bits_debugInfo_writebackTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_13_bits_debugInfo_runahead_checkpoint_id,io_writeback_13_bits_debugInfo_runahead_checkpoint_id,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_13_bits_debugInfo_tlbFirstReqTime,io_writeback_13_bits_debugInfo_tlbFirstReqTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_13_bits_debugInfo_tlbRespTime,io_writeback_13_bits_debugInfo_tlbRespTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_13_bits_debug_seqNum,io_writeback_13_bits_debug_seqNum,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_valid,io_writeback_7_valid,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_data_0,io_writeback_7_bits_data_0,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_data_1,io_writeback_7_bits_data_1,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_pdest,io_writeback_7_bits_pdest,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_robIdx_flag,io_writeback_7_bits_robIdx_flag,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_robIdx_value,io_writeback_7_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_intWen,io_writeback_7_bits_intWen,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_valid,io_writeback_7_bits_redirect_valid,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_isRVC,io_writeback_7_bits_redirect_bits_isRVC,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_robIdx_flag,io_writeback_7_bits_redirect_bits_robIdx_flag,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_robIdx_value,io_writeback_7_bits_redirect_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_ftqIdx_flag,io_writeback_7_bits_redirect_bits_ftqIdx_flag,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_ftqIdx_value,io_writeback_7_bits_redirect_bits_ftqIdx_value,6);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_ftqOffset,io_writeback_7_bits_redirect_bits_ftqOffset,4);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_level,io_writeback_7_bits_redirect_bits_level,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_interrupt,io_writeback_7_bits_redirect_bits_interrupt,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_pc,io_writeback_7_bits_redirect_bits_cfiUpdate_pc,50);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid,io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC,io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType,io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType,2);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall,io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet,io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_ssp,io_writeback_7_bits_redirect_bits_cfiUpdate_ssp,4);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_sctr,io_writeback_7_bits_redirect_bits_cfiUpdate_sctr,3);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag,io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value,io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value,5);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag,io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value,io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value,5);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag,io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value,io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value,5);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr,io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr,50);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist,io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist,11);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist,io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist,11);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist,io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist,7);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist,io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist,io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist,9);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist,io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist,4);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist,io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist,io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist,9);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist,io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist,7);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist,io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist,io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist,7);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist,io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist,9);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist,io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist,7);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist,io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist,io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist,io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist,io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist,11);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist,io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0,io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1,io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2,io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3,io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0,io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1,io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2,io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3,io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0,io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1,io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2,io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3,io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0,io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1,io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2,io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3,io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0,io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1,io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2,io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3,io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0,io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1,io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2,io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3,io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH,io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH,3);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_ghr,io_writeback_7_bits_redirect_bits_cfiUpdate_ghr,4);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag,io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value,io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value,8);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0,io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0,10);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1,io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1,10);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit,io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit,io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit,io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken,io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_target,io_writeback_7_bits_redirect_bits_cfiUpdate_target,50);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_taken,io_writeback_7_bits_redirect_bits_cfiUpdate_taken,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred,io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_shift,io_writeback_7_bits_redirect_bits_cfiUpdate_shift,2);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist,io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF,io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF,io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF,io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_fullTarget,io_writeback_7_bits_redirect_bits_fullTarget,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_stFtqIdx_flag,io_writeback_7_bits_redirect_bits_stFtqIdx_flag,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_stFtqIdx_value,io_writeback_7_bits_redirect_bits_stFtqIdx_value,6);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_stFtqOffset,io_writeback_7_bits_redirect_bits_stFtqOffset,4);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id,io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_debugIsCtrl,io_writeback_7_bits_redirect_bits_debugIsCtrl,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_redirect_bits_debugIsMemVio,io_writeback_7_bits_redirect_bits_debugIsMemVio,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_exceptionVec_2,io_writeback_7_bits_exceptionVec_2,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_exceptionVec_3,io_writeback_7_bits_exceptionVec_3,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_exceptionVec_8,io_writeback_7_bits_exceptionVec_8,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_exceptionVec_9,io_writeback_7_bits_exceptionVec_9,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_exceptionVec_10,io_writeback_7_bits_exceptionVec_10,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_exceptionVec_11,io_writeback_7_bits_exceptionVec_11,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_exceptionVec_22,io_writeback_7_bits_exceptionVec_22,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_flushPipe,io_writeback_7_bits_flushPipe,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_predecodeInfo_valid,io_writeback_7_bits_predecodeInfo_valid,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_predecodeInfo_isRVC,io_writeback_7_bits_predecodeInfo_isRVC,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_predecodeInfo_brType,io_writeback_7_bits_predecodeInfo_brType,2);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_predecodeInfo_isCall,io_writeback_7_bits_predecodeInfo_isCall,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_predecodeInfo_isRet,io_writeback_7_bits_predecodeInfo_isRet,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_debug_isPerfCnt,io_writeback_7_bits_debug_isPerfCnt,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_debugInfo_eliminatedMove,io_writeback_7_bits_debugInfo_eliminatedMove,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_debugInfo_renameTime,io_writeback_7_bits_debugInfo_renameTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_debugInfo_dispatchTime,io_writeback_7_bits_debugInfo_dispatchTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_debugInfo_enqRsTime,io_writeback_7_bits_debugInfo_enqRsTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_debugInfo_selectTime,io_writeback_7_bits_debugInfo_selectTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_debugInfo_issueTime,io_writeback_7_bits_debugInfo_issueTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_debugInfo_writebackTime,io_writeback_7_bits_debugInfo_writebackTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_debugInfo_runahead_checkpoint_id,io_writeback_7_bits_debugInfo_runahead_checkpoint_id,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_debugInfo_tlbFirstReqTime,io_writeback_7_bits_debugInfo_tlbFirstReqTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_debugInfo_tlbRespTime,io_writeback_7_bits_debugInfo_tlbRespTime,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_7_bits_debug_seqNum,io_writeback_7_bits_debug_seqNum,64);
            `TCNT_CHECK_SIG_XZ(io_writeback_5_valid,io_writeback_5_valid,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_5_bits_redirect_valid,io_writeback_5_bits_redirect_valid,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred,io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_3_valid,io_writeback_3_valid,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_3_bits_redirect_valid,io_writeback_3_bits_redirect_valid,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred,io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_1_valid,io_writeback_1_valid,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_1_bits_redirect_valid,io_writeback_1_bits_redirect_valid,1);
            `TCNT_CHECK_SIG_XZ(io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred,io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_26_valid,io_exuWriteback_26_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_26_bits_robIdx_value,io_exuWriteback_26_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_25_valid,io_exuWriteback_25_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_25_bits_robIdx_value,io_exuWriteback_25_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_24_valid,io_exuWriteback_24_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_24_bits_data_0,io_exuWriteback_24_bits_data_0,128);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_24_bits_pdest,io_exuWriteback_24_bits_pdest,7);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_24_bits_robIdx_value,io_exuWriteback_24_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_24_bits_vecWen,io_exuWriteback_24_bits_vecWen,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_24_bits_v0Wen,io_exuWriteback_24_bits_v0Wen,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_24_bits_vls_vdIdx,io_exuWriteback_24_bits_vls_vdIdx,3);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_24_bits_debug_isMMIO,io_exuWriteback_24_bits_debug_isMMIO,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_24_bits_debug_isNCIO,io_exuWriteback_24_bits_debug_isNCIO,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_24_bits_debug_isPerfCnt,io_exuWriteback_24_bits_debug_isPerfCnt,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_24_bits_debug_paddr,io_exuWriteback_24_bits_debug_paddr,48);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_23_valid,io_exuWriteback_23_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_23_bits_data_0,io_exuWriteback_23_bits_data_0,128);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_23_bits_pdest,io_exuWriteback_23_bits_pdest,7);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_23_bits_robIdx_value,io_exuWriteback_23_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_23_bits_vecWen,io_exuWriteback_23_bits_vecWen,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_23_bits_v0Wen,io_exuWriteback_23_bits_v0Wen,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_23_bits_vls_vdIdx,io_exuWriteback_23_bits_vls_vdIdx,3);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_23_bits_debug_isMMIO,io_exuWriteback_23_bits_debug_isMMIO,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_23_bits_debug_isNCIO,io_exuWriteback_23_bits_debug_isNCIO,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_23_bits_debug_isPerfCnt,io_exuWriteback_23_bits_debug_isPerfCnt,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_23_bits_debug_paddr,io_exuWriteback_23_bits_debug_paddr,48);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_22_valid,io_exuWriteback_22_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_22_bits_data_0,io_exuWriteback_22_bits_data_0,64);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_22_bits_robIdx_value,io_exuWriteback_22_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_22_bits_lqIdx_value,io_exuWriteback_22_bits_lqIdx_value,7);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_22_bits_debug_isMMIO,io_exuWriteback_22_bits_debug_isMMIO,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_22_bits_debug_isNCIO,io_exuWriteback_22_bits_debug_isNCIO,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_22_bits_debug_isPerfCnt,io_exuWriteback_22_bits_debug_isPerfCnt,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_22_bits_debug_paddr,io_exuWriteback_22_bits_debug_paddr,48);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_21_valid,io_exuWriteback_21_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_21_bits_data_0,io_exuWriteback_21_bits_data_0,64);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_21_bits_robIdx_value,io_exuWriteback_21_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_21_bits_lqIdx_value,io_exuWriteback_21_bits_lqIdx_value,7);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_21_bits_debug_isMMIO,io_exuWriteback_21_bits_debug_isMMIO,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_21_bits_debug_isNCIO,io_exuWriteback_21_bits_debug_isNCIO,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_21_bits_debug_isPerfCnt,io_exuWriteback_21_bits_debug_isPerfCnt,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_21_bits_debug_paddr,io_exuWriteback_21_bits_debug_paddr,48);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_20_valid,io_exuWriteback_20_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_20_bits_data_0,io_exuWriteback_20_bits_data_0,64);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_20_bits_robIdx_value,io_exuWriteback_20_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_20_bits_lqIdx_value,io_exuWriteback_20_bits_lqIdx_value,7);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_20_bits_debug_isMMIO,io_exuWriteback_20_bits_debug_isMMIO,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_20_bits_debug_isNCIO,io_exuWriteback_20_bits_debug_isNCIO,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_20_bits_debug_isPerfCnt,io_exuWriteback_20_bits_debug_isPerfCnt,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_20_bits_debug_paddr,io_exuWriteback_20_bits_debug_paddr,48);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_19_valid,io_exuWriteback_19_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_19_bits_data_0,io_exuWriteback_19_bits_data_0,64);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_19_bits_robIdx_value,io_exuWriteback_19_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_19_bits_sqIdx_value,io_exuWriteback_19_bits_sqIdx_value,6);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_19_bits_debug_isMMIO,io_exuWriteback_19_bits_debug_isMMIO,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_19_bits_debug_isNCIO,io_exuWriteback_19_bits_debug_isNCIO,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_19_bits_debug_isPerfCnt,io_exuWriteback_19_bits_debug_isPerfCnt,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_19_bits_debug_paddr,io_exuWriteback_19_bits_debug_paddr,48);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_18_valid,io_exuWriteback_18_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_18_bits_data_0,io_exuWriteback_18_bits_data_0,64);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_18_bits_robIdx_value,io_exuWriteback_18_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_18_bits_sqIdx_value,io_exuWriteback_18_bits_sqIdx_value,6);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_18_bits_debug_isMMIO,io_exuWriteback_18_bits_debug_isMMIO,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_18_bits_debug_isNCIO,io_exuWriteback_18_bits_debug_isNCIO,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_18_bits_debug_isPerfCnt,io_exuWriteback_18_bits_debug_isPerfCnt,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_18_bits_debug_paddr,io_exuWriteback_18_bits_debug_paddr,48);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_17_valid,io_exuWriteback_17_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_17_bits_data_0,io_exuWriteback_17_bits_data_0,128);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_17_bits_robIdx_value,io_exuWriteback_17_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_17_bits_fflags,io_exuWriteback_17_bits_fflags,5);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_17_bits_wflags,io_exuWriteback_17_bits_wflags,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_16_valid,io_exuWriteback_16_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_16_bits_data_0,io_exuWriteback_16_bits_data_0,128);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_16_bits_robIdx_value,io_exuWriteback_16_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_16_bits_fflags,io_exuWriteback_16_bits_fflags,5);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_16_bits_wflags,io_exuWriteback_16_bits_wflags,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_15_valid,io_exuWriteback_15_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_15_bits_data_0,io_exuWriteback_15_bits_data_0,128);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_15_bits_robIdx_value,io_exuWriteback_15_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_15_bits_fflags,io_exuWriteback_15_bits_fflags,5);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_15_bits_wflags,io_exuWriteback_15_bits_wflags,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_15_bits_vxsat,io_exuWriteback_15_bits_vxsat,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_14_valid,io_exuWriteback_14_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_14_bits_data_0,io_exuWriteback_14_bits_data_0,128);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_14_bits_robIdx_value,io_exuWriteback_14_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_14_bits_fflags,io_exuWriteback_14_bits_fflags,5);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_14_bits_wflags,io_exuWriteback_14_bits_wflags,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_13_valid,io_exuWriteback_13_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_13_bits_data_0,io_exuWriteback_13_bits_data_0,128);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_13_bits_robIdx_value,io_exuWriteback_13_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_13_bits_fflags,io_exuWriteback_13_bits_fflags,5);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_13_bits_wflags,io_exuWriteback_13_bits_wflags,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_13_bits_vxsat,io_exuWriteback_13_bits_vxsat,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_12_valid,io_exuWriteback_12_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_12_bits_data_0,io_exuWriteback_12_bits_data_0,64);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_12_bits_robIdx_value,io_exuWriteback_12_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_12_bits_fflags,io_exuWriteback_12_bits_fflags,5);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_12_bits_wflags,io_exuWriteback_12_bits_wflags,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_11_valid,io_exuWriteback_11_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_11_bits_data_0,io_exuWriteback_11_bits_data_0,64);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_11_bits_robIdx_value,io_exuWriteback_11_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_11_bits_fflags,io_exuWriteback_11_bits_fflags,5);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_11_bits_wflags,io_exuWriteback_11_bits_wflags,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_10_valid,io_exuWriteback_10_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_10_bits_data_0,io_exuWriteback_10_bits_data_0,64);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_10_bits_robIdx_value,io_exuWriteback_10_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_10_bits_fflags,io_exuWriteback_10_bits_fflags,5);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_10_bits_wflags,io_exuWriteback_10_bits_wflags,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_9_valid,io_exuWriteback_9_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_9_bits_data_0,io_exuWriteback_9_bits_data_0,64);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_9_bits_robIdx_value,io_exuWriteback_9_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_9_bits_fflags,io_exuWriteback_9_bits_fflags,5);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_9_bits_wflags,io_exuWriteback_9_bits_wflags,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_8_valid,io_exuWriteback_8_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_8_bits_data_0,io_exuWriteback_8_bits_data_0,128);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_8_bits_robIdx_value,io_exuWriteback_8_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_8_bits_fflags,io_exuWriteback_8_bits_fflags,5);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_8_bits_wflags,io_exuWriteback_8_bits_wflags,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_7_valid,io_exuWriteback_7_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_7_bits_data_0,io_exuWriteback_7_bits_data_0,64);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_7_bits_robIdx_value,io_exuWriteback_7_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_7_bits_debug_isPerfCnt,io_exuWriteback_7_bits_debug_isPerfCnt,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_6_valid,io_exuWriteback_6_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_6_bits_data_0,io_exuWriteback_6_bits_data_0,64);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_6_bits_robIdx_value,io_exuWriteback_6_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_5_valid,io_exuWriteback_5_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_5_bits_data_0,io_exuWriteback_5_bits_data_0,128);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_5_bits_robIdx_value,io_exuWriteback_5_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_5_bits_redirect_valid,io_exuWriteback_5_bits_redirect_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken,io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_5_bits_fflags,io_exuWriteback_5_bits_fflags,5);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_5_bits_wflags,io_exuWriteback_5_bits_wflags,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_4_valid,io_exuWriteback_4_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_4_bits_data_0,io_exuWriteback_4_bits_data_0,64);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_4_bits_robIdx_value,io_exuWriteback_4_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_3_valid,io_exuWriteback_3_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_3_bits_data_0,io_exuWriteback_3_bits_data_0,64);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_3_bits_robIdx_value,io_exuWriteback_3_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_3_bits_redirect_valid,io_exuWriteback_3_bits_redirect_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken,io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_2_valid,io_exuWriteback_2_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_2_bits_data_0,io_exuWriteback_2_bits_data_0,64);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_2_bits_robIdx_value,io_exuWriteback_2_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_1_valid,io_exuWriteback_1_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_1_bits_data_0,io_exuWriteback_1_bits_data_0,64);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_1_bits_robIdx_value,io_exuWriteback_1_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_1_bits_redirect_valid,io_exuWriteback_1_bits_redirect_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken,io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_0_valid,io_exuWriteback_0_valid,1);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_0_bits_data_0,io_exuWriteback_0_bits_data_0,64);
            `TCNT_CHECK_SIG_XZ(io_exuWriteback_0_bits_robIdx_value,io_exuWriteback_0_bits_robIdx_value,8);
            `TCNT_CHECK_SIG_XZ(io_writebackNums_0_bits,io_writebackNums_0_bits,5);
            `TCNT_CHECK_SIG_XZ(io_writebackNums_1_bits,io_writebackNums_1_bits,5);
            `TCNT_CHECK_SIG_XZ(io_writebackNums_2_bits,io_writebackNums_2_bits,5);
            `TCNT_CHECK_SIG_XZ(io_writebackNums_3_bits,io_writebackNums_3_bits,5);
            `TCNT_CHECK_SIG_XZ(io_writebackNums_4_bits,io_writebackNums_4_bits,5);
            `TCNT_CHECK_SIG_XZ(io_writebackNums_5_bits,io_writebackNums_5_bits,5);
            `TCNT_CHECK_SIG_XZ(io_writebackNums_6_bits,io_writebackNums_6_bits,5);
            `TCNT_CHECK_SIG_XZ(io_writebackNums_7_bits,io_writebackNums_7_bits,5);
            `TCNT_CHECK_SIG_XZ(io_writebackNums_8_bits,io_writebackNums_8_bits,5);
            `TCNT_CHECK_SIG_XZ(io_writebackNums_9_bits,io_writebackNums_9_bits,5);
            `TCNT_CHECK_SIG_XZ(io_writebackNums_10_bits,io_writebackNums_10_bits,5);
            `TCNT_CHECK_SIG_XZ(io_writebackNums_11_bits,io_writebackNums_11_bits,5);
            `TCNT_CHECK_SIG_XZ(io_writebackNums_12_bits,io_writebackNums_12_bits,5);
            `TCNT_CHECK_SIG_XZ(io_writebackNums_13_bits,io_writebackNums_13_bits,5);
            `TCNT_CHECK_SIG_XZ(io_writebackNums_14_bits,io_writebackNums_14_bits,5);
            `TCNT_CHECK_SIG_XZ(io_writebackNums_15_bits,io_writebackNums_15_bits,5);
            `TCNT_CHECK_SIG_XZ(io_writebackNums_16_bits,io_writebackNums_16_bits,5);
            `TCNT_CHECK_SIG_XZ(io_writebackNums_17_bits,io_writebackNums_17_bits,5);
            `TCNT_CHECK_SIG_XZ(io_writebackNums_18_bits,io_writebackNums_18_bits,5);
            `TCNT_CHECK_SIG_XZ(io_writebackNums_19_bits,io_writebackNums_19_bits,5);
            `TCNT_CHECK_SIG_XZ(io_writebackNums_20_bits,io_writebackNums_20_bits,5);
            `TCNT_CHECK_SIG_XZ(io_writebackNums_21_bits,io_writebackNums_21_bits,5);
            `TCNT_CHECK_SIG_XZ(io_writebackNums_22_bits,io_writebackNums_22_bits,5);
            `TCNT_CHECK_SIG_XZ(io_writebackNums_23_bits,io_writebackNums_23_bits,5);
            `TCNT_CHECK_SIG_XZ(io_writebackNums_24_bits,io_writebackNums_24_bits,5);
            `TCNT_CHECK_SIG_XZ(io_writebackNeedFlush_0,io_writebackNeedFlush_0,1);
            `TCNT_CHECK_SIG_XZ(io_writebackNeedFlush_1,io_writebackNeedFlush_1,1);
            `TCNT_CHECK_SIG_XZ(io_writebackNeedFlush_2,io_writebackNeedFlush_2,1);
            `TCNT_CHECK_SIG_XZ(io_writebackNeedFlush_6,io_writebackNeedFlush_6,1);
            `TCNT_CHECK_SIG_XZ(io_writebackNeedFlush_7,io_writebackNeedFlush_7,1);
            `TCNT_CHECK_SIG_XZ(io_writebackNeedFlush_8,io_writebackNeedFlush_8,1);
            `TCNT_CHECK_SIG_XZ(io_writebackNeedFlush_9,io_writebackNeedFlush_9,1);
            `TCNT_CHECK_SIG_XZ(io_writebackNeedFlush_10,io_writebackNeedFlush_10,1);
            `TCNT_CHECK_SIG_XZ(io_writebackNeedFlush_11,io_writebackNeedFlush_11,1);
            `TCNT_CHECK_SIG_XZ(io_writebackNeedFlush_12,io_writebackNeedFlush_12,1);

        end
        //if(xxxTODOxxx==1'b1) begin
        //    mon_tr = WriteBack_in_agent_xaction::type_id::create("mon_tr");
        //    mon_tr.io_writeback_24_valid = io_writeback_24_valid;
        //    mon_tr.io_writeback_24_bits_data_0 = io_writeback_24_bits_data_0;
        //    mon_tr.io_writeback_24_bits_pdest = io_writeback_24_bits_pdest;
        //    mon_tr.io_writeback_24_bits_robIdx_flag = io_writeback_24_bits_robIdx_flag;
        //    mon_tr.io_writeback_24_bits_robIdx_value = io_writeback_24_bits_robIdx_value;
        //    mon_tr.io_writeback_24_bits_vecWen = io_writeback_24_bits_vecWen;
        //    mon_tr.io_writeback_24_bits_v0Wen = io_writeback_24_bits_v0Wen;
        //    mon_tr.io_writeback_24_bits_vlWen = io_writeback_24_bits_vlWen;
        //    mon_tr.io_writeback_24_bits_exceptionVec_0 = io_writeback_24_bits_exceptionVec_0;
        //    mon_tr.io_writeback_24_bits_exceptionVec_1 = io_writeback_24_bits_exceptionVec_1;
        //    mon_tr.io_writeback_24_bits_exceptionVec_2 = io_writeback_24_bits_exceptionVec_2;
        //    mon_tr.io_writeback_24_bits_exceptionVec_3 = io_writeback_24_bits_exceptionVec_3;
        //    mon_tr.io_writeback_24_bits_exceptionVec_4 = io_writeback_24_bits_exceptionVec_4;
        //    mon_tr.io_writeback_24_bits_exceptionVec_5 = io_writeback_24_bits_exceptionVec_5;
        //    mon_tr.io_writeback_24_bits_exceptionVec_6 = io_writeback_24_bits_exceptionVec_6;
        //    mon_tr.io_writeback_24_bits_exceptionVec_7 = io_writeback_24_bits_exceptionVec_7;
        //    mon_tr.io_writeback_24_bits_exceptionVec_8 = io_writeback_24_bits_exceptionVec_8;
        //    mon_tr.io_writeback_24_bits_exceptionVec_9 = io_writeback_24_bits_exceptionVec_9;
        //    mon_tr.io_writeback_24_bits_exceptionVec_10 = io_writeback_24_bits_exceptionVec_10;
        //    mon_tr.io_writeback_24_bits_exceptionVec_11 = io_writeback_24_bits_exceptionVec_11;
        //    mon_tr.io_writeback_24_bits_exceptionVec_12 = io_writeback_24_bits_exceptionVec_12;
        //    mon_tr.io_writeback_24_bits_exceptionVec_13 = io_writeback_24_bits_exceptionVec_13;
        //    mon_tr.io_writeback_24_bits_exceptionVec_14 = io_writeback_24_bits_exceptionVec_14;
        //    mon_tr.io_writeback_24_bits_exceptionVec_15 = io_writeback_24_bits_exceptionVec_15;
        //    mon_tr.io_writeback_24_bits_exceptionVec_16 = io_writeback_24_bits_exceptionVec_16;
        //    mon_tr.io_writeback_24_bits_exceptionVec_17 = io_writeback_24_bits_exceptionVec_17;
        //    mon_tr.io_writeback_24_bits_exceptionVec_18 = io_writeback_24_bits_exceptionVec_18;
        //    mon_tr.io_writeback_24_bits_exceptionVec_19 = io_writeback_24_bits_exceptionVec_19;
        //    mon_tr.io_writeback_24_bits_exceptionVec_20 = io_writeback_24_bits_exceptionVec_20;
        //    mon_tr.io_writeback_24_bits_exceptionVec_21 = io_writeback_24_bits_exceptionVec_21;
        //    mon_tr.io_writeback_24_bits_exceptionVec_22 = io_writeback_24_bits_exceptionVec_22;
        //    mon_tr.io_writeback_24_bits_exceptionVec_23 = io_writeback_24_bits_exceptionVec_23;
        //    mon_tr.io_writeback_24_bits_flushPipe = io_writeback_24_bits_flushPipe;
        //    mon_tr.io_writeback_24_bits_replay = io_writeback_24_bits_replay;
        //    mon_tr.io_writeback_24_bits_trigger = io_writeback_24_bits_trigger;
        //    mon_tr.io_writeback_24_bits_vls_vpu_vill = io_writeback_24_bits_vls_vpu_vill;
        //    mon_tr.io_writeback_24_bits_vls_vpu_vma = io_writeback_24_bits_vls_vpu_vma;
        //    mon_tr.io_writeback_24_bits_vls_vpu_vta = io_writeback_24_bits_vls_vpu_vta;
        //    mon_tr.io_writeback_24_bits_vls_vpu_vsew = io_writeback_24_bits_vls_vpu_vsew;
        //    mon_tr.io_writeback_24_bits_vls_vpu_vlmul = io_writeback_24_bits_vls_vpu_vlmul;
        //    mon_tr.io_writeback_24_bits_vls_vpu_specVill = io_writeback_24_bits_vls_vpu_specVill;
        //    mon_tr.io_writeback_24_bits_vls_vpu_specVma = io_writeback_24_bits_vls_vpu_specVma;
        //    mon_tr.io_writeback_24_bits_vls_vpu_specVta = io_writeback_24_bits_vls_vpu_specVta;
        //    mon_tr.io_writeback_24_bits_vls_vpu_specVsew = io_writeback_24_bits_vls_vpu_specVsew;
        //    mon_tr.io_writeback_24_bits_vls_vpu_specVlmul = io_writeback_24_bits_vls_vpu_specVlmul;
        //    mon_tr.io_writeback_24_bits_vls_vpu_vm = io_writeback_24_bits_vls_vpu_vm;
        //    mon_tr.io_writeback_24_bits_vls_vpu_vstart = io_writeback_24_bits_vls_vpu_vstart;
        //    mon_tr.io_writeback_24_bits_vls_vpu_frm = io_writeback_24_bits_vls_vpu_frm;
        //    mon_tr.io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst = io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst;
        //    mon_tr.io_writeback_24_bits_vls_vpu_fpu_isFP32Instr = io_writeback_24_bits_vls_vpu_fpu_isFP32Instr;
        //    mon_tr.io_writeback_24_bits_vls_vpu_fpu_isFP64Instr = io_writeback_24_bits_vls_vpu_fpu_isFP64Instr;
        //    mon_tr.io_writeback_24_bits_vls_vpu_fpu_isReduction = io_writeback_24_bits_vls_vpu_fpu_isReduction;
        //    mon_tr.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2 = io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2;
        //    mon_tr.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4 = io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4;
        //    mon_tr.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8 = io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8;
        //    mon_tr.io_writeback_24_bits_vls_vpu_vxrm = io_writeback_24_bits_vls_vpu_vxrm;
        //    mon_tr.io_writeback_24_bits_vls_vpu_vuopIdx = io_writeback_24_bits_vls_vpu_vuopIdx;
        //    mon_tr.io_writeback_24_bits_vls_vpu_lastUop = io_writeback_24_bits_vls_vpu_lastUop;
        //    mon_tr.io_writeback_24_bits_vls_vpu_vmask = io_writeback_24_bits_vls_vpu_vmask;
        //    mon_tr.io_writeback_24_bits_vls_vpu_vl = io_writeback_24_bits_vls_vpu_vl;
        //    mon_tr.io_writeback_24_bits_vls_vpu_nf = io_writeback_24_bits_vls_vpu_nf;
        //    mon_tr.io_writeback_24_bits_vls_vpu_veew = io_writeback_24_bits_vls_vpu_veew;
        //    mon_tr.io_writeback_24_bits_vls_vpu_isReverse = io_writeback_24_bits_vls_vpu_isReverse;
        //    mon_tr.io_writeback_24_bits_vls_vpu_isExt = io_writeback_24_bits_vls_vpu_isExt;
        //    mon_tr.io_writeback_24_bits_vls_vpu_isNarrow = io_writeback_24_bits_vls_vpu_isNarrow;
        //    mon_tr.io_writeback_24_bits_vls_vpu_isDstMask = io_writeback_24_bits_vls_vpu_isDstMask;
        //    mon_tr.io_writeback_24_bits_vls_vpu_isOpMask = io_writeback_24_bits_vls_vpu_isOpMask;
        //    mon_tr.io_writeback_24_bits_vls_vpu_isMove = io_writeback_24_bits_vls_vpu_isMove;
        //    mon_tr.io_writeback_24_bits_vls_vpu_isDependOldVd = io_writeback_24_bits_vls_vpu_isDependOldVd;
        //    mon_tr.io_writeback_24_bits_vls_vpu_isWritePartVd = io_writeback_24_bits_vls_vpu_isWritePartVd;
        //    mon_tr.io_writeback_24_bits_vls_vpu_isVleff = io_writeback_24_bits_vls_vpu_isVleff;
        //    mon_tr.io_writeback_24_bits_vls_oldVdPsrc = io_writeback_24_bits_vls_oldVdPsrc;
        //    mon_tr.io_writeback_24_bits_vls_vdIdx = io_writeback_24_bits_vls_vdIdx;
        //    mon_tr.io_writeback_24_bits_vls_vdIdxInField = io_writeback_24_bits_vls_vdIdxInField;
        //    mon_tr.io_writeback_24_bits_vls_isIndexed = io_writeback_24_bits_vls_isIndexed;
        //    mon_tr.io_writeback_24_bits_vls_isMasked = io_writeback_24_bits_vls_isMasked;
        //    mon_tr.io_writeback_24_bits_vls_isStrided = io_writeback_24_bits_vls_isStrided;
        //    mon_tr.io_writeback_24_bits_vls_isWhole = io_writeback_24_bits_vls_isWhole;
        //    mon_tr.io_writeback_24_bits_vls_isVecLoad = io_writeback_24_bits_vls_isVecLoad;
        //    mon_tr.io_writeback_24_bits_vls_isVlm = io_writeback_24_bits_vls_isVlm;
        //    mon_tr.io_writeback_24_bits_debug_isMMIO = io_writeback_24_bits_debug_isMMIO;
        //    mon_tr.io_writeback_24_bits_debug_isNCIO = io_writeback_24_bits_debug_isNCIO;
        //    mon_tr.io_writeback_24_bits_debug_isPerfCnt = io_writeback_24_bits_debug_isPerfCnt;
        //    mon_tr.io_writeback_24_bits_debug_paddr = io_writeback_24_bits_debug_paddr;
        //    mon_tr.io_writeback_24_bits_debug_vaddr = io_writeback_24_bits_debug_vaddr;
        //    mon_tr.io_writeback_24_bits_debugInfo_eliminatedMove = io_writeback_24_bits_debugInfo_eliminatedMove;
        //    mon_tr.io_writeback_24_bits_debugInfo_renameTime = io_writeback_24_bits_debugInfo_renameTime;
        //    mon_tr.io_writeback_24_bits_debugInfo_dispatchTime = io_writeback_24_bits_debugInfo_dispatchTime;
        //    mon_tr.io_writeback_24_bits_debugInfo_enqRsTime = io_writeback_24_bits_debugInfo_enqRsTime;
        //    mon_tr.io_writeback_24_bits_debugInfo_selectTime = io_writeback_24_bits_debugInfo_selectTime;
        //    mon_tr.io_writeback_24_bits_debugInfo_issueTime = io_writeback_24_bits_debugInfo_issueTime;
        //    mon_tr.io_writeback_24_bits_debugInfo_writebackTime = io_writeback_24_bits_debugInfo_writebackTime;
        //    mon_tr.io_writeback_24_bits_debugInfo_runahead_checkpoint_id = io_writeback_24_bits_debugInfo_runahead_checkpoint_id;
        //    mon_tr.io_writeback_24_bits_debugInfo_tlbFirstReqTime = io_writeback_24_bits_debugInfo_tlbFirstReqTime;
        //    mon_tr.io_writeback_24_bits_debugInfo_tlbRespTime = io_writeback_24_bits_debugInfo_tlbRespTime;
        //    mon_tr.io_writeback_24_bits_debug_seqNum = io_writeback_24_bits_debug_seqNum;
        //    mon_tr.io_writeback_23_valid = io_writeback_23_valid;
        //    mon_tr.io_writeback_23_bits_data_0 = io_writeback_23_bits_data_0;
        //    mon_tr.io_writeback_23_bits_pdest = io_writeback_23_bits_pdest;
        //    mon_tr.io_writeback_23_bits_robIdx_flag = io_writeback_23_bits_robIdx_flag;
        //    mon_tr.io_writeback_23_bits_robIdx_value = io_writeback_23_bits_robIdx_value;
        //    mon_tr.io_writeback_23_bits_vecWen = io_writeback_23_bits_vecWen;
        //    mon_tr.io_writeback_23_bits_v0Wen = io_writeback_23_bits_v0Wen;
        //    mon_tr.io_writeback_23_bits_vlWen = io_writeback_23_bits_vlWen;
        //    mon_tr.io_writeback_23_bits_exceptionVec_0 = io_writeback_23_bits_exceptionVec_0;
        //    mon_tr.io_writeback_23_bits_exceptionVec_1 = io_writeback_23_bits_exceptionVec_1;
        //    mon_tr.io_writeback_23_bits_exceptionVec_2 = io_writeback_23_bits_exceptionVec_2;
        //    mon_tr.io_writeback_23_bits_exceptionVec_3 = io_writeback_23_bits_exceptionVec_3;
        //    mon_tr.io_writeback_23_bits_exceptionVec_4 = io_writeback_23_bits_exceptionVec_4;
        //    mon_tr.io_writeback_23_bits_exceptionVec_5 = io_writeback_23_bits_exceptionVec_5;
        //    mon_tr.io_writeback_23_bits_exceptionVec_6 = io_writeback_23_bits_exceptionVec_6;
        //    mon_tr.io_writeback_23_bits_exceptionVec_7 = io_writeback_23_bits_exceptionVec_7;
        //    mon_tr.io_writeback_23_bits_exceptionVec_8 = io_writeback_23_bits_exceptionVec_8;
        //    mon_tr.io_writeback_23_bits_exceptionVec_9 = io_writeback_23_bits_exceptionVec_9;
        //    mon_tr.io_writeback_23_bits_exceptionVec_10 = io_writeback_23_bits_exceptionVec_10;
        //    mon_tr.io_writeback_23_bits_exceptionVec_11 = io_writeback_23_bits_exceptionVec_11;
        //    mon_tr.io_writeback_23_bits_exceptionVec_12 = io_writeback_23_bits_exceptionVec_12;
        //    mon_tr.io_writeback_23_bits_exceptionVec_13 = io_writeback_23_bits_exceptionVec_13;
        //    mon_tr.io_writeback_23_bits_exceptionVec_14 = io_writeback_23_bits_exceptionVec_14;
        //    mon_tr.io_writeback_23_bits_exceptionVec_15 = io_writeback_23_bits_exceptionVec_15;
        //    mon_tr.io_writeback_23_bits_exceptionVec_16 = io_writeback_23_bits_exceptionVec_16;
        //    mon_tr.io_writeback_23_bits_exceptionVec_17 = io_writeback_23_bits_exceptionVec_17;
        //    mon_tr.io_writeback_23_bits_exceptionVec_18 = io_writeback_23_bits_exceptionVec_18;
        //    mon_tr.io_writeback_23_bits_exceptionVec_19 = io_writeback_23_bits_exceptionVec_19;
        //    mon_tr.io_writeback_23_bits_exceptionVec_20 = io_writeback_23_bits_exceptionVec_20;
        //    mon_tr.io_writeback_23_bits_exceptionVec_21 = io_writeback_23_bits_exceptionVec_21;
        //    mon_tr.io_writeback_23_bits_exceptionVec_22 = io_writeback_23_bits_exceptionVec_22;
        //    mon_tr.io_writeback_23_bits_exceptionVec_23 = io_writeback_23_bits_exceptionVec_23;
        //    mon_tr.io_writeback_23_bits_flushPipe = io_writeback_23_bits_flushPipe;
        //    mon_tr.io_writeback_23_bits_replay = io_writeback_23_bits_replay;
        //    mon_tr.io_writeback_23_bits_trigger = io_writeback_23_bits_trigger;
        //    mon_tr.io_writeback_23_bits_vls_vpu_vill = io_writeback_23_bits_vls_vpu_vill;
        //    mon_tr.io_writeback_23_bits_vls_vpu_vma = io_writeback_23_bits_vls_vpu_vma;
        //    mon_tr.io_writeback_23_bits_vls_vpu_vta = io_writeback_23_bits_vls_vpu_vta;
        //    mon_tr.io_writeback_23_bits_vls_vpu_vsew = io_writeback_23_bits_vls_vpu_vsew;
        //    mon_tr.io_writeback_23_bits_vls_vpu_vlmul = io_writeback_23_bits_vls_vpu_vlmul;
        //    mon_tr.io_writeback_23_bits_vls_vpu_specVill = io_writeback_23_bits_vls_vpu_specVill;
        //    mon_tr.io_writeback_23_bits_vls_vpu_specVma = io_writeback_23_bits_vls_vpu_specVma;
        //    mon_tr.io_writeback_23_bits_vls_vpu_specVta = io_writeback_23_bits_vls_vpu_specVta;
        //    mon_tr.io_writeback_23_bits_vls_vpu_specVsew = io_writeback_23_bits_vls_vpu_specVsew;
        //    mon_tr.io_writeback_23_bits_vls_vpu_specVlmul = io_writeback_23_bits_vls_vpu_specVlmul;
        //    mon_tr.io_writeback_23_bits_vls_vpu_vm = io_writeback_23_bits_vls_vpu_vm;
        //    mon_tr.io_writeback_23_bits_vls_vpu_vstart = io_writeback_23_bits_vls_vpu_vstart;
        //    mon_tr.io_writeback_23_bits_vls_vpu_frm = io_writeback_23_bits_vls_vpu_frm;
        //    mon_tr.io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst = io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst;
        //    mon_tr.io_writeback_23_bits_vls_vpu_fpu_isFP32Instr = io_writeback_23_bits_vls_vpu_fpu_isFP32Instr;
        //    mon_tr.io_writeback_23_bits_vls_vpu_fpu_isFP64Instr = io_writeback_23_bits_vls_vpu_fpu_isFP64Instr;
        //    mon_tr.io_writeback_23_bits_vls_vpu_fpu_isReduction = io_writeback_23_bits_vls_vpu_fpu_isReduction;
        //    mon_tr.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2 = io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2;
        //    mon_tr.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4 = io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4;
        //    mon_tr.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8 = io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8;
        //    mon_tr.io_writeback_23_bits_vls_vpu_vxrm = io_writeback_23_bits_vls_vpu_vxrm;
        //    mon_tr.io_writeback_23_bits_vls_vpu_vuopIdx = io_writeback_23_bits_vls_vpu_vuopIdx;
        //    mon_tr.io_writeback_23_bits_vls_vpu_lastUop = io_writeback_23_bits_vls_vpu_lastUop;
        //    mon_tr.io_writeback_23_bits_vls_vpu_vmask = io_writeback_23_bits_vls_vpu_vmask;
        //    mon_tr.io_writeback_23_bits_vls_vpu_vl = io_writeback_23_bits_vls_vpu_vl;
        //    mon_tr.io_writeback_23_bits_vls_vpu_nf = io_writeback_23_bits_vls_vpu_nf;
        //    mon_tr.io_writeback_23_bits_vls_vpu_veew = io_writeback_23_bits_vls_vpu_veew;
        //    mon_tr.io_writeback_23_bits_vls_vpu_isReverse = io_writeback_23_bits_vls_vpu_isReverse;
        //    mon_tr.io_writeback_23_bits_vls_vpu_isExt = io_writeback_23_bits_vls_vpu_isExt;
        //    mon_tr.io_writeback_23_bits_vls_vpu_isNarrow = io_writeback_23_bits_vls_vpu_isNarrow;
        //    mon_tr.io_writeback_23_bits_vls_vpu_isDstMask = io_writeback_23_bits_vls_vpu_isDstMask;
        //    mon_tr.io_writeback_23_bits_vls_vpu_isOpMask = io_writeback_23_bits_vls_vpu_isOpMask;
        //    mon_tr.io_writeback_23_bits_vls_vpu_isMove = io_writeback_23_bits_vls_vpu_isMove;
        //    mon_tr.io_writeback_23_bits_vls_vpu_isDependOldVd = io_writeback_23_bits_vls_vpu_isDependOldVd;
        //    mon_tr.io_writeback_23_bits_vls_vpu_isWritePartVd = io_writeback_23_bits_vls_vpu_isWritePartVd;
        //    mon_tr.io_writeback_23_bits_vls_vpu_isVleff = io_writeback_23_bits_vls_vpu_isVleff;
        //    mon_tr.io_writeback_23_bits_vls_oldVdPsrc = io_writeback_23_bits_vls_oldVdPsrc;
        //    mon_tr.io_writeback_23_bits_vls_vdIdx = io_writeback_23_bits_vls_vdIdx;
        //    mon_tr.io_writeback_23_bits_vls_vdIdxInField = io_writeback_23_bits_vls_vdIdxInField;
        //    mon_tr.io_writeback_23_bits_vls_isIndexed = io_writeback_23_bits_vls_isIndexed;
        //    mon_tr.io_writeback_23_bits_vls_isMasked = io_writeback_23_bits_vls_isMasked;
        //    mon_tr.io_writeback_23_bits_vls_isStrided = io_writeback_23_bits_vls_isStrided;
        //    mon_tr.io_writeback_23_bits_vls_isWhole = io_writeback_23_bits_vls_isWhole;
        //    mon_tr.io_writeback_23_bits_vls_isVecLoad = io_writeback_23_bits_vls_isVecLoad;
        //    mon_tr.io_writeback_23_bits_vls_isVlm = io_writeback_23_bits_vls_isVlm;
        //    mon_tr.io_writeback_23_bits_debug_isMMIO = io_writeback_23_bits_debug_isMMIO;
        //    mon_tr.io_writeback_23_bits_debug_isNCIO = io_writeback_23_bits_debug_isNCIO;
        //    mon_tr.io_writeback_23_bits_debug_isPerfCnt = io_writeback_23_bits_debug_isPerfCnt;
        //    mon_tr.io_writeback_23_bits_debug_paddr = io_writeback_23_bits_debug_paddr;
        //    mon_tr.io_writeback_23_bits_debug_vaddr = io_writeback_23_bits_debug_vaddr;
        //    mon_tr.io_writeback_23_bits_debugInfo_eliminatedMove = io_writeback_23_bits_debugInfo_eliminatedMove;
        //    mon_tr.io_writeback_23_bits_debugInfo_renameTime = io_writeback_23_bits_debugInfo_renameTime;
        //    mon_tr.io_writeback_23_bits_debugInfo_dispatchTime = io_writeback_23_bits_debugInfo_dispatchTime;
        //    mon_tr.io_writeback_23_bits_debugInfo_enqRsTime = io_writeback_23_bits_debugInfo_enqRsTime;
        //    mon_tr.io_writeback_23_bits_debugInfo_selectTime = io_writeback_23_bits_debugInfo_selectTime;
        //    mon_tr.io_writeback_23_bits_debugInfo_issueTime = io_writeback_23_bits_debugInfo_issueTime;
        //    mon_tr.io_writeback_23_bits_debugInfo_writebackTime = io_writeback_23_bits_debugInfo_writebackTime;
        //    mon_tr.io_writeback_23_bits_debugInfo_runahead_checkpoint_id = io_writeback_23_bits_debugInfo_runahead_checkpoint_id;
        //    mon_tr.io_writeback_23_bits_debugInfo_tlbFirstReqTime = io_writeback_23_bits_debugInfo_tlbFirstReqTime;
        //    mon_tr.io_writeback_23_bits_debugInfo_tlbRespTime = io_writeback_23_bits_debugInfo_tlbRespTime;
        //    mon_tr.io_writeback_23_bits_debug_seqNum = io_writeback_23_bits_debug_seqNum;
        //    mon_tr.io_writeback_22_valid = io_writeback_22_valid;
        //    mon_tr.io_writeback_22_bits_data_0 = io_writeback_22_bits_data_0;
        //    mon_tr.io_writeback_22_bits_pdest = io_writeback_22_bits_pdest;
        //    mon_tr.io_writeback_22_bits_robIdx_flag = io_writeback_22_bits_robIdx_flag;
        //    mon_tr.io_writeback_22_bits_robIdx_value = io_writeback_22_bits_robIdx_value;
        //    mon_tr.io_writeback_22_bits_intWen = io_writeback_22_bits_intWen;
        //    mon_tr.io_writeback_22_bits_fpWen = io_writeback_22_bits_fpWen;
        //    mon_tr.io_writeback_22_bits_exceptionVec_0 = io_writeback_22_bits_exceptionVec_0;
        //    mon_tr.io_writeback_22_bits_exceptionVec_1 = io_writeback_22_bits_exceptionVec_1;
        //    mon_tr.io_writeback_22_bits_exceptionVec_2 = io_writeback_22_bits_exceptionVec_2;
        //    mon_tr.io_writeback_22_bits_exceptionVec_3 = io_writeback_22_bits_exceptionVec_3;
        //    mon_tr.io_writeback_22_bits_exceptionVec_4 = io_writeback_22_bits_exceptionVec_4;
        //    mon_tr.io_writeback_22_bits_exceptionVec_5 = io_writeback_22_bits_exceptionVec_5;
        //    mon_tr.io_writeback_22_bits_exceptionVec_6 = io_writeback_22_bits_exceptionVec_6;
        //    mon_tr.io_writeback_22_bits_exceptionVec_7 = io_writeback_22_bits_exceptionVec_7;
        //    mon_tr.io_writeback_22_bits_exceptionVec_8 = io_writeback_22_bits_exceptionVec_8;
        //    mon_tr.io_writeback_22_bits_exceptionVec_9 = io_writeback_22_bits_exceptionVec_9;
        //    mon_tr.io_writeback_22_bits_exceptionVec_10 = io_writeback_22_bits_exceptionVec_10;
        //    mon_tr.io_writeback_22_bits_exceptionVec_11 = io_writeback_22_bits_exceptionVec_11;
        //    mon_tr.io_writeback_22_bits_exceptionVec_12 = io_writeback_22_bits_exceptionVec_12;
        //    mon_tr.io_writeback_22_bits_exceptionVec_13 = io_writeback_22_bits_exceptionVec_13;
        //    mon_tr.io_writeback_22_bits_exceptionVec_14 = io_writeback_22_bits_exceptionVec_14;
        //    mon_tr.io_writeback_22_bits_exceptionVec_15 = io_writeback_22_bits_exceptionVec_15;
        //    mon_tr.io_writeback_22_bits_exceptionVec_16 = io_writeback_22_bits_exceptionVec_16;
        //    mon_tr.io_writeback_22_bits_exceptionVec_17 = io_writeback_22_bits_exceptionVec_17;
        //    mon_tr.io_writeback_22_bits_exceptionVec_18 = io_writeback_22_bits_exceptionVec_18;
        //    mon_tr.io_writeback_22_bits_exceptionVec_19 = io_writeback_22_bits_exceptionVec_19;
        //    mon_tr.io_writeback_22_bits_exceptionVec_20 = io_writeback_22_bits_exceptionVec_20;
        //    mon_tr.io_writeback_22_bits_exceptionVec_21 = io_writeback_22_bits_exceptionVec_21;
        //    mon_tr.io_writeback_22_bits_exceptionVec_22 = io_writeback_22_bits_exceptionVec_22;
        //    mon_tr.io_writeback_22_bits_exceptionVec_23 = io_writeback_22_bits_exceptionVec_23;
        //    mon_tr.io_writeback_22_bits_flushPipe = io_writeback_22_bits_flushPipe;
        //    mon_tr.io_writeback_22_bits_replay = io_writeback_22_bits_replay;
        //    mon_tr.io_writeback_22_bits_lqIdx_flag = io_writeback_22_bits_lqIdx_flag;
        //    mon_tr.io_writeback_22_bits_lqIdx_value = io_writeback_22_bits_lqIdx_value;
        //    mon_tr.io_writeback_22_bits_trigger = io_writeback_22_bits_trigger;
        //    mon_tr.io_writeback_22_bits_predecodeInfo_valid = io_writeback_22_bits_predecodeInfo_valid;
        //    mon_tr.io_writeback_22_bits_predecodeInfo_isRVC = io_writeback_22_bits_predecodeInfo_isRVC;
        //    mon_tr.io_writeback_22_bits_predecodeInfo_brType = io_writeback_22_bits_predecodeInfo_brType;
        //    mon_tr.io_writeback_22_bits_predecodeInfo_isCall = io_writeback_22_bits_predecodeInfo_isCall;
        //    mon_tr.io_writeback_22_bits_predecodeInfo_isRet = io_writeback_22_bits_predecodeInfo_isRet;
        //    mon_tr.io_writeback_22_bits_debug_isMMIO = io_writeback_22_bits_debug_isMMIO;
        //    mon_tr.io_writeback_22_bits_debug_isNCIO = io_writeback_22_bits_debug_isNCIO;
        //    mon_tr.io_writeback_22_bits_debug_isPerfCnt = io_writeback_22_bits_debug_isPerfCnt;
        //    mon_tr.io_writeback_22_bits_debug_paddr = io_writeback_22_bits_debug_paddr;
        //    mon_tr.io_writeback_22_bits_debug_vaddr = io_writeback_22_bits_debug_vaddr;
        //    mon_tr.io_writeback_22_bits_debugInfo_eliminatedMove = io_writeback_22_bits_debugInfo_eliminatedMove;
        //    mon_tr.io_writeback_22_bits_debugInfo_renameTime = io_writeback_22_bits_debugInfo_renameTime;
        //    mon_tr.io_writeback_22_bits_debugInfo_dispatchTime = io_writeback_22_bits_debugInfo_dispatchTime;
        //    mon_tr.io_writeback_22_bits_debugInfo_enqRsTime = io_writeback_22_bits_debugInfo_enqRsTime;
        //    mon_tr.io_writeback_22_bits_debugInfo_selectTime = io_writeback_22_bits_debugInfo_selectTime;
        //    mon_tr.io_writeback_22_bits_debugInfo_issueTime = io_writeback_22_bits_debugInfo_issueTime;
        //    mon_tr.io_writeback_22_bits_debugInfo_writebackTime = io_writeback_22_bits_debugInfo_writebackTime;
        //    mon_tr.io_writeback_22_bits_debugInfo_runahead_checkpoint_id = io_writeback_22_bits_debugInfo_runahead_checkpoint_id;
        //    mon_tr.io_writeback_22_bits_debugInfo_tlbFirstReqTime = io_writeback_22_bits_debugInfo_tlbFirstReqTime;
        //    mon_tr.io_writeback_22_bits_debugInfo_tlbRespTime = io_writeback_22_bits_debugInfo_tlbRespTime;
        //    mon_tr.io_writeback_22_bits_debug_seqNum = io_writeback_22_bits_debug_seqNum;
        //    mon_tr.io_writeback_21_valid = io_writeback_21_valid;
        //    mon_tr.io_writeback_21_bits_data_0 = io_writeback_21_bits_data_0;
        //    mon_tr.io_writeback_21_bits_pdest = io_writeback_21_bits_pdest;
        //    mon_tr.io_writeback_21_bits_robIdx_flag = io_writeback_21_bits_robIdx_flag;
        //    mon_tr.io_writeback_21_bits_robIdx_value = io_writeback_21_bits_robIdx_value;
        //    mon_tr.io_writeback_21_bits_intWen = io_writeback_21_bits_intWen;
        //    mon_tr.io_writeback_21_bits_fpWen = io_writeback_21_bits_fpWen;
        //    mon_tr.io_writeback_21_bits_exceptionVec_0 = io_writeback_21_bits_exceptionVec_0;
        //    mon_tr.io_writeback_21_bits_exceptionVec_1 = io_writeback_21_bits_exceptionVec_1;
        //    mon_tr.io_writeback_21_bits_exceptionVec_2 = io_writeback_21_bits_exceptionVec_2;
        //    mon_tr.io_writeback_21_bits_exceptionVec_3 = io_writeback_21_bits_exceptionVec_3;
        //    mon_tr.io_writeback_21_bits_exceptionVec_4 = io_writeback_21_bits_exceptionVec_4;
        //    mon_tr.io_writeback_21_bits_exceptionVec_5 = io_writeback_21_bits_exceptionVec_5;
        //    mon_tr.io_writeback_21_bits_exceptionVec_6 = io_writeback_21_bits_exceptionVec_6;
        //    mon_tr.io_writeback_21_bits_exceptionVec_7 = io_writeback_21_bits_exceptionVec_7;
        //    mon_tr.io_writeback_21_bits_exceptionVec_8 = io_writeback_21_bits_exceptionVec_8;
        //    mon_tr.io_writeback_21_bits_exceptionVec_9 = io_writeback_21_bits_exceptionVec_9;
        //    mon_tr.io_writeback_21_bits_exceptionVec_10 = io_writeback_21_bits_exceptionVec_10;
        //    mon_tr.io_writeback_21_bits_exceptionVec_11 = io_writeback_21_bits_exceptionVec_11;
        //    mon_tr.io_writeback_21_bits_exceptionVec_12 = io_writeback_21_bits_exceptionVec_12;
        //    mon_tr.io_writeback_21_bits_exceptionVec_13 = io_writeback_21_bits_exceptionVec_13;
        //    mon_tr.io_writeback_21_bits_exceptionVec_14 = io_writeback_21_bits_exceptionVec_14;
        //    mon_tr.io_writeback_21_bits_exceptionVec_15 = io_writeback_21_bits_exceptionVec_15;
        //    mon_tr.io_writeback_21_bits_exceptionVec_16 = io_writeback_21_bits_exceptionVec_16;
        //    mon_tr.io_writeback_21_bits_exceptionVec_17 = io_writeback_21_bits_exceptionVec_17;
        //    mon_tr.io_writeback_21_bits_exceptionVec_18 = io_writeback_21_bits_exceptionVec_18;
        //    mon_tr.io_writeback_21_bits_exceptionVec_19 = io_writeback_21_bits_exceptionVec_19;
        //    mon_tr.io_writeback_21_bits_exceptionVec_20 = io_writeback_21_bits_exceptionVec_20;
        //    mon_tr.io_writeback_21_bits_exceptionVec_21 = io_writeback_21_bits_exceptionVec_21;
        //    mon_tr.io_writeback_21_bits_exceptionVec_22 = io_writeback_21_bits_exceptionVec_22;
        //    mon_tr.io_writeback_21_bits_exceptionVec_23 = io_writeback_21_bits_exceptionVec_23;
        //    mon_tr.io_writeback_21_bits_flushPipe = io_writeback_21_bits_flushPipe;
        //    mon_tr.io_writeback_21_bits_replay = io_writeback_21_bits_replay;
        //    mon_tr.io_writeback_21_bits_lqIdx_flag = io_writeback_21_bits_lqIdx_flag;
        //    mon_tr.io_writeback_21_bits_lqIdx_value = io_writeback_21_bits_lqIdx_value;
        //    mon_tr.io_writeback_21_bits_trigger = io_writeback_21_bits_trigger;
        //    mon_tr.io_writeback_21_bits_predecodeInfo_valid = io_writeback_21_bits_predecodeInfo_valid;
        //    mon_tr.io_writeback_21_bits_predecodeInfo_isRVC = io_writeback_21_bits_predecodeInfo_isRVC;
        //    mon_tr.io_writeback_21_bits_predecodeInfo_brType = io_writeback_21_bits_predecodeInfo_brType;
        //    mon_tr.io_writeback_21_bits_predecodeInfo_isCall = io_writeback_21_bits_predecodeInfo_isCall;
        //    mon_tr.io_writeback_21_bits_predecodeInfo_isRet = io_writeback_21_bits_predecodeInfo_isRet;
        //    mon_tr.io_writeback_21_bits_debug_isMMIO = io_writeback_21_bits_debug_isMMIO;
        //    mon_tr.io_writeback_21_bits_debug_isNCIO = io_writeback_21_bits_debug_isNCIO;
        //    mon_tr.io_writeback_21_bits_debug_isPerfCnt = io_writeback_21_bits_debug_isPerfCnt;
        //    mon_tr.io_writeback_21_bits_debug_paddr = io_writeback_21_bits_debug_paddr;
        //    mon_tr.io_writeback_21_bits_debug_vaddr = io_writeback_21_bits_debug_vaddr;
        //    mon_tr.io_writeback_21_bits_debugInfo_eliminatedMove = io_writeback_21_bits_debugInfo_eliminatedMove;
        //    mon_tr.io_writeback_21_bits_debugInfo_renameTime = io_writeback_21_bits_debugInfo_renameTime;
        //    mon_tr.io_writeback_21_bits_debugInfo_dispatchTime = io_writeback_21_bits_debugInfo_dispatchTime;
        //    mon_tr.io_writeback_21_bits_debugInfo_enqRsTime = io_writeback_21_bits_debugInfo_enqRsTime;
        //    mon_tr.io_writeback_21_bits_debugInfo_selectTime = io_writeback_21_bits_debugInfo_selectTime;
        //    mon_tr.io_writeback_21_bits_debugInfo_issueTime = io_writeback_21_bits_debugInfo_issueTime;
        //    mon_tr.io_writeback_21_bits_debugInfo_writebackTime = io_writeback_21_bits_debugInfo_writebackTime;
        //    mon_tr.io_writeback_21_bits_debugInfo_runahead_checkpoint_id = io_writeback_21_bits_debugInfo_runahead_checkpoint_id;
        //    mon_tr.io_writeback_21_bits_debugInfo_tlbFirstReqTime = io_writeback_21_bits_debugInfo_tlbFirstReqTime;
        //    mon_tr.io_writeback_21_bits_debugInfo_tlbRespTime = io_writeback_21_bits_debugInfo_tlbRespTime;
        //    mon_tr.io_writeback_21_bits_debug_seqNum = io_writeback_21_bits_debug_seqNum;
        //    mon_tr.io_writeback_20_valid = io_writeback_20_valid;
        //    mon_tr.io_writeback_20_bits_data_0 = io_writeback_20_bits_data_0;
        //    mon_tr.io_writeback_20_bits_pdest = io_writeback_20_bits_pdest;
        //    mon_tr.io_writeback_20_bits_robIdx_flag = io_writeback_20_bits_robIdx_flag;
        //    mon_tr.io_writeback_20_bits_robIdx_value = io_writeback_20_bits_robIdx_value;
        //    mon_tr.io_writeback_20_bits_intWen = io_writeback_20_bits_intWen;
        //    mon_tr.io_writeback_20_bits_fpWen = io_writeback_20_bits_fpWen;
        //    mon_tr.io_writeback_20_bits_exceptionVec_0 = io_writeback_20_bits_exceptionVec_0;
        //    mon_tr.io_writeback_20_bits_exceptionVec_1 = io_writeback_20_bits_exceptionVec_1;
        //    mon_tr.io_writeback_20_bits_exceptionVec_2 = io_writeback_20_bits_exceptionVec_2;
        //    mon_tr.io_writeback_20_bits_exceptionVec_3 = io_writeback_20_bits_exceptionVec_3;
        //    mon_tr.io_writeback_20_bits_exceptionVec_4 = io_writeback_20_bits_exceptionVec_4;
        //    mon_tr.io_writeback_20_bits_exceptionVec_5 = io_writeback_20_bits_exceptionVec_5;
        //    mon_tr.io_writeback_20_bits_exceptionVec_6 = io_writeback_20_bits_exceptionVec_6;
        //    mon_tr.io_writeback_20_bits_exceptionVec_7 = io_writeback_20_bits_exceptionVec_7;
        //    mon_tr.io_writeback_20_bits_exceptionVec_8 = io_writeback_20_bits_exceptionVec_8;
        //    mon_tr.io_writeback_20_bits_exceptionVec_9 = io_writeback_20_bits_exceptionVec_9;
        //    mon_tr.io_writeback_20_bits_exceptionVec_10 = io_writeback_20_bits_exceptionVec_10;
        //    mon_tr.io_writeback_20_bits_exceptionVec_11 = io_writeback_20_bits_exceptionVec_11;
        //    mon_tr.io_writeback_20_bits_exceptionVec_12 = io_writeback_20_bits_exceptionVec_12;
        //    mon_tr.io_writeback_20_bits_exceptionVec_13 = io_writeback_20_bits_exceptionVec_13;
        //    mon_tr.io_writeback_20_bits_exceptionVec_14 = io_writeback_20_bits_exceptionVec_14;
        //    mon_tr.io_writeback_20_bits_exceptionVec_15 = io_writeback_20_bits_exceptionVec_15;
        //    mon_tr.io_writeback_20_bits_exceptionVec_16 = io_writeback_20_bits_exceptionVec_16;
        //    mon_tr.io_writeback_20_bits_exceptionVec_17 = io_writeback_20_bits_exceptionVec_17;
        //    mon_tr.io_writeback_20_bits_exceptionVec_18 = io_writeback_20_bits_exceptionVec_18;
        //    mon_tr.io_writeback_20_bits_exceptionVec_19 = io_writeback_20_bits_exceptionVec_19;
        //    mon_tr.io_writeback_20_bits_exceptionVec_20 = io_writeback_20_bits_exceptionVec_20;
        //    mon_tr.io_writeback_20_bits_exceptionVec_21 = io_writeback_20_bits_exceptionVec_21;
        //    mon_tr.io_writeback_20_bits_exceptionVec_22 = io_writeback_20_bits_exceptionVec_22;
        //    mon_tr.io_writeback_20_bits_exceptionVec_23 = io_writeback_20_bits_exceptionVec_23;
        //    mon_tr.io_writeback_20_bits_flushPipe = io_writeback_20_bits_flushPipe;
        //    mon_tr.io_writeback_20_bits_replay = io_writeback_20_bits_replay;
        //    mon_tr.io_writeback_20_bits_lqIdx_flag = io_writeback_20_bits_lqIdx_flag;
        //    mon_tr.io_writeback_20_bits_lqIdx_value = io_writeback_20_bits_lqIdx_value;
        //    mon_tr.io_writeback_20_bits_trigger = io_writeback_20_bits_trigger;
        //    mon_tr.io_writeback_20_bits_predecodeInfo_valid = io_writeback_20_bits_predecodeInfo_valid;
        //    mon_tr.io_writeback_20_bits_predecodeInfo_isRVC = io_writeback_20_bits_predecodeInfo_isRVC;
        //    mon_tr.io_writeback_20_bits_predecodeInfo_brType = io_writeback_20_bits_predecodeInfo_brType;
        //    mon_tr.io_writeback_20_bits_predecodeInfo_isCall = io_writeback_20_bits_predecodeInfo_isCall;
        //    mon_tr.io_writeback_20_bits_predecodeInfo_isRet = io_writeback_20_bits_predecodeInfo_isRet;
        //    mon_tr.io_writeback_20_bits_debug_isMMIO = io_writeback_20_bits_debug_isMMIO;
        //    mon_tr.io_writeback_20_bits_debug_isNCIO = io_writeback_20_bits_debug_isNCIO;
        //    mon_tr.io_writeback_20_bits_debug_isPerfCnt = io_writeback_20_bits_debug_isPerfCnt;
        //    mon_tr.io_writeback_20_bits_debug_paddr = io_writeback_20_bits_debug_paddr;
        //    mon_tr.io_writeback_20_bits_debug_vaddr = io_writeback_20_bits_debug_vaddr;
        //    mon_tr.io_writeback_20_bits_debugInfo_eliminatedMove = io_writeback_20_bits_debugInfo_eliminatedMove;
        //    mon_tr.io_writeback_20_bits_debugInfo_renameTime = io_writeback_20_bits_debugInfo_renameTime;
        //    mon_tr.io_writeback_20_bits_debugInfo_dispatchTime = io_writeback_20_bits_debugInfo_dispatchTime;
        //    mon_tr.io_writeback_20_bits_debugInfo_enqRsTime = io_writeback_20_bits_debugInfo_enqRsTime;
        //    mon_tr.io_writeback_20_bits_debugInfo_selectTime = io_writeback_20_bits_debugInfo_selectTime;
        //    mon_tr.io_writeback_20_bits_debugInfo_issueTime = io_writeback_20_bits_debugInfo_issueTime;
        //    mon_tr.io_writeback_20_bits_debugInfo_writebackTime = io_writeback_20_bits_debugInfo_writebackTime;
        //    mon_tr.io_writeback_20_bits_debugInfo_runahead_checkpoint_id = io_writeback_20_bits_debugInfo_runahead_checkpoint_id;
        //    mon_tr.io_writeback_20_bits_debugInfo_tlbFirstReqTime = io_writeback_20_bits_debugInfo_tlbFirstReqTime;
        //    mon_tr.io_writeback_20_bits_debugInfo_tlbRespTime = io_writeback_20_bits_debugInfo_tlbRespTime;
        //    mon_tr.io_writeback_20_bits_debug_seqNum = io_writeback_20_bits_debug_seqNum;
        //    mon_tr.io_writeback_19_valid = io_writeback_19_valid;
        //    mon_tr.io_writeback_19_bits_data_0 = io_writeback_19_bits_data_0;
        //    mon_tr.io_writeback_19_bits_pdest = io_writeback_19_bits_pdest;
        //    mon_tr.io_writeback_19_bits_robIdx_flag = io_writeback_19_bits_robIdx_flag;
        //    mon_tr.io_writeback_19_bits_robIdx_value = io_writeback_19_bits_robIdx_value;
        //    mon_tr.io_writeback_19_bits_intWen = io_writeback_19_bits_intWen;
        //    mon_tr.io_writeback_19_bits_exceptionVec_0 = io_writeback_19_bits_exceptionVec_0;
        //    mon_tr.io_writeback_19_bits_exceptionVec_1 = io_writeback_19_bits_exceptionVec_1;
        //    mon_tr.io_writeback_19_bits_exceptionVec_2 = io_writeback_19_bits_exceptionVec_2;
        //    mon_tr.io_writeback_19_bits_exceptionVec_3 = io_writeback_19_bits_exceptionVec_3;
        //    mon_tr.io_writeback_19_bits_exceptionVec_4 = io_writeback_19_bits_exceptionVec_4;
        //    mon_tr.io_writeback_19_bits_exceptionVec_5 = io_writeback_19_bits_exceptionVec_5;
        //    mon_tr.io_writeback_19_bits_exceptionVec_6 = io_writeback_19_bits_exceptionVec_6;
        //    mon_tr.io_writeback_19_bits_exceptionVec_7 = io_writeback_19_bits_exceptionVec_7;
        //    mon_tr.io_writeback_19_bits_exceptionVec_8 = io_writeback_19_bits_exceptionVec_8;
        //    mon_tr.io_writeback_19_bits_exceptionVec_9 = io_writeback_19_bits_exceptionVec_9;
        //    mon_tr.io_writeback_19_bits_exceptionVec_10 = io_writeback_19_bits_exceptionVec_10;
        //    mon_tr.io_writeback_19_bits_exceptionVec_11 = io_writeback_19_bits_exceptionVec_11;
        //    mon_tr.io_writeback_19_bits_exceptionVec_12 = io_writeback_19_bits_exceptionVec_12;
        //    mon_tr.io_writeback_19_bits_exceptionVec_13 = io_writeback_19_bits_exceptionVec_13;
        //    mon_tr.io_writeback_19_bits_exceptionVec_14 = io_writeback_19_bits_exceptionVec_14;
        //    mon_tr.io_writeback_19_bits_exceptionVec_15 = io_writeback_19_bits_exceptionVec_15;
        //    mon_tr.io_writeback_19_bits_exceptionVec_16 = io_writeback_19_bits_exceptionVec_16;
        //    mon_tr.io_writeback_19_bits_exceptionVec_17 = io_writeback_19_bits_exceptionVec_17;
        //    mon_tr.io_writeback_19_bits_exceptionVec_18 = io_writeback_19_bits_exceptionVec_18;
        //    mon_tr.io_writeback_19_bits_exceptionVec_19 = io_writeback_19_bits_exceptionVec_19;
        //    mon_tr.io_writeback_19_bits_exceptionVec_20 = io_writeback_19_bits_exceptionVec_20;
        //    mon_tr.io_writeback_19_bits_exceptionVec_21 = io_writeback_19_bits_exceptionVec_21;
        //    mon_tr.io_writeback_19_bits_exceptionVec_22 = io_writeback_19_bits_exceptionVec_22;
        //    mon_tr.io_writeback_19_bits_exceptionVec_23 = io_writeback_19_bits_exceptionVec_23;
        //    mon_tr.io_writeback_19_bits_flushPipe = io_writeback_19_bits_flushPipe;
        //    mon_tr.io_writeback_19_bits_sqIdx_flag = io_writeback_19_bits_sqIdx_flag;
        //    mon_tr.io_writeback_19_bits_sqIdx_value = io_writeback_19_bits_sqIdx_value;
        //    mon_tr.io_writeback_19_bits_trigger = io_writeback_19_bits_trigger;
        //    mon_tr.io_writeback_19_bits_debug_isMMIO = io_writeback_19_bits_debug_isMMIO;
        //    mon_tr.io_writeback_19_bits_debug_isNCIO = io_writeback_19_bits_debug_isNCIO;
        //    mon_tr.io_writeback_19_bits_debug_isPerfCnt = io_writeback_19_bits_debug_isPerfCnt;
        //    mon_tr.io_writeback_19_bits_debug_paddr = io_writeback_19_bits_debug_paddr;
        //    mon_tr.io_writeback_19_bits_debug_vaddr = io_writeback_19_bits_debug_vaddr;
        //    mon_tr.io_writeback_19_bits_debugInfo_eliminatedMove = io_writeback_19_bits_debugInfo_eliminatedMove;
        //    mon_tr.io_writeback_19_bits_debugInfo_renameTime = io_writeback_19_bits_debugInfo_renameTime;
        //    mon_tr.io_writeback_19_bits_debugInfo_dispatchTime = io_writeback_19_bits_debugInfo_dispatchTime;
        //    mon_tr.io_writeback_19_bits_debugInfo_enqRsTime = io_writeback_19_bits_debugInfo_enqRsTime;
        //    mon_tr.io_writeback_19_bits_debugInfo_selectTime = io_writeback_19_bits_debugInfo_selectTime;
        //    mon_tr.io_writeback_19_bits_debugInfo_issueTime = io_writeback_19_bits_debugInfo_issueTime;
        //    mon_tr.io_writeback_19_bits_debugInfo_writebackTime = io_writeback_19_bits_debugInfo_writebackTime;
        //    mon_tr.io_writeback_19_bits_debugInfo_runahead_checkpoint_id = io_writeback_19_bits_debugInfo_runahead_checkpoint_id;
        //    mon_tr.io_writeback_19_bits_debugInfo_tlbFirstReqTime = io_writeback_19_bits_debugInfo_tlbFirstReqTime;
        //    mon_tr.io_writeback_19_bits_debugInfo_tlbRespTime = io_writeback_19_bits_debugInfo_tlbRespTime;
        //    mon_tr.io_writeback_19_bits_debug_seqNum = io_writeback_19_bits_debug_seqNum;
        //    mon_tr.io_writeback_18_valid = io_writeback_18_valid;
        //    mon_tr.io_writeback_18_bits_data_0 = io_writeback_18_bits_data_0;
        //    mon_tr.io_writeback_18_bits_pdest = io_writeback_18_bits_pdest;
        //    mon_tr.io_writeback_18_bits_robIdx_flag = io_writeback_18_bits_robIdx_flag;
        //    mon_tr.io_writeback_18_bits_robIdx_value = io_writeback_18_bits_robIdx_value;
        //    mon_tr.io_writeback_18_bits_intWen = io_writeback_18_bits_intWen;
        //    mon_tr.io_writeback_18_bits_exceptionVec_0 = io_writeback_18_bits_exceptionVec_0;
        //    mon_tr.io_writeback_18_bits_exceptionVec_1 = io_writeback_18_bits_exceptionVec_1;
        //    mon_tr.io_writeback_18_bits_exceptionVec_2 = io_writeback_18_bits_exceptionVec_2;
        //    mon_tr.io_writeback_18_bits_exceptionVec_3 = io_writeback_18_bits_exceptionVec_3;
        //    mon_tr.io_writeback_18_bits_exceptionVec_4 = io_writeback_18_bits_exceptionVec_4;
        //    mon_tr.io_writeback_18_bits_exceptionVec_5 = io_writeback_18_bits_exceptionVec_5;
        //    mon_tr.io_writeback_18_bits_exceptionVec_6 = io_writeback_18_bits_exceptionVec_6;
        //    mon_tr.io_writeback_18_bits_exceptionVec_7 = io_writeback_18_bits_exceptionVec_7;
        //    mon_tr.io_writeback_18_bits_exceptionVec_8 = io_writeback_18_bits_exceptionVec_8;
        //    mon_tr.io_writeback_18_bits_exceptionVec_9 = io_writeback_18_bits_exceptionVec_9;
        //    mon_tr.io_writeback_18_bits_exceptionVec_10 = io_writeback_18_bits_exceptionVec_10;
        //    mon_tr.io_writeback_18_bits_exceptionVec_11 = io_writeback_18_bits_exceptionVec_11;
        //    mon_tr.io_writeback_18_bits_exceptionVec_12 = io_writeback_18_bits_exceptionVec_12;
        //    mon_tr.io_writeback_18_bits_exceptionVec_13 = io_writeback_18_bits_exceptionVec_13;
        //    mon_tr.io_writeback_18_bits_exceptionVec_14 = io_writeback_18_bits_exceptionVec_14;
        //    mon_tr.io_writeback_18_bits_exceptionVec_15 = io_writeback_18_bits_exceptionVec_15;
        //    mon_tr.io_writeback_18_bits_exceptionVec_16 = io_writeback_18_bits_exceptionVec_16;
        //    mon_tr.io_writeback_18_bits_exceptionVec_17 = io_writeback_18_bits_exceptionVec_17;
        //    mon_tr.io_writeback_18_bits_exceptionVec_18 = io_writeback_18_bits_exceptionVec_18;
        //    mon_tr.io_writeback_18_bits_exceptionVec_19 = io_writeback_18_bits_exceptionVec_19;
        //    mon_tr.io_writeback_18_bits_exceptionVec_20 = io_writeback_18_bits_exceptionVec_20;
        //    mon_tr.io_writeback_18_bits_exceptionVec_21 = io_writeback_18_bits_exceptionVec_21;
        //    mon_tr.io_writeback_18_bits_exceptionVec_22 = io_writeback_18_bits_exceptionVec_22;
        //    mon_tr.io_writeback_18_bits_exceptionVec_23 = io_writeback_18_bits_exceptionVec_23;
        //    mon_tr.io_writeback_18_bits_flushPipe = io_writeback_18_bits_flushPipe;
        //    mon_tr.io_writeback_18_bits_sqIdx_flag = io_writeback_18_bits_sqIdx_flag;
        //    mon_tr.io_writeback_18_bits_sqIdx_value = io_writeback_18_bits_sqIdx_value;
        //    mon_tr.io_writeback_18_bits_trigger = io_writeback_18_bits_trigger;
        //    mon_tr.io_writeback_18_bits_debug_isMMIO = io_writeback_18_bits_debug_isMMIO;
        //    mon_tr.io_writeback_18_bits_debug_isNCIO = io_writeback_18_bits_debug_isNCIO;
        //    mon_tr.io_writeback_18_bits_debug_isPerfCnt = io_writeback_18_bits_debug_isPerfCnt;
        //    mon_tr.io_writeback_18_bits_debug_paddr = io_writeback_18_bits_debug_paddr;
        //    mon_tr.io_writeback_18_bits_debug_vaddr = io_writeback_18_bits_debug_vaddr;
        //    mon_tr.io_writeback_18_bits_debugInfo_eliminatedMove = io_writeback_18_bits_debugInfo_eliminatedMove;
        //    mon_tr.io_writeback_18_bits_debugInfo_renameTime = io_writeback_18_bits_debugInfo_renameTime;
        //    mon_tr.io_writeback_18_bits_debugInfo_dispatchTime = io_writeback_18_bits_debugInfo_dispatchTime;
        //    mon_tr.io_writeback_18_bits_debugInfo_enqRsTime = io_writeback_18_bits_debugInfo_enqRsTime;
        //    mon_tr.io_writeback_18_bits_debugInfo_selectTime = io_writeback_18_bits_debugInfo_selectTime;
        //    mon_tr.io_writeback_18_bits_debugInfo_issueTime = io_writeback_18_bits_debugInfo_issueTime;
        //    mon_tr.io_writeback_18_bits_debugInfo_writebackTime = io_writeback_18_bits_debugInfo_writebackTime;
        //    mon_tr.io_writeback_18_bits_debugInfo_runahead_checkpoint_id = io_writeback_18_bits_debugInfo_runahead_checkpoint_id;
        //    mon_tr.io_writeback_18_bits_debugInfo_tlbFirstReqTime = io_writeback_18_bits_debugInfo_tlbFirstReqTime;
        //    mon_tr.io_writeback_18_bits_debugInfo_tlbRespTime = io_writeback_18_bits_debugInfo_tlbRespTime;
        //    mon_tr.io_writeback_18_bits_debug_seqNum = io_writeback_18_bits_debug_seqNum;
        //    mon_tr.io_writeback_17_valid = io_writeback_17_valid;
        //    mon_tr.io_writeback_17_bits_data_0 = io_writeback_17_bits_data_0;
        //    mon_tr.io_writeback_17_bits_data_1 = io_writeback_17_bits_data_1;
        //    mon_tr.io_writeback_17_bits_data_2 = io_writeback_17_bits_data_2;
        //    mon_tr.io_writeback_17_bits_pdest = io_writeback_17_bits_pdest;
        //    mon_tr.io_writeback_17_bits_robIdx_flag = io_writeback_17_bits_robIdx_flag;
        //    mon_tr.io_writeback_17_bits_robIdx_value = io_writeback_17_bits_robIdx_value;
        //    mon_tr.io_writeback_17_bits_vecWen = io_writeback_17_bits_vecWen;
        //    mon_tr.io_writeback_17_bits_v0Wen = io_writeback_17_bits_v0Wen;
        //    mon_tr.io_writeback_17_bits_fflags = io_writeback_17_bits_fflags;
        //    mon_tr.io_writeback_17_bits_wflags = io_writeback_17_bits_wflags;
        //    mon_tr.io_writeback_17_bits_debugInfo_eliminatedMove = io_writeback_17_bits_debugInfo_eliminatedMove;
        //    mon_tr.io_writeback_17_bits_debugInfo_renameTime = io_writeback_17_bits_debugInfo_renameTime;
        //    mon_tr.io_writeback_17_bits_debugInfo_dispatchTime = io_writeback_17_bits_debugInfo_dispatchTime;
        //    mon_tr.io_writeback_17_bits_debugInfo_enqRsTime = io_writeback_17_bits_debugInfo_enqRsTime;
        //    mon_tr.io_writeback_17_bits_debugInfo_selectTime = io_writeback_17_bits_debugInfo_selectTime;
        //    mon_tr.io_writeback_17_bits_debugInfo_issueTime = io_writeback_17_bits_debugInfo_issueTime;
        //    mon_tr.io_writeback_17_bits_debugInfo_writebackTime = io_writeback_17_bits_debugInfo_writebackTime;
        //    mon_tr.io_writeback_17_bits_debugInfo_runahead_checkpoint_id = io_writeback_17_bits_debugInfo_runahead_checkpoint_id;
        //    mon_tr.io_writeback_17_bits_debugInfo_tlbFirstReqTime = io_writeback_17_bits_debugInfo_tlbFirstReqTime;
        //    mon_tr.io_writeback_17_bits_debugInfo_tlbRespTime = io_writeback_17_bits_debugInfo_tlbRespTime;
        //    mon_tr.io_writeback_17_bits_debug_seqNum = io_writeback_17_bits_debug_seqNum;
        //    mon_tr.io_writeback_16_valid = io_writeback_16_valid;
        //    mon_tr.io_writeback_16_bits_data_0 = io_writeback_16_bits_data_0;
        //    mon_tr.io_writeback_16_bits_data_1 = io_writeback_16_bits_data_1;
        //    mon_tr.io_writeback_16_bits_data_2 = io_writeback_16_bits_data_2;
        //    mon_tr.io_writeback_16_bits_data_3 = io_writeback_16_bits_data_3;
        //    mon_tr.io_writeback_16_bits_pdest = io_writeback_16_bits_pdest;
        //    mon_tr.io_writeback_16_bits_robIdx_flag = io_writeback_16_bits_robIdx_flag;
        //    mon_tr.io_writeback_16_bits_robIdx_value = io_writeback_16_bits_robIdx_value;
        //    mon_tr.io_writeback_16_bits_fpWen = io_writeback_16_bits_fpWen;
        //    mon_tr.io_writeback_16_bits_vecWen = io_writeback_16_bits_vecWen;
        //    mon_tr.io_writeback_16_bits_v0Wen = io_writeback_16_bits_v0Wen;
        //    mon_tr.io_writeback_16_bits_fflags = io_writeback_16_bits_fflags;
        //    mon_tr.io_writeback_16_bits_wflags = io_writeback_16_bits_wflags;
        //    mon_tr.io_writeback_16_bits_debugInfo_eliminatedMove = io_writeback_16_bits_debugInfo_eliminatedMove;
        //    mon_tr.io_writeback_16_bits_debugInfo_renameTime = io_writeback_16_bits_debugInfo_renameTime;
        //    mon_tr.io_writeback_16_bits_debugInfo_dispatchTime = io_writeback_16_bits_debugInfo_dispatchTime;
        //    mon_tr.io_writeback_16_bits_debugInfo_enqRsTime = io_writeback_16_bits_debugInfo_enqRsTime;
        //    mon_tr.io_writeback_16_bits_debugInfo_selectTime = io_writeback_16_bits_debugInfo_selectTime;
        //    mon_tr.io_writeback_16_bits_debugInfo_issueTime = io_writeback_16_bits_debugInfo_issueTime;
        //    mon_tr.io_writeback_16_bits_debugInfo_writebackTime = io_writeback_16_bits_debugInfo_writebackTime;
        //    mon_tr.io_writeback_16_bits_debugInfo_runahead_checkpoint_id = io_writeback_16_bits_debugInfo_runahead_checkpoint_id;
        //    mon_tr.io_writeback_16_bits_debugInfo_tlbFirstReqTime = io_writeback_16_bits_debugInfo_tlbFirstReqTime;
        //    mon_tr.io_writeback_16_bits_debugInfo_tlbRespTime = io_writeback_16_bits_debugInfo_tlbRespTime;
        //    mon_tr.io_writeback_16_bits_debug_seqNum = io_writeback_16_bits_debug_seqNum;
        //    mon_tr.io_writeback_15_valid = io_writeback_15_valid;
        //    mon_tr.io_writeback_15_bits_data_0 = io_writeback_15_bits_data_0;
        //    mon_tr.io_writeback_15_bits_data_1 = io_writeback_15_bits_data_1;
        //    mon_tr.io_writeback_15_bits_data_2 = io_writeback_15_bits_data_2;
        //    mon_tr.io_writeback_15_bits_pdest = io_writeback_15_bits_pdest;
        //    mon_tr.io_writeback_15_bits_robIdx_flag = io_writeback_15_bits_robIdx_flag;
        //    mon_tr.io_writeback_15_bits_robIdx_value = io_writeback_15_bits_robIdx_value;
        //    mon_tr.io_writeback_15_bits_vecWen = io_writeback_15_bits_vecWen;
        //    mon_tr.io_writeback_15_bits_v0Wen = io_writeback_15_bits_v0Wen;
        //    mon_tr.io_writeback_15_bits_fflags = io_writeback_15_bits_fflags;
        //    mon_tr.io_writeback_15_bits_wflags = io_writeback_15_bits_wflags;
        //    mon_tr.io_writeback_15_bits_vxsat = io_writeback_15_bits_vxsat;
        //    mon_tr.io_writeback_15_bits_debugInfo_eliminatedMove = io_writeback_15_bits_debugInfo_eliminatedMove;
        //    mon_tr.io_writeback_15_bits_debugInfo_renameTime = io_writeback_15_bits_debugInfo_renameTime;
        //    mon_tr.io_writeback_15_bits_debugInfo_dispatchTime = io_writeback_15_bits_debugInfo_dispatchTime;
        //    mon_tr.io_writeback_15_bits_debugInfo_enqRsTime = io_writeback_15_bits_debugInfo_enqRsTime;
        //    mon_tr.io_writeback_15_bits_debugInfo_selectTime = io_writeback_15_bits_debugInfo_selectTime;
        //    mon_tr.io_writeback_15_bits_debugInfo_issueTime = io_writeback_15_bits_debugInfo_issueTime;
        //    mon_tr.io_writeback_15_bits_debugInfo_writebackTime = io_writeback_15_bits_debugInfo_writebackTime;
        //    mon_tr.io_writeback_15_bits_debugInfo_runahead_checkpoint_id = io_writeback_15_bits_debugInfo_runahead_checkpoint_id;
        //    mon_tr.io_writeback_15_bits_debugInfo_tlbFirstReqTime = io_writeback_15_bits_debugInfo_tlbFirstReqTime;
        //    mon_tr.io_writeback_15_bits_debugInfo_tlbRespTime = io_writeback_15_bits_debugInfo_tlbRespTime;
        //    mon_tr.io_writeback_15_bits_debug_seqNum = io_writeback_15_bits_debug_seqNum;
        //    mon_tr.io_writeback_14_valid = io_writeback_14_valid;
        //    mon_tr.io_writeback_14_bits_data_0 = io_writeback_14_bits_data_0;
        //    mon_tr.io_writeback_14_bits_data_1 = io_writeback_14_bits_data_1;
        //    mon_tr.io_writeback_14_bits_data_2 = io_writeback_14_bits_data_2;
        //    mon_tr.io_writeback_14_bits_data_3 = io_writeback_14_bits_data_3;
        //    mon_tr.io_writeback_14_bits_data_4 = io_writeback_14_bits_data_4;
        //    mon_tr.io_writeback_14_bits_data_5 = io_writeback_14_bits_data_5;
        //    mon_tr.io_writeback_14_bits_pdest = io_writeback_14_bits_pdest;
        //    mon_tr.io_writeback_14_bits_robIdx_flag = io_writeback_14_bits_robIdx_flag;
        //    mon_tr.io_writeback_14_bits_robIdx_value = io_writeback_14_bits_robIdx_value;
        //    mon_tr.io_writeback_14_bits_intWen = io_writeback_14_bits_intWen;
        //    mon_tr.io_writeback_14_bits_fpWen = io_writeback_14_bits_fpWen;
        //    mon_tr.io_writeback_14_bits_vecWen = io_writeback_14_bits_vecWen;
        //    mon_tr.io_writeback_14_bits_v0Wen = io_writeback_14_bits_v0Wen;
        //    mon_tr.io_writeback_14_bits_vlWen = io_writeback_14_bits_vlWen;
        //    mon_tr.io_writeback_14_bits_fflags = io_writeback_14_bits_fflags;
        //    mon_tr.io_writeback_14_bits_wflags = io_writeback_14_bits_wflags;
        //    mon_tr.io_writeback_14_bits_exceptionVec_2 = io_writeback_14_bits_exceptionVec_2;
        //    mon_tr.io_writeback_14_bits_debugInfo_eliminatedMove = io_writeback_14_bits_debugInfo_eliminatedMove;
        //    mon_tr.io_writeback_14_bits_debugInfo_renameTime = io_writeback_14_bits_debugInfo_renameTime;
        //    mon_tr.io_writeback_14_bits_debugInfo_dispatchTime = io_writeback_14_bits_debugInfo_dispatchTime;
        //    mon_tr.io_writeback_14_bits_debugInfo_enqRsTime = io_writeback_14_bits_debugInfo_enqRsTime;
        //    mon_tr.io_writeback_14_bits_debugInfo_selectTime = io_writeback_14_bits_debugInfo_selectTime;
        //    mon_tr.io_writeback_14_bits_debugInfo_issueTime = io_writeback_14_bits_debugInfo_issueTime;
        //    mon_tr.io_writeback_14_bits_debugInfo_writebackTime = io_writeback_14_bits_debugInfo_writebackTime;
        //    mon_tr.io_writeback_14_bits_debugInfo_runahead_checkpoint_id = io_writeback_14_bits_debugInfo_runahead_checkpoint_id;
        //    mon_tr.io_writeback_14_bits_debugInfo_tlbFirstReqTime = io_writeback_14_bits_debugInfo_tlbFirstReqTime;
        //    mon_tr.io_writeback_14_bits_debugInfo_tlbRespTime = io_writeback_14_bits_debugInfo_tlbRespTime;
        //    mon_tr.io_writeback_14_bits_debug_seqNum = io_writeback_14_bits_debug_seqNum;
        //    mon_tr.io_writeback_13_valid = io_writeback_13_valid;
        //    mon_tr.io_writeback_13_bits_data_0 = io_writeback_13_bits_data_0;
        //    mon_tr.io_writeback_13_bits_data_1 = io_writeback_13_bits_data_1;
        //    mon_tr.io_writeback_13_bits_data_2 = io_writeback_13_bits_data_2;
        //    mon_tr.io_writeback_13_bits_pdest = io_writeback_13_bits_pdest;
        //    mon_tr.io_writeback_13_bits_robIdx_flag = io_writeback_13_bits_robIdx_flag;
        //    mon_tr.io_writeback_13_bits_robIdx_value = io_writeback_13_bits_robIdx_value;
        //    mon_tr.io_writeback_13_bits_vecWen = io_writeback_13_bits_vecWen;
        //    mon_tr.io_writeback_13_bits_v0Wen = io_writeback_13_bits_v0Wen;
        //    mon_tr.io_writeback_13_bits_fflags = io_writeback_13_bits_fflags;
        //    mon_tr.io_writeback_13_bits_wflags = io_writeback_13_bits_wflags;
        //    mon_tr.io_writeback_13_bits_vxsat = io_writeback_13_bits_vxsat;
        //    mon_tr.io_writeback_13_bits_exceptionVec_2 = io_writeback_13_bits_exceptionVec_2;
        //    mon_tr.io_writeback_13_bits_debugInfo_eliminatedMove = io_writeback_13_bits_debugInfo_eliminatedMove;
        //    mon_tr.io_writeback_13_bits_debugInfo_renameTime = io_writeback_13_bits_debugInfo_renameTime;
        //    mon_tr.io_writeback_13_bits_debugInfo_dispatchTime = io_writeback_13_bits_debugInfo_dispatchTime;
        //    mon_tr.io_writeback_13_bits_debugInfo_enqRsTime = io_writeback_13_bits_debugInfo_enqRsTime;
        //    mon_tr.io_writeback_13_bits_debugInfo_selectTime = io_writeback_13_bits_debugInfo_selectTime;
        //    mon_tr.io_writeback_13_bits_debugInfo_issueTime = io_writeback_13_bits_debugInfo_issueTime;
        //    mon_tr.io_writeback_13_bits_debugInfo_writebackTime = io_writeback_13_bits_debugInfo_writebackTime;
        //    mon_tr.io_writeback_13_bits_debugInfo_runahead_checkpoint_id = io_writeback_13_bits_debugInfo_runahead_checkpoint_id;
        //    mon_tr.io_writeback_13_bits_debugInfo_tlbFirstReqTime = io_writeback_13_bits_debugInfo_tlbFirstReqTime;
        //    mon_tr.io_writeback_13_bits_debugInfo_tlbRespTime = io_writeback_13_bits_debugInfo_tlbRespTime;
        //    mon_tr.io_writeback_13_bits_debug_seqNum = io_writeback_13_bits_debug_seqNum;
        //    mon_tr.io_writeback_7_valid = io_writeback_7_valid;
        //    mon_tr.io_writeback_7_bits_data_0 = io_writeback_7_bits_data_0;
        //    mon_tr.io_writeback_7_bits_data_1 = io_writeback_7_bits_data_1;
        //    mon_tr.io_writeback_7_bits_pdest = io_writeback_7_bits_pdest;
        //    mon_tr.io_writeback_7_bits_robIdx_flag = io_writeback_7_bits_robIdx_flag;
        //    mon_tr.io_writeback_7_bits_robIdx_value = io_writeback_7_bits_robIdx_value;
        //    mon_tr.io_writeback_7_bits_intWen = io_writeback_7_bits_intWen;
        //    mon_tr.io_writeback_7_bits_redirect_valid = io_writeback_7_bits_redirect_valid;
        //    mon_tr.io_writeback_7_bits_redirect_bits_isRVC = io_writeback_7_bits_redirect_bits_isRVC;
        //    mon_tr.io_writeback_7_bits_redirect_bits_robIdx_flag = io_writeback_7_bits_redirect_bits_robIdx_flag;
        //    mon_tr.io_writeback_7_bits_redirect_bits_robIdx_value = io_writeback_7_bits_redirect_bits_robIdx_value;
        //    mon_tr.io_writeback_7_bits_redirect_bits_ftqIdx_flag = io_writeback_7_bits_redirect_bits_ftqIdx_flag;
        //    mon_tr.io_writeback_7_bits_redirect_bits_ftqIdx_value = io_writeback_7_bits_redirect_bits_ftqIdx_value;
        //    mon_tr.io_writeback_7_bits_redirect_bits_ftqOffset = io_writeback_7_bits_redirect_bits_ftqOffset;
        //    mon_tr.io_writeback_7_bits_redirect_bits_level = io_writeback_7_bits_redirect_bits_level;
        //    mon_tr.io_writeback_7_bits_redirect_bits_interrupt = io_writeback_7_bits_redirect_bits_interrupt;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_pc = io_writeback_7_bits_redirect_bits_cfiUpdate_pc;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid = io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC = io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType = io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall = io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet = io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_ssp = io_writeback_7_bits_redirect_bits_cfiUpdate_ssp;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_sctr = io_writeback_7_bits_redirect_bits_cfiUpdate_sctr;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag = io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value = io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag = io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value = io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag = io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value = io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr = io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist = io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist = io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist = io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist = io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist = io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist = io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist = io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist = io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist = io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist = io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist = io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist = io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist = io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist = io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist = io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist = io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist = io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist = io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0 = io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1 = io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2 = io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3 = io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0 = io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1 = io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2 = io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3 = io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0 = io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1 = io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2 = io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3 = io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0 = io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1 = io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2 = io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3 = io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0 = io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1 = io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2 = io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3 = io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0 = io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1 = io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2 = io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3 = io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH = io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_ghr = io_writeback_7_bits_redirect_bits_cfiUpdate_ghr;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag = io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value = io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0 = io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1 = io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit = io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit = io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit = io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken = io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_target = io_writeback_7_bits_redirect_bits_cfiUpdate_target;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_taken = io_writeback_7_bits_redirect_bits_cfiUpdate_taken;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred = io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_shift = io_writeback_7_bits_redirect_bits_cfiUpdate_shift;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist = io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF = io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF = io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF;
        //    mon_tr.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF = io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF;
        //    mon_tr.io_writeback_7_bits_redirect_bits_fullTarget = io_writeback_7_bits_redirect_bits_fullTarget;
        //    mon_tr.io_writeback_7_bits_redirect_bits_stFtqIdx_flag = io_writeback_7_bits_redirect_bits_stFtqIdx_flag;
        //    mon_tr.io_writeback_7_bits_redirect_bits_stFtqIdx_value = io_writeback_7_bits_redirect_bits_stFtqIdx_value;
        //    mon_tr.io_writeback_7_bits_redirect_bits_stFtqOffset = io_writeback_7_bits_redirect_bits_stFtqOffset;
        //    mon_tr.io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id = io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id;
        //    mon_tr.io_writeback_7_bits_redirect_bits_debugIsCtrl = io_writeback_7_bits_redirect_bits_debugIsCtrl;
        //    mon_tr.io_writeback_7_bits_redirect_bits_debugIsMemVio = io_writeback_7_bits_redirect_bits_debugIsMemVio;
        //    mon_tr.io_writeback_7_bits_exceptionVec_2 = io_writeback_7_bits_exceptionVec_2;
        //    mon_tr.io_writeback_7_bits_exceptionVec_3 = io_writeback_7_bits_exceptionVec_3;
        //    mon_tr.io_writeback_7_bits_exceptionVec_8 = io_writeback_7_bits_exceptionVec_8;
        //    mon_tr.io_writeback_7_bits_exceptionVec_9 = io_writeback_7_bits_exceptionVec_9;
        //    mon_tr.io_writeback_7_bits_exceptionVec_10 = io_writeback_7_bits_exceptionVec_10;
        //    mon_tr.io_writeback_7_bits_exceptionVec_11 = io_writeback_7_bits_exceptionVec_11;
        //    mon_tr.io_writeback_7_bits_exceptionVec_22 = io_writeback_7_bits_exceptionVec_22;
        //    mon_tr.io_writeback_7_bits_flushPipe = io_writeback_7_bits_flushPipe;
        //    mon_tr.io_writeback_7_bits_predecodeInfo_valid = io_writeback_7_bits_predecodeInfo_valid;
        //    mon_tr.io_writeback_7_bits_predecodeInfo_isRVC = io_writeback_7_bits_predecodeInfo_isRVC;
        //    mon_tr.io_writeback_7_bits_predecodeInfo_brType = io_writeback_7_bits_predecodeInfo_brType;
        //    mon_tr.io_writeback_7_bits_predecodeInfo_isCall = io_writeback_7_bits_predecodeInfo_isCall;
        //    mon_tr.io_writeback_7_bits_predecodeInfo_isRet = io_writeback_7_bits_predecodeInfo_isRet;
        //    mon_tr.io_writeback_7_bits_debug_isPerfCnt = io_writeback_7_bits_debug_isPerfCnt;
        //    mon_tr.io_writeback_7_bits_debugInfo_eliminatedMove = io_writeback_7_bits_debugInfo_eliminatedMove;
        //    mon_tr.io_writeback_7_bits_debugInfo_renameTime = io_writeback_7_bits_debugInfo_renameTime;
        //    mon_tr.io_writeback_7_bits_debugInfo_dispatchTime = io_writeback_7_bits_debugInfo_dispatchTime;
        //    mon_tr.io_writeback_7_bits_debugInfo_enqRsTime = io_writeback_7_bits_debugInfo_enqRsTime;
        //    mon_tr.io_writeback_7_bits_debugInfo_selectTime = io_writeback_7_bits_debugInfo_selectTime;
        //    mon_tr.io_writeback_7_bits_debugInfo_issueTime = io_writeback_7_bits_debugInfo_issueTime;
        //    mon_tr.io_writeback_7_bits_debugInfo_writebackTime = io_writeback_7_bits_debugInfo_writebackTime;
        //    mon_tr.io_writeback_7_bits_debugInfo_runahead_checkpoint_id = io_writeback_7_bits_debugInfo_runahead_checkpoint_id;
        //    mon_tr.io_writeback_7_bits_debugInfo_tlbFirstReqTime = io_writeback_7_bits_debugInfo_tlbFirstReqTime;
        //    mon_tr.io_writeback_7_bits_debugInfo_tlbRespTime = io_writeback_7_bits_debugInfo_tlbRespTime;
        //    mon_tr.io_writeback_7_bits_debug_seqNum = io_writeback_7_bits_debug_seqNum;
        //    mon_tr.io_writeback_5_valid = io_writeback_5_valid;
        //    mon_tr.io_writeback_5_bits_redirect_valid = io_writeback_5_bits_redirect_valid;
        //    mon_tr.io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred = io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred;
        //    mon_tr.io_writeback_3_valid = io_writeback_3_valid;
        //    mon_tr.io_writeback_3_bits_redirect_valid = io_writeback_3_bits_redirect_valid;
        //    mon_tr.io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred = io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred;
        //    mon_tr.io_writeback_1_valid = io_writeback_1_valid;
        //    mon_tr.io_writeback_1_bits_redirect_valid = io_writeback_1_bits_redirect_valid;
        //    mon_tr.io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred = io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred;
        //    mon_tr.io_exuWriteback_26_valid = io_exuWriteback_26_valid;
        //    mon_tr.io_exuWriteback_26_bits_robIdx_value = io_exuWriteback_26_bits_robIdx_value;
        //    mon_tr.io_exuWriteback_25_valid = io_exuWriteback_25_valid;
        //    mon_tr.io_exuWriteback_25_bits_robIdx_value = io_exuWriteback_25_bits_robIdx_value;
        //    mon_tr.io_exuWriteback_24_valid = io_exuWriteback_24_valid;
        //    mon_tr.io_exuWriteback_24_bits_data_0 = io_exuWriteback_24_bits_data_0;
        //    mon_tr.io_exuWriteback_24_bits_pdest = io_exuWriteback_24_bits_pdest;
        //    mon_tr.io_exuWriteback_24_bits_robIdx_value = io_exuWriteback_24_bits_robIdx_value;
        //    mon_tr.io_exuWriteback_24_bits_vecWen = io_exuWriteback_24_bits_vecWen;
        //    mon_tr.io_exuWriteback_24_bits_v0Wen = io_exuWriteback_24_bits_v0Wen;
        //    mon_tr.io_exuWriteback_24_bits_vls_vdIdx = io_exuWriteback_24_bits_vls_vdIdx;
        //    mon_tr.io_exuWriteback_24_bits_debug_isMMIO = io_exuWriteback_24_bits_debug_isMMIO;
        //    mon_tr.io_exuWriteback_24_bits_debug_isNCIO = io_exuWriteback_24_bits_debug_isNCIO;
        //    mon_tr.io_exuWriteback_24_bits_debug_isPerfCnt = io_exuWriteback_24_bits_debug_isPerfCnt;
        //    mon_tr.io_exuWriteback_24_bits_debug_paddr = io_exuWriteback_24_bits_debug_paddr;
        //    mon_tr.io_exuWriteback_23_valid = io_exuWriteback_23_valid;
        //    mon_tr.io_exuWriteback_23_bits_data_0 = io_exuWriteback_23_bits_data_0;
        //    mon_tr.io_exuWriteback_23_bits_pdest = io_exuWriteback_23_bits_pdest;
        //    mon_tr.io_exuWriteback_23_bits_robIdx_value = io_exuWriteback_23_bits_robIdx_value;
        //    mon_tr.io_exuWriteback_23_bits_vecWen = io_exuWriteback_23_bits_vecWen;
        //    mon_tr.io_exuWriteback_23_bits_v0Wen = io_exuWriteback_23_bits_v0Wen;
        //    mon_tr.io_exuWriteback_23_bits_vls_vdIdx = io_exuWriteback_23_bits_vls_vdIdx;
        //    mon_tr.io_exuWriteback_23_bits_debug_isMMIO = io_exuWriteback_23_bits_debug_isMMIO;
        //    mon_tr.io_exuWriteback_23_bits_debug_isNCIO = io_exuWriteback_23_bits_debug_isNCIO;
        //    mon_tr.io_exuWriteback_23_bits_debug_isPerfCnt = io_exuWriteback_23_bits_debug_isPerfCnt;
        //    mon_tr.io_exuWriteback_23_bits_debug_paddr = io_exuWriteback_23_bits_debug_paddr;
        //    mon_tr.io_exuWriteback_22_valid = io_exuWriteback_22_valid;
        //    mon_tr.io_exuWriteback_22_bits_data_0 = io_exuWriteback_22_bits_data_0;
        //    mon_tr.io_exuWriteback_22_bits_robIdx_value = io_exuWriteback_22_bits_robIdx_value;
        //    mon_tr.io_exuWriteback_22_bits_lqIdx_value = io_exuWriteback_22_bits_lqIdx_value;
        //    mon_tr.io_exuWriteback_22_bits_debug_isMMIO = io_exuWriteback_22_bits_debug_isMMIO;
        //    mon_tr.io_exuWriteback_22_bits_debug_isNCIO = io_exuWriteback_22_bits_debug_isNCIO;
        //    mon_tr.io_exuWriteback_22_bits_debug_isPerfCnt = io_exuWriteback_22_bits_debug_isPerfCnt;
        //    mon_tr.io_exuWriteback_22_bits_debug_paddr = io_exuWriteback_22_bits_debug_paddr;
        //    mon_tr.io_exuWriteback_21_valid = io_exuWriteback_21_valid;
        //    mon_tr.io_exuWriteback_21_bits_data_0 = io_exuWriteback_21_bits_data_0;
        //    mon_tr.io_exuWriteback_21_bits_robIdx_value = io_exuWriteback_21_bits_robIdx_value;
        //    mon_tr.io_exuWriteback_21_bits_lqIdx_value = io_exuWriteback_21_bits_lqIdx_value;
        //    mon_tr.io_exuWriteback_21_bits_debug_isMMIO = io_exuWriteback_21_bits_debug_isMMIO;
        //    mon_tr.io_exuWriteback_21_bits_debug_isNCIO = io_exuWriteback_21_bits_debug_isNCIO;
        //    mon_tr.io_exuWriteback_21_bits_debug_isPerfCnt = io_exuWriteback_21_bits_debug_isPerfCnt;
        //    mon_tr.io_exuWriteback_21_bits_debug_paddr = io_exuWriteback_21_bits_debug_paddr;
        //    mon_tr.io_exuWriteback_20_valid = io_exuWriteback_20_valid;
        //    mon_tr.io_exuWriteback_20_bits_data_0 = io_exuWriteback_20_bits_data_0;
        //    mon_tr.io_exuWriteback_20_bits_robIdx_value = io_exuWriteback_20_bits_robIdx_value;
        //    mon_tr.io_exuWriteback_20_bits_lqIdx_value = io_exuWriteback_20_bits_lqIdx_value;
        //    mon_tr.io_exuWriteback_20_bits_debug_isMMIO = io_exuWriteback_20_bits_debug_isMMIO;
        //    mon_tr.io_exuWriteback_20_bits_debug_isNCIO = io_exuWriteback_20_bits_debug_isNCIO;
        //    mon_tr.io_exuWriteback_20_bits_debug_isPerfCnt = io_exuWriteback_20_bits_debug_isPerfCnt;
        //    mon_tr.io_exuWriteback_20_bits_debug_paddr = io_exuWriteback_20_bits_debug_paddr;
        //    mon_tr.io_exuWriteback_19_valid = io_exuWriteback_19_valid;
        //    mon_tr.io_exuWriteback_19_bits_data_0 = io_exuWriteback_19_bits_data_0;
        //    mon_tr.io_exuWriteback_19_bits_robIdx_value = io_exuWriteback_19_bits_robIdx_value;
        //    mon_tr.io_exuWriteback_19_bits_sqIdx_value = io_exuWriteback_19_bits_sqIdx_value;
        //    mon_tr.io_exuWriteback_19_bits_debug_isMMIO = io_exuWriteback_19_bits_debug_isMMIO;
        //    mon_tr.io_exuWriteback_19_bits_debug_isNCIO = io_exuWriteback_19_bits_debug_isNCIO;
        //    mon_tr.io_exuWriteback_19_bits_debug_isPerfCnt = io_exuWriteback_19_bits_debug_isPerfCnt;
        //    mon_tr.io_exuWriteback_19_bits_debug_paddr = io_exuWriteback_19_bits_debug_paddr;
        //    mon_tr.io_exuWriteback_18_valid = io_exuWriteback_18_valid;
        //    mon_tr.io_exuWriteback_18_bits_data_0 = io_exuWriteback_18_bits_data_0;
        //    mon_tr.io_exuWriteback_18_bits_robIdx_value = io_exuWriteback_18_bits_robIdx_value;
        //    mon_tr.io_exuWriteback_18_bits_sqIdx_value = io_exuWriteback_18_bits_sqIdx_value;
        //    mon_tr.io_exuWriteback_18_bits_debug_isMMIO = io_exuWriteback_18_bits_debug_isMMIO;
        //    mon_tr.io_exuWriteback_18_bits_debug_isNCIO = io_exuWriteback_18_bits_debug_isNCIO;
        //    mon_tr.io_exuWriteback_18_bits_debug_isPerfCnt = io_exuWriteback_18_bits_debug_isPerfCnt;
        //    mon_tr.io_exuWriteback_18_bits_debug_paddr = io_exuWriteback_18_bits_debug_paddr;
        //    mon_tr.io_exuWriteback_17_valid = io_exuWriteback_17_valid;
        //    mon_tr.io_exuWriteback_17_bits_data_0 = io_exuWriteback_17_bits_data_0;
        //    mon_tr.io_exuWriteback_17_bits_robIdx_value = io_exuWriteback_17_bits_robIdx_value;
        //    mon_tr.io_exuWriteback_17_bits_fflags = io_exuWriteback_17_bits_fflags;
        //    mon_tr.io_exuWriteback_17_bits_wflags = io_exuWriteback_17_bits_wflags;
        //    mon_tr.io_exuWriteback_16_valid = io_exuWriteback_16_valid;
        //    mon_tr.io_exuWriteback_16_bits_data_0 = io_exuWriteback_16_bits_data_0;
        //    mon_tr.io_exuWriteback_16_bits_robIdx_value = io_exuWriteback_16_bits_robIdx_value;
        //    mon_tr.io_exuWriteback_16_bits_fflags = io_exuWriteback_16_bits_fflags;
        //    mon_tr.io_exuWriteback_16_bits_wflags = io_exuWriteback_16_bits_wflags;
        //    mon_tr.io_exuWriteback_15_valid = io_exuWriteback_15_valid;
        //    mon_tr.io_exuWriteback_15_bits_data_0 = io_exuWriteback_15_bits_data_0;
        //    mon_tr.io_exuWriteback_15_bits_robIdx_value = io_exuWriteback_15_bits_robIdx_value;
        //    mon_tr.io_exuWriteback_15_bits_fflags = io_exuWriteback_15_bits_fflags;
        //    mon_tr.io_exuWriteback_15_bits_wflags = io_exuWriteback_15_bits_wflags;
        //    mon_tr.io_exuWriteback_15_bits_vxsat = io_exuWriteback_15_bits_vxsat;
        //    mon_tr.io_exuWriteback_14_valid = io_exuWriteback_14_valid;
        //    mon_tr.io_exuWriteback_14_bits_data_0 = io_exuWriteback_14_bits_data_0;
        //    mon_tr.io_exuWriteback_14_bits_robIdx_value = io_exuWriteback_14_bits_robIdx_value;
        //    mon_tr.io_exuWriteback_14_bits_fflags = io_exuWriteback_14_bits_fflags;
        //    mon_tr.io_exuWriteback_14_bits_wflags = io_exuWriteback_14_bits_wflags;
        //    mon_tr.io_exuWriteback_13_valid = io_exuWriteback_13_valid;
        //    mon_tr.io_exuWriteback_13_bits_data_0 = io_exuWriteback_13_bits_data_0;
        //    mon_tr.io_exuWriteback_13_bits_robIdx_value = io_exuWriteback_13_bits_robIdx_value;
        //    mon_tr.io_exuWriteback_13_bits_fflags = io_exuWriteback_13_bits_fflags;
        //    mon_tr.io_exuWriteback_13_bits_wflags = io_exuWriteback_13_bits_wflags;
        //    mon_tr.io_exuWriteback_13_bits_vxsat = io_exuWriteback_13_bits_vxsat;
        //    mon_tr.io_exuWriteback_12_valid = io_exuWriteback_12_valid;
        //    mon_tr.io_exuWriteback_12_bits_data_0 = io_exuWriteback_12_bits_data_0;
        //    mon_tr.io_exuWriteback_12_bits_robIdx_value = io_exuWriteback_12_bits_robIdx_value;
        //    mon_tr.io_exuWriteback_12_bits_fflags = io_exuWriteback_12_bits_fflags;
        //    mon_tr.io_exuWriteback_12_bits_wflags = io_exuWriteback_12_bits_wflags;
        //    mon_tr.io_exuWriteback_11_valid = io_exuWriteback_11_valid;
        //    mon_tr.io_exuWriteback_11_bits_data_0 = io_exuWriteback_11_bits_data_0;
        //    mon_tr.io_exuWriteback_11_bits_robIdx_value = io_exuWriteback_11_bits_robIdx_value;
        //    mon_tr.io_exuWriteback_11_bits_fflags = io_exuWriteback_11_bits_fflags;
        //    mon_tr.io_exuWriteback_11_bits_wflags = io_exuWriteback_11_bits_wflags;
        //    mon_tr.io_exuWriteback_10_valid = io_exuWriteback_10_valid;
        //    mon_tr.io_exuWriteback_10_bits_data_0 = io_exuWriteback_10_bits_data_0;
        //    mon_tr.io_exuWriteback_10_bits_robIdx_value = io_exuWriteback_10_bits_robIdx_value;
        //    mon_tr.io_exuWriteback_10_bits_fflags = io_exuWriteback_10_bits_fflags;
        //    mon_tr.io_exuWriteback_10_bits_wflags = io_exuWriteback_10_bits_wflags;
        //    mon_tr.io_exuWriteback_9_valid = io_exuWriteback_9_valid;
        //    mon_tr.io_exuWriteback_9_bits_data_0 = io_exuWriteback_9_bits_data_0;
        //    mon_tr.io_exuWriteback_9_bits_robIdx_value = io_exuWriteback_9_bits_robIdx_value;
        //    mon_tr.io_exuWriteback_9_bits_fflags = io_exuWriteback_9_bits_fflags;
        //    mon_tr.io_exuWriteback_9_bits_wflags = io_exuWriteback_9_bits_wflags;
        //    mon_tr.io_exuWriteback_8_valid = io_exuWriteback_8_valid;
        //    mon_tr.io_exuWriteback_8_bits_data_0 = io_exuWriteback_8_bits_data_0;
        //    mon_tr.io_exuWriteback_8_bits_robIdx_value = io_exuWriteback_8_bits_robIdx_value;
        //    mon_tr.io_exuWriteback_8_bits_fflags = io_exuWriteback_8_bits_fflags;
        //    mon_tr.io_exuWriteback_8_bits_wflags = io_exuWriteback_8_bits_wflags;
        //    mon_tr.io_exuWriteback_7_valid = io_exuWriteback_7_valid;
        //    mon_tr.io_exuWriteback_7_bits_data_0 = io_exuWriteback_7_bits_data_0;
        //    mon_tr.io_exuWriteback_7_bits_robIdx_value = io_exuWriteback_7_bits_robIdx_value;
        //    mon_tr.io_exuWriteback_7_bits_debug_isPerfCnt = io_exuWriteback_7_bits_debug_isPerfCnt;
        //    mon_tr.io_exuWriteback_6_valid = io_exuWriteback_6_valid;
        //    mon_tr.io_exuWriteback_6_bits_data_0 = io_exuWriteback_6_bits_data_0;
        //    mon_tr.io_exuWriteback_6_bits_robIdx_value = io_exuWriteback_6_bits_robIdx_value;
        //    mon_tr.io_exuWriteback_5_valid = io_exuWriteback_5_valid;
        //    mon_tr.io_exuWriteback_5_bits_data_0 = io_exuWriteback_5_bits_data_0;
        //    mon_tr.io_exuWriteback_5_bits_robIdx_value = io_exuWriteback_5_bits_robIdx_value;
        //    mon_tr.io_exuWriteback_5_bits_redirect_valid = io_exuWriteback_5_bits_redirect_valid;
        //    mon_tr.io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken = io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken;
        //    mon_tr.io_exuWriteback_5_bits_fflags = io_exuWriteback_5_bits_fflags;
        //    mon_tr.io_exuWriteback_5_bits_wflags = io_exuWriteback_5_bits_wflags;
        //    mon_tr.io_exuWriteback_4_valid = io_exuWriteback_4_valid;
        //    mon_tr.io_exuWriteback_4_bits_data_0 = io_exuWriteback_4_bits_data_0;
        //    mon_tr.io_exuWriteback_4_bits_robIdx_value = io_exuWriteback_4_bits_robIdx_value;
        //    mon_tr.io_exuWriteback_3_valid = io_exuWriteback_3_valid;
        //    mon_tr.io_exuWriteback_3_bits_data_0 = io_exuWriteback_3_bits_data_0;
        //    mon_tr.io_exuWriteback_3_bits_robIdx_value = io_exuWriteback_3_bits_robIdx_value;
        //    mon_tr.io_exuWriteback_3_bits_redirect_valid = io_exuWriteback_3_bits_redirect_valid;
        //    mon_tr.io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken = io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken;
        //    mon_tr.io_exuWriteback_2_valid = io_exuWriteback_2_valid;
        //    mon_tr.io_exuWriteback_2_bits_data_0 = io_exuWriteback_2_bits_data_0;
        //    mon_tr.io_exuWriteback_2_bits_robIdx_value = io_exuWriteback_2_bits_robIdx_value;
        //    mon_tr.io_exuWriteback_1_valid = io_exuWriteback_1_valid;
        //    mon_tr.io_exuWriteback_1_bits_data_0 = io_exuWriteback_1_bits_data_0;
        //    mon_tr.io_exuWriteback_1_bits_robIdx_value = io_exuWriteback_1_bits_robIdx_value;
        //    mon_tr.io_exuWriteback_1_bits_redirect_valid = io_exuWriteback_1_bits_redirect_valid;
        //    mon_tr.io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken = io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken;
        //    mon_tr.io_exuWriteback_0_valid = io_exuWriteback_0_valid;
        //    mon_tr.io_exuWriteback_0_bits_data_0 = io_exuWriteback_0_bits_data_0;
        //    mon_tr.io_exuWriteback_0_bits_robIdx_value = io_exuWriteback_0_bits_robIdx_value;
        //    mon_tr.io_writebackNums_0_bits = io_writebackNums_0_bits;
        //    mon_tr.io_writebackNums_1_bits = io_writebackNums_1_bits;
        //    mon_tr.io_writebackNums_2_bits = io_writebackNums_2_bits;
        //    mon_tr.io_writebackNums_3_bits = io_writebackNums_3_bits;
        //    mon_tr.io_writebackNums_4_bits = io_writebackNums_4_bits;
        //    mon_tr.io_writebackNums_5_bits = io_writebackNums_5_bits;
        //    mon_tr.io_writebackNums_6_bits = io_writebackNums_6_bits;
        //    mon_tr.io_writebackNums_7_bits = io_writebackNums_7_bits;
        //    mon_tr.io_writebackNums_8_bits = io_writebackNums_8_bits;
        //    mon_tr.io_writebackNums_9_bits = io_writebackNums_9_bits;
        //    mon_tr.io_writebackNums_10_bits = io_writebackNums_10_bits;
        //    mon_tr.io_writebackNums_11_bits = io_writebackNums_11_bits;
        //    mon_tr.io_writebackNums_12_bits = io_writebackNums_12_bits;
        //    mon_tr.io_writebackNums_13_bits = io_writebackNums_13_bits;
        //    mon_tr.io_writebackNums_14_bits = io_writebackNums_14_bits;
        //    mon_tr.io_writebackNums_15_bits = io_writebackNums_15_bits;
        //    mon_tr.io_writebackNums_16_bits = io_writebackNums_16_bits;
        //    mon_tr.io_writebackNums_17_bits = io_writebackNums_17_bits;
        //    mon_tr.io_writebackNums_18_bits = io_writebackNums_18_bits;
        //    mon_tr.io_writebackNums_19_bits = io_writebackNums_19_bits;
        //    mon_tr.io_writebackNums_20_bits = io_writebackNums_20_bits;
        //    mon_tr.io_writebackNums_21_bits = io_writebackNums_21_bits;
        //    mon_tr.io_writebackNums_22_bits = io_writebackNums_22_bits;
        //    mon_tr.io_writebackNums_23_bits = io_writebackNums_23_bits;
        //    mon_tr.io_writebackNums_24_bits = io_writebackNums_24_bits;
        //    mon_tr.io_writebackNeedFlush_0 = io_writebackNeedFlush_0;
        //    mon_tr.io_writebackNeedFlush_1 = io_writebackNeedFlush_1;
        //    mon_tr.io_writebackNeedFlush_2 = io_writebackNeedFlush_2;
        //    mon_tr.io_writebackNeedFlush_6 = io_writebackNeedFlush_6;
        //    mon_tr.io_writebackNeedFlush_7 = io_writebackNeedFlush_7;
        //    mon_tr.io_writebackNeedFlush_8 = io_writebackNeedFlush_8;
        //    mon_tr.io_writebackNeedFlush_9 = io_writebackNeedFlush_9;
        //    mon_tr.io_writebackNeedFlush_10 = io_writebackNeedFlush_10;
        //    mon_tr.io_writebackNeedFlush_11 = io_writebackNeedFlush_11;
        //    mon_tr.io_writebackNeedFlush_12 = io_writebackNeedFlush_12;

        //    mon_tr.channel_id = this.cfg.channel_id;
        //    mon_tr.unpack();
        //    this.mon_item_port.write(mon_tr);
        //end
    end
endtask:mon_data

`endif


//=========================================================
//File name    : WriteBack_in_agent_dec.sv
//Author       : nanyunhao
//Module name  : WriteBack_in_agent_dec
//Discribution : WriteBack_in_agent_dec : parameter
//Date         : 2026-01-22
//=========================================================
`ifndef WRITEBACK_IN_AGENT_DEC__SV
`define WRITEBACK_IN_AGENT_DEC__SV

package WriteBack_in_agent_dec;

endpackage:WriteBack_in_agent_dec

import WriteBack_in_agent_dec::*;

`endif


//=========================================================
//File name    : Rob_output_connect.sv
//Author       : nanyunhao
//Module name  : Rob_output_connect
//Discribution : Rob_output_connect : Rob_output Interface connection macro
//Date         : 2026-01-22
//=========================================================
`ifndef ROB_OUTPUT_CONNECT__SV
`define ROB_OUTPUT_CONNECT__SV

`define ROB__ROB_OUTPUT_CONNECT(U_IF_NAME,AGENT_PATH,RTL_PATH) \
    Rob_output_agent_interface  U_IF_NAME (clk,tc_if.rst_n); \
    initial begin \
        uvm_config_db#(virtual Rob_output_agent_interface)::set(null,`"*AGENT_PATH*`", "vif", U_IF_NAME); \
    end \
    `ifdef ROB_UT \
    initial begin \
        force U_IF_NAME.io_enq_canAccept = RTL_PATH.io_enq_canAccept; \
        force U_IF_NAME.io_enq_canAcceptForDispatch = RTL_PATH.io_enq_canAcceptForDispatch; \
        force U_IF_NAME.io_enq_isEmpty = RTL_PATH.io_enq_isEmpty; \
        force U_IF_NAME.io_flushOut_valid = RTL_PATH.io_flushOut_valid; \
        force U_IF_NAME.io_flushOut_bits_isRVC = RTL_PATH.io_flushOut_bits_isRVC; \
        force U_IF_NAME.io_flushOut_bits_robIdx_flag = RTL_PATH.io_flushOut_bits_robIdx_flag; \
        force U_IF_NAME.io_flushOut_bits_robIdx_value = RTL_PATH.io_flushOut_bits_robIdx_value; \
        force U_IF_NAME.io_flushOut_bits_ftqIdx_flag = RTL_PATH.io_flushOut_bits_ftqIdx_flag; \
        force U_IF_NAME.io_flushOut_bits_ftqIdx_value = RTL_PATH.io_flushOut_bits_ftqIdx_value; \
        force U_IF_NAME.io_flushOut_bits_ftqOffset = RTL_PATH.io_flushOut_bits_ftqOffset; \
        force U_IF_NAME.io_flushOut_bits_level = RTL_PATH.io_flushOut_bits_level; \
        force U_IF_NAME.io_exception_valid = RTL_PATH.io_exception_valid; \
        force U_IF_NAME.io_exception_bits_instr = RTL_PATH.io_exception_bits_instr; \
        force U_IF_NAME.io_exception_bits_commitType = RTL_PATH.io_exception_bits_commitType; \
        force U_IF_NAME.io_exception_bits_exceptionVec_0 = RTL_PATH.io_exception_bits_exceptionVec_0; \
        force U_IF_NAME.io_exception_bits_exceptionVec_1 = RTL_PATH.io_exception_bits_exceptionVec_1; \
        force U_IF_NAME.io_exception_bits_exceptionVec_2 = RTL_PATH.io_exception_bits_exceptionVec_2; \
        force U_IF_NAME.io_exception_bits_exceptionVec_3 = RTL_PATH.io_exception_bits_exceptionVec_3; \
        force U_IF_NAME.io_exception_bits_exceptionVec_4 = RTL_PATH.io_exception_bits_exceptionVec_4; \
        force U_IF_NAME.io_exception_bits_exceptionVec_5 = RTL_PATH.io_exception_bits_exceptionVec_5; \
        force U_IF_NAME.io_exception_bits_exceptionVec_6 = RTL_PATH.io_exception_bits_exceptionVec_6; \
        force U_IF_NAME.io_exception_bits_exceptionVec_7 = RTL_PATH.io_exception_bits_exceptionVec_7; \
        force U_IF_NAME.io_exception_bits_exceptionVec_8 = RTL_PATH.io_exception_bits_exceptionVec_8; \
        force U_IF_NAME.io_exception_bits_exceptionVec_9 = RTL_PATH.io_exception_bits_exceptionVec_9; \
        force U_IF_NAME.io_exception_bits_exceptionVec_10 = RTL_PATH.io_exception_bits_exceptionVec_10; \
        force U_IF_NAME.io_exception_bits_exceptionVec_11 = RTL_PATH.io_exception_bits_exceptionVec_11; \
        force U_IF_NAME.io_exception_bits_exceptionVec_12 = RTL_PATH.io_exception_bits_exceptionVec_12; \
        force U_IF_NAME.io_exception_bits_exceptionVec_13 = RTL_PATH.io_exception_bits_exceptionVec_13; \
        force U_IF_NAME.io_exception_bits_exceptionVec_14 = RTL_PATH.io_exception_bits_exceptionVec_14; \
        force U_IF_NAME.io_exception_bits_exceptionVec_15 = RTL_PATH.io_exception_bits_exceptionVec_15; \
        force U_IF_NAME.io_exception_bits_exceptionVec_16 = RTL_PATH.io_exception_bits_exceptionVec_16; \
        force U_IF_NAME.io_exception_bits_exceptionVec_17 = RTL_PATH.io_exception_bits_exceptionVec_17; \
        force U_IF_NAME.io_exception_bits_exceptionVec_18 = RTL_PATH.io_exception_bits_exceptionVec_18; \
        force U_IF_NAME.io_exception_bits_exceptionVec_19 = RTL_PATH.io_exception_bits_exceptionVec_19; \
        force U_IF_NAME.io_exception_bits_exceptionVec_20 = RTL_PATH.io_exception_bits_exceptionVec_20; \
        force U_IF_NAME.io_exception_bits_exceptionVec_21 = RTL_PATH.io_exception_bits_exceptionVec_21; \
        force U_IF_NAME.io_exception_bits_exceptionVec_22 = RTL_PATH.io_exception_bits_exceptionVec_22; \
        force U_IF_NAME.io_exception_bits_exceptionVec_23 = RTL_PATH.io_exception_bits_exceptionVec_23; \
        force U_IF_NAME.io_exception_bits_isPcBkpt = RTL_PATH.io_exception_bits_isPcBkpt; \
        force U_IF_NAME.io_exception_bits_isFetchMalAddr = RTL_PATH.io_exception_bits_isFetchMalAddr; \
        force U_IF_NAME.io_exception_bits_gpaddr = RTL_PATH.io_exception_bits_gpaddr; \
        force U_IF_NAME.io_exception_bits_singleStep = RTL_PATH.io_exception_bits_singleStep; \
        force U_IF_NAME.io_exception_bits_crossPageIPFFix = RTL_PATH.io_exception_bits_crossPageIPFFix; \
        force U_IF_NAME.io_exception_bits_isInterrupt = RTL_PATH.io_exception_bits_isInterrupt; \
        force U_IF_NAME.io_exception_bits_isHls = RTL_PATH.io_exception_bits_isHls; \
        force U_IF_NAME.io_exception_bits_trigger = RTL_PATH.io_exception_bits_trigger; \
        force U_IF_NAME.io_exception_bits_isForVSnonLeafPTE = RTL_PATH.io_exception_bits_isForVSnonLeafPTE; \
        force U_IF_NAME.io_commits_isCommit = RTL_PATH.io_commits_isCommit; \
        force U_IF_NAME.io_commits_commitValid_0 = RTL_PATH.io_commits_commitValid_0; \
        force U_IF_NAME.io_commits_commitValid_1 = RTL_PATH.io_commits_commitValid_1; \
        force U_IF_NAME.io_commits_commitValid_2 = RTL_PATH.io_commits_commitValid_2; \
        force U_IF_NAME.io_commits_commitValid_3 = RTL_PATH.io_commits_commitValid_3; \
        force U_IF_NAME.io_commits_commitValid_4 = RTL_PATH.io_commits_commitValid_4; \
        force U_IF_NAME.io_commits_commitValid_5 = RTL_PATH.io_commits_commitValid_5; \
        force U_IF_NAME.io_commits_commitValid_6 = RTL_PATH.io_commits_commitValid_6; \
        force U_IF_NAME.io_commits_commitValid_7 = RTL_PATH.io_commits_commitValid_7; \
        force U_IF_NAME.io_commits_isWalk = RTL_PATH.io_commits_isWalk; \
        force U_IF_NAME.io_commits_walkValid_0 = RTL_PATH.io_commits_walkValid_0; \
        force U_IF_NAME.io_commits_walkValid_1 = RTL_PATH.io_commits_walkValid_1; \
        force U_IF_NAME.io_commits_walkValid_2 = RTL_PATH.io_commits_walkValid_2; \
        force U_IF_NAME.io_commits_walkValid_3 = RTL_PATH.io_commits_walkValid_3; \
        force U_IF_NAME.io_commits_walkValid_4 = RTL_PATH.io_commits_walkValid_4; \
        force U_IF_NAME.io_commits_walkValid_5 = RTL_PATH.io_commits_walkValid_5; \
        force U_IF_NAME.io_commits_walkValid_6 = RTL_PATH.io_commits_walkValid_6; \
        force U_IF_NAME.io_commits_walkValid_7 = RTL_PATH.io_commits_walkValid_7; \
        force U_IF_NAME.io_commits_info_0_walk_v = RTL_PATH.io_commits_info_0_walk_v; \
        force U_IF_NAME.io_commits_info_0_commit_v = RTL_PATH.io_commits_info_0_commit_v; \
        force U_IF_NAME.io_commits_info_0_commit_w = RTL_PATH.io_commits_info_0_commit_w; \
        force U_IF_NAME.io_commits_info_0_realDestSize = RTL_PATH.io_commits_info_0_realDestSize; \
        force U_IF_NAME.io_commits_info_0_interrupt_safe = RTL_PATH.io_commits_info_0_interrupt_safe; \
        force U_IF_NAME.io_commits_info_0_wflags = RTL_PATH.io_commits_info_0_wflags; \
        force U_IF_NAME.io_commits_info_0_fflags = RTL_PATH.io_commits_info_0_fflags; \
        force U_IF_NAME.io_commits_info_0_vxsat = RTL_PATH.io_commits_info_0_vxsat; \
        force U_IF_NAME.io_commits_info_0_isRVC = RTL_PATH.io_commits_info_0_isRVC; \
        force U_IF_NAME.io_commits_info_0_isVset = RTL_PATH.io_commits_info_0_isVset; \
        force U_IF_NAME.io_commits_info_0_isHls = RTL_PATH.io_commits_info_0_isHls; \
        force U_IF_NAME.io_commits_info_0_isVls = RTL_PATH.io_commits_info_0_isVls; \
        force U_IF_NAME.io_commits_info_0_vls = RTL_PATH.io_commits_info_0_vls; \
        force U_IF_NAME.io_commits_info_0_mmio = RTL_PATH.io_commits_info_0_mmio; \
        force U_IF_NAME.io_commits_info_0_commitType = RTL_PATH.io_commits_info_0_commitType; \
        force U_IF_NAME.io_commits_info_0_ftqIdx_flag = RTL_PATH.io_commits_info_0_ftqIdx_flag; \
        force U_IF_NAME.io_commits_info_0_ftqIdx_value = RTL_PATH.io_commits_info_0_ftqIdx_value; \
        force U_IF_NAME.io_commits_info_0_ftqOffset = RTL_PATH.io_commits_info_0_ftqOffset; \
        force U_IF_NAME.io_commits_info_0_instrSize = RTL_PATH.io_commits_info_0_instrSize; \
        force U_IF_NAME.io_commits_info_0_fpWen = RTL_PATH.io_commits_info_0_fpWen; \
        force U_IF_NAME.io_commits_info_0_rfWen = RTL_PATH.io_commits_info_0_rfWen; \
        force U_IF_NAME.io_commits_info_0_needFlush = RTL_PATH.io_commits_info_0_needFlush; \
        force U_IF_NAME.io_commits_info_0_traceBlockInPipe_itype = RTL_PATH.io_commits_info_0_traceBlockInPipe_itype; \
        force U_IF_NAME.io_commits_info_0_traceBlockInPipe_iretire = RTL_PATH.io_commits_info_0_traceBlockInPipe_iretire; \
        force U_IF_NAME.io_commits_info_0_traceBlockInPipe_ilastsize = RTL_PATH.io_commits_info_0_traceBlockInPipe_ilastsize; \
        force U_IF_NAME.io_commits_info_0_debug_pc = RTL_PATH.io_commits_info_0_debug_pc; \
        force U_IF_NAME.io_commits_info_0_debug_instr = RTL_PATH.io_commits_info_0_debug_instr; \
        force U_IF_NAME.io_commits_info_0_debug_ldest = RTL_PATH.io_commits_info_0_debug_ldest; \
        force U_IF_NAME.io_commits_info_0_debug_pdest = RTL_PATH.io_commits_info_0_debug_pdest; \
        force U_IF_NAME.io_commits_info_0_debug_otherPdest_0 = RTL_PATH.io_commits_info_0_debug_otherPdest_0; \
        force U_IF_NAME.io_commits_info_0_debug_otherPdest_1 = RTL_PATH.io_commits_info_0_debug_otherPdest_1; \
        force U_IF_NAME.io_commits_info_0_debug_otherPdest_2 = RTL_PATH.io_commits_info_0_debug_otherPdest_2; \
        force U_IF_NAME.io_commits_info_0_debug_otherPdest_3 = RTL_PATH.io_commits_info_0_debug_otherPdest_3; \
        force U_IF_NAME.io_commits_info_0_debug_otherPdest_4 = RTL_PATH.io_commits_info_0_debug_otherPdest_4; \
        force U_IF_NAME.io_commits_info_0_debug_otherPdest_5 = RTL_PATH.io_commits_info_0_debug_otherPdest_5; \
        force U_IF_NAME.io_commits_info_0_debug_otherPdest_6 = RTL_PATH.io_commits_info_0_debug_otherPdest_6; \
        force U_IF_NAME.io_commits_info_0_debug_fuType = RTL_PATH.io_commits_info_0_debug_fuType; \
        force U_IF_NAME.io_commits_info_0_dirtyFs = RTL_PATH.io_commits_info_0_dirtyFs; \
        force U_IF_NAME.io_commits_info_0_dirtyVs = RTL_PATH.io_commits_info_0_dirtyVs; \
        force U_IF_NAME.io_commits_info_1_walk_v = RTL_PATH.io_commits_info_1_walk_v; \
        force U_IF_NAME.io_commits_info_1_commit_v = RTL_PATH.io_commits_info_1_commit_v; \
        force U_IF_NAME.io_commits_info_1_commit_w = RTL_PATH.io_commits_info_1_commit_w; \
        force U_IF_NAME.io_commits_info_1_realDestSize = RTL_PATH.io_commits_info_1_realDestSize; \
        force U_IF_NAME.io_commits_info_1_interrupt_safe = RTL_PATH.io_commits_info_1_interrupt_safe; \
        force U_IF_NAME.io_commits_info_1_wflags = RTL_PATH.io_commits_info_1_wflags; \
        force U_IF_NAME.io_commits_info_1_fflags = RTL_PATH.io_commits_info_1_fflags; \
        force U_IF_NAME.io_commits_info_1_vxsat = RTL_PATH.io_commits_info_1_vxsat; \
        force U_IF_NAME.io_commits_info_1_isRVC = RTL_PATH.io_commits_info_1_isRVC; \
        force U_IF_NAME.io_commits_info_1_isVset = RTL_PATH.io_commits_info_1_isVset; \
        force U_IF_NAME.io_commits_info_1_isHls = RTL_PATH.io_commits_info_1_isHls; \
        force U_IF_NAME.io_commits_info_1_isVls = RTL_PATH.io_commits_info_1_isVls; \
        force U_IF_NAME.io_commits_info_1_vls = RTL_PATH.io_commits_info_1_vls; \
        force U_IF_NAME.io_commits_info_1_mmio = RTL_PATH.io_commits_info_1_mmio; \
        force U_IF_NAME.io_commits_info_1_commitType = RTL_PATH.io_commits_info_1_commitType; \
        force U_IF_NAME.io_commits_info_1_ftqIdx_flag = RTL_PATH.io_commits_info_1_ftqIdx_flag; \
        force U_IF_NAME.io_commits_info_1_ftqIdx_value = RTL_PATH.io_commits_info_1_ftqIdx_value; \
        force U_IF_NAME.io_commits_info_1_ftqOffset = RTL_PATH.io_commits_info_1_ftqOffset; \
        force U_IF_NAME.io_commits_info_1_instrSize = RTL_PATH.io_commits_info_1_instrSize; \
        force U_IF_NAME.io_commits_info_1_fpWen = RTL_PATH.io_commits_info_1_fpWen; \
        force U_IF_NAME.io_commits_info_1_rfWen = RTL_PATH.io_commits_info_1_rfWen; \
        force U_IF_NAME.io_commits_info_1_needFlush = RTL_PATH.io_commits_info_1_needFlush; \
        force U_IF_NAME.io_commits_info_1_traceBlockInPipe_itype = RTL_PATH.io_commits_info_1_traceBlockInPipe_itype; \
        force U_IF_NAME.io_commits_info_1_traceBlockInPipe_iretire = RTL_PATH.io_commits_info_1_traceBlockInPipe_iretire; \
        force U_IF_NAME.io_commits_info_1_traceBlockInPipe_ilastsize = RTL_PATH.io_commits_info_1_traceBlockInPipe_ilastsize; \
        force U_IF_NAME.io_commits_info_1_debug_pc = RTL_PATH.io_commits_info_1_debug_pc; \
        force U_IF_NAME.io_commits_info_1_debug_instr = RTL_PATH.io_commits_info_1_debug_instr; \
        force U_IF_NAME.io_commits_info_1_debug_ldest = RTL_PATH.io_commits_info_1_debug_ldest; \
        force U_IF_NAME.io_commits_info_1_debug_pdest = RTL_PATH.io_commits_info_1_debug_pdest; \
        force U_IF_NAME.io_commits_info_1_debug_otherPdest_0 = RTL_PATH.io_commits_info_1_debug_otherPdest_0; \
        force U_IF_NAME.io_commits_info_1_debug_otherPdest_1 = RTL_PATH.io_commits_info_1_debug_otherPdest_1; \
        force U_IF_NAME.io_commits_info_1_debug_otherPdest_2 = RTL_PATH.io_commits_info_1_debug_otherPdest_2; \
        force U_IF_NAME.io_commits_info_1_debug_otherPdest_3 = RTL_PATH.io_commits_info_1_debug_otherPdest_3; \
        force U_IF_NAME.io_commits_info_1_debug_otherPdest_4 = RTL_PATH.io_commits_info_1_debug_otherPdest_4; \
        force U_IF_NAME.io_commits_info_1_debug_otherPdest_5 = RTL_PATH.io_commits_info_1_debug_otherPdest_5; \
        force U_IF_NAME.io_commits_info_1_debug_otherPdest_6 = RTL_PATH.io_commits_info_1_debug_otherPdest_6; \
        force U_IF_NAME.io_commits_info_1_debug_fuType = RTL_PATH.io_commits_info_1_debug_fuType; \
        force U_IF_NAME.io_commits_info_1_dirtyFs = RTL_PATH.io_commits_info_1_dirtyFs; \
        force U_IF_NAME.io_commits_info_1_dirtyVs = RTL_PATH.io_commits_info_1_dirtyVs; \
        force U_IF_NAME.io_commits_info_2_walk_v = RTL_PATH.io_commits_info_2_walk_v; \
        force U_IF_NAME.io_commits_info_2_commit_v = RTL_PATH.io_commits_info_2_commit_v; \
        force U_IF_NAME.io_commits_info_2_commit_w = RTL_PATH.io_commits_info_2_commit_w; \
        force U_IF_NAME.io_commits_info_2_realDestSize = RTL_PATH.io_commits_info_2_realDestSize; \
        force U_IF_NAME.io_commits_info_2_interrupt_safe = RTL_PATH.io_commits_info_2_interrupt_safe; \
        force U_IF_NAME.io_commits_info_2_wflags = RTL_PATH.io_commits_info_2_wflags; \
        force U_IF_NAME.io_commits_info_2_fflags = RTL_PATH.io_commits_info_2_fflags; \
        force U_IF_NAME.io_commits_info_2_vxsat = RTL_PATH.io_commits_info_2_vxsat; \
        force U_IF_NAME.io_commits_info_2_isRVC = RTL_PATH.io_commits_info_2_isRVC; \
        force U_IF_NAME.io_commits_info_2_isVset = RTL_PATH.io_commits_info_2_isVset; \
        force U_IF_NAME.io_commits_info_2_isHls = RTL_PATH.io_commits_info_2_isHls; \
        force U_IF_NAME.io_commits_info_2_isVls = RTL_PATH.io_commits_info_2_isVls; \
        force U_IF_NAME.io_commits_info_2_vls = RTL_PATH.io_commits_info_2_vls; \
        force U_IF_NAME.io_commits_info_2_mmio = RTL_PATH.io_commits_info_2_mmio; \
        force U_IF_NAME.io_commits_info_2_commitType = RTL_PATH.io_commits_info_2_commitType; \
        force U_IF_NAME.io_commits_info_2_ftqIdx_flag = RTL_PATH.io_commits_info_2_ftqIdx_flag; \
        force U_IF_NAME.io_commits_info_2_ftqIdx_value = RTL_PATH.io_commits_info_2_ftqIdx_value; \
        force U_IF_NAME.io_commits_info_2_ftqOffset = RTL_PATH.io_commits_info_2_ftqOffset; \
        force U_IF_NAME.io_commits_info_2_instrSize = RTL_PATH.io_commits_info_2_instrSize; \
        force U_IF_NAME.io_commits_info_2_fpWen = RTL_PATH.io_commits_info_2_fpWen; \
        force U_IF_NAME.io_commits_info_2_rfWen = RTL_PATH.io_commits_info_2_rfWen; \
        force U_IF_NAME.io_commits_info_2_needFlush = RTL_PATH.io_commits_info_2_needFlush; \
        force U_IF_NAME.io_commits_info_2_traceBlockInPipe_itype = RTL_PATH.io_commits_info_2_traceBlockInPipe_itype; \
        force U_IF_NAME.io_commits_info_2_traceBlockInPipe_iretire = RTL_PATH.io_commits_info_2_traceBlockInPipe_iretire; \
        force U_IF_NAME.io_commits_info_2_traceBlockInPipe_ilastsize = RTL_PATH.io_commits_info_2_traceBlockInPipe_ilastsize; \
        force U_IF_NAME.io_commits_info_2_debug_pc = RTL_PATH.io_commits_info_2_debug_pc; \
        force U_IF_NAME.io_commits_info_2_debug_instr = RTL_PATH.io_commits_info_2_debug_instr; \
        force U_IF_NAME.io_commits_info_2_debug_ldest = RTL_PATH.io_commits_info_2_debug_ldest; \
        force U_IF_NAME.io_commits_info_2_debug_pdest = RTL_PATH.io_commits_info_2_debug_pdest; \
        force U_IF_NAME.io_commits_info_2_debug_otherPdest_0 = RTL_PATH.io_commits_info_2_debug_otherPdest_0; \
        force U_IF_NAME.io_commits_info_2_debug_otherPdest_1 = RTL_PATH.io_commits_info_2_debug_otherPdest_1; \
        force U_IF_NAME.io_commits_info_2_debug_otherPdest_2 = RTL_PATH.io_commits_info_2_debug_otherPdest_2; \
        force U_IF_NAME.io_commits_info_2_debug_otherPdest_3 = RTL_PATH.io_commits_info_2_debug_otherPdest_3; \
        force U_IF_NAME.io_commits_info_2_debug_otherPdest_4 = RTL_PATH.io_commits_info_2_debug_otherPdest_4; \
        force U_IF_NAME.io_commits_info_2_debug_otherPdest_5 = RTL_PATH.io_commits_info_2_debug_otherPdest_5; \
        force U_IF_NAME.io_commits_info_2_debug_otherPdest_6 = RTL_PATH.io_commits_info_2_debug_otherPdest_6; \
        force U_IF_NAME.io_commits_info_2_debug_fuType = RTL_PATH.io_commits_info_2_debug_fuType; \
        force U_IF_NAME.io_commits_info_2_dirtyFs = RTL_PATH.io_commits_info_2_dirtyFs; \
        force U_IF_NAME.io_commits_info_2_dirtyVs = RTL_PATH.io_commits_info_2_dirtyVs; \
        force U_IF_NAME.io_commits_info_3_walk_v = RTL_PATH.io_commits_info_3_walk_v; \
        force U_IF_NAME.io_commits_info_3_commit_v = RTL_PATH.io_commits_info_3_commit_v; \
        force U_IF_NAME.io_commits_info_3_commit_w = RTL_PATH.io_commits_info_3_commit_w; \
        force U_IF_NAME.io_commits_info_3_realDestSize = RTL_PATH.io_commits_info_3_realDestSize; \
        force U_IF_NAME.io_commits_info_3_interrupt_safe = RTL_PATH.io_commits_info_3_interrupt_safe; \
        force U_IF_NAME.io_commits_info_3_wflags = RTL_PATH.io_commits_info_3_wflags; \
        force U_IF_NAME.io_commits_info_3_fflags = RTL_PATH.io_commits_info_3_fflags; \
        force U_IF_NAME.io_commits_info_3_vxsat = RTL_PATH.io_commits_info_3_vxsat; \
        force U_IF_NAME.io_commits_info_3_isRVC = RTL_PATH.io_commits_info_3_isRVC; \
        force U_IF_NAME.io_commits_info_3_isVset = RTL_PATH.io_commits_info_3_isVset; \
        force U_IF_NAME.io_commits_info_3_isHls = RTL_PATH.io_commits_info_3_isHls; \
        force U_IF_NAME.io_commits_info_3_isVls = RTL_PATH.io_commits_info_3_isVls; \
        force U_IF_NAME.io_commits_info_3_vls = RTL_PATH.io_commits_info_3_vls; \
        force U_IF_NAME.io_commits_info_3_mmio = RTL_PATH.io_commits_info_3_mmio; \
        force U_IF_NAME.io_commits_info_3_commitType = RTL_PATH.io_commits_info_3_commitType; \
        force U_IF_NAME.io_commits_info_3_ftqIdx_flag = RTL_PATH.io_commits_info_3_ftqIdx_flag; \
        force U_IF_NAME.io_commits_info_3_ftqIdx_value = RTL_PATH.io_commits_info_3_ftqIdx_value; \
        force U_IF_NAME.io_commits_info_3_ftqOffset = RTL_PATH.io_commits_info_3_ftqOffset; \
        force U_IF_NAME.io_commits_info_3_instrSize = RTL_PATH.io_commits_info_3_instrSize; \
        force U_IF_NAME.io_commits_info_3_fpWen = RTL_PATH.io_commits_info_3_fpWen; \
        force U_IF_NAME.io_commits_info_3_rfWen = RTL_PATH.io_commits_info_3_rfWen; \
        force U_IF_NAME.io_commits_info_3_needFlush = RTL_PATH.io_commits_info_3_needFlush; \
        force U_IF_NAME.io_commits_info_3_traceBlockInPipe_itype = RTL_PATH.io_commits_info_3_traceBlockInPipe_itype; \
        force U_IF_NAME.io_commits_info_3_traceBlockInPipe_iretire = RTL_PATH.io_commits_info_3_traceBlockInPipe_iretire; \
        force U_IF_NAME.io_commits_info_3_traceBlockInPipe_ilastsize = RTL_PATH.io_commits_info_3_traceBlockInPipe_ilastsize; \
        force U_IF_NAME.io_commits_info_3_debug_pc = RTL_PATH.io_commits_info_3_debug_pc; \
        force U_IF_NAME.io_commits_info_3_debug_instr = RTL_PATH.io_commits_info_3_debug_instr; \
        force U_IF_NAME.io_commits_info_3_debug_ldest = RTL_PATH.io_commits_info_3_debug_ldest; \
        force U_IF_NAME.io_commits_info_3_debug_pdest = RTL_PATH.io_commits_info_3_debug_pdest; \
        force U_IF_NAME.io_commits_info_3_debug_otherPdest_0 = RTL_PATH.io_commits_info_3_debug_otherPdest_0; \
        force U_IF_NAME.io_commits_info_3_debug_otherPdest_1 = RTL_PATH.io_commits_info_3_debug_otherPdest_1; \
        force U_IF_NAME.io_commits_info_3_debug_otherPdest_2 = RTL_PATH.io_commits_info_3_debug_otherPdest_2; \
        force U_IF_NAME.io_commits_info_3_debug_otherPdest_3 = RTL_PATH.io_commits_info_3_debug_otherPdest_3; \
        force U_IF_NAME.io_commits_info_3_debug_otherPdest_4 = RTL_PATH.io_commits_info_3_debug_otherPdest_4; \
        force U_IF_NAME.io_commits_info_3_debug_otherPdest_5 = RTL_PATH.io_commits_info_3_debug_otherPdest_5; \
        force U_IF_NAME.io_commits_info_3_debug_otherPdest_6 = RTL_PATH.io_commits_info_3_debug_otherPdest_6; \
        force U_IF_NAME.io_commits_info_3_debug_fuType = RTL_PATH.io_commits_info_3_debug_fuType; \
        force U_IF_NAME.io_commits_info_3_dirtyFs = RTL_PATH.io_commits_info_3_dirtyFs; \
        force U_IF_NAME.io_commits_info_3_dirtyVs = RTL_PATH.io_commits_info_3_dirtyVs; \
        force U_IF_NAME.io_commits_info_4_walk_v = RTL_PATH.io_commits_info_4_walk_v; \
        force U_IF_NAME.io_commits_info_4_commit_v = RTL_PATH.io_commits_info_4_commit_v; \
        force U_IF_NAME.io_commits_info_4_commit_w = RTL_PATH.io_commits_info_4_commit_w; \
        force U_IF_NAME.io_commits_info_4_realDestSize = RTL_PATH.io_commits_info_4_realDestSize; \
        force U_IF_NAME.io_commits_info_4_interrupt_safe = RTL_PATH.io_commits_info_4_interrupt_safe; \
        force U_IF_NAME.io_commits_info_4_wflags = RTL_PATH.io_commits_info_4_wflags; \
        force U_IF_NAME.io_commits_info_4_fflags = RTL_PATH.io_commits_info_4_fflags; \
        force U_IF_NAME.io_commits_info_4_vxsat = RTL_PATH.io_commits_info_4_vxsat; \
        force U_IF_NAME.io_commits_info_4_isRVC = RTL_PATH.io_commits_info_4_isRVC; \
        force U_IF_NAME.io_commits_info_4_isVset = RTL_PATH.io_commits_info_4_isVset; \
        force U_IF_NAME.io_commits_info_4_isHls = RTL_PATH.io_commits_info_4_isHls; \
        force U_IF_NAME.io_commits_info_4_isVls = RTL_PATH.io_commits_info_4_isVls; \
        force U_IF_NAME.io_commits_info_4_vls = RTL_PATH.io_commits_info_4_vls; \
        force U_IF_NAME.io_commits_info_4_mmio = RTL_PATH.io_commits_info_4_mmio; \
        force U_IF_NAME.io_commits_info_4_commitType = RTL_PATH.io_commits_info_4_commitType; \
        force U_IF_NAME.io_commits_info_4_ftqIdx_flag = RTL_PATH.io_commits_info_4_ftqIdx_flag; \
        force U_IF_NAME.io_commits_info_4_ftqIdx_value = RTL_PATH.io_commits_info_4_ftqIdx_value; \
        force U_IF_NAME.io_commits_info_4_ftqOffset = RTL_PATH.io_commits_info_4_ftqOffset; \
        force U_IF_NAME.io_commits_info_4_instrSize = RTL_PATH.io_commits_info_4_instrSize; \
        force U_IF_NAME.io_commits_info_4_fpWen = RTL_PATH.io_commits_info_4_fpWen; \
        force U_IF_NAME.io_commits_info_4_rfWen = RTL_PATH.io_commits_info_4_rfWen; \
        force U_IF_NAME.io_commits_info_4_needFlush = RTL_PATH.io_commits_info_4_needFlush; \
        force U_IF_NAME.io_commits_info_4_traceBlockInPipe_itype = RTL_PATH.io_commits_info_4_traceBlockInPipe_itype; \
        force U_IF_NAME.io_commits_info_4_traceBlockInPipe_iretire = RTL_PATH.io_commits_info_4_traceBlockInPipe_iretire; \
        force U_IF_NAME.io_commits_info_4_traceBlockInPipe_ilastsize = RTL_PATH.io_commits_info_4_traceBlockInPipe_ilastsize; \
        force U_IF_NAME.io_commits_info_4_debug_pc = RTL_PATH.io_commits_info_4_debug_pc; \
        force U_IF_NAME.io_commits_info_4_debug_instr = RTL_PATH.io_commits_info_4_debug_instr; \
        force U_IF_NAME.io_commits_info_4_debug_ldest = RTL_PATH.io_commits_info_4_debug_ldest; \
        force U_IF_NAME.io_commits_info_4_debug_pdest = RTL_PATH.io_commits_info_4_debug_pdest; \
        force U_IF_NAME.io_commits_info_4_debug_otherPdest_0 = RTL_PATH.io_commits_info_4_debug_otherPdest_0; \
        force U_IF_NAME.io_commits_info_4_debug_otherPdest_1 = RTL_PATH.io_commits_info_4_debug_otherPdest_1; \
        force U_IF_NAME.io_commits_info_4_debug_otherPdest_2 = RTL_PATH.io_commits_info_4_debug_otherPdest_2; \
        force U_IF_NAME.io_commits_info_4_debug_otherPdest_3 = RTL_PATH.io_commits_info_4_debug_otherPdest_3; \
        force U_IF_NAME.io_commits_info_4_debug_otherPdest_4 = RTL_PATH.io_commits_info_4_debug_otherPdest_4; \
        force U_IF_NAME.io_commits_info_4_debug_otherPdest_5 = RTL_PATH.io_commits_info_4_debug_otherPdest_5; \
        force U_IF_NAME.io_commits_info_4_debug_otherPdest_6 = RTL_PATH.io_commits_info_4_debug_otherPdest_6; \
        force U_IF_NAME.io_commits_info_4_debug_fuType = RTL_PATH.io_commits_info_4_debug_fuType; \
        force U_IF_NAME.io_commits_info_4_dirtyFs = RTL_PATH.io_commits_info_4_dirtyFs; \
        force U_IF_NAME.io_commits_info_4_dirtyVs = RTL_PATH.io_commits_info_4_dirtyVs; \
        force U_IF_NAME.io_commits_info_5_walk_v = RTL_PATH.io_commits_info_5_walk_v; \
        force U_IF_NAME.io_commits_info_5_commit_v = RTL_PATH.io_commits_info_5_commit_v; \
        force U_IF_NAME.io_commits_info_5_commit_w = RTL_PATH.io_commits_info_5_commit_w; \
        force U_IF_NAME.io_commits_info_5_realDestSize = RTL_PATH.io_commits_info_5_realDestSize; \
        force U_IF_NAME.io_commits_info_5_interrupt_safe = RTL_PATH.io_commits_info_5_interrupt_safe; \
        force U_IF_NAME.io_commits_info_5_wflags = RTL_PATH.io_commits_info_5_wflags; \
        force U_IF_NAME.io_commits_info_5_fflags = RTL_PATH.io_commits_info_5_fflags; \
        force U_IF_NAME.io_commits_info_5_vxsat = RTL_PATH.io_commits_info_5_vxsat; \
        force U_IF_NAME.io_commits_info_5_isRVC = RTL_PATH.io_commits_info_5_isRVC; \
        force U_IF_NAME.io_commits_info_5_isVset = RTL_PATH.io_commits_info_5_isVset; \
        force U_IF_NAME.io_commits_info_5_isHls = RTL_PATH.io_commits_info_5_isHls; \
        force U_IF_NAME.io_commits_info_5_isVls = RTL_PATH.io_commits_info_5_isVls; \
        force U_IF_NAME.io_commits_info_5_vls = RTL_PATH.io_commits_info_5_vls; \
        force U_IF_NAME.io_commits_info_5_mmio = RTL_PATH.io_commits_info_5_mmio; \
        force U_IF_NAME.io_commits_info_5_commitType = RTL_PATH.io_commits_info_5_commitType; \
        force U_IF_NAME.io_commits_info_5_ftqIdx_flag = RTL_PATH.io_commits_info_5_ftqIdx_flag; \
        force U_IF_NAME.io_commits_info_5_ftqIdx_value = RTL_PATH.io_commits_info_5_ftqIdx_value; \
        force U_IF_NAME.io_commits_info_5_ftqOffset = RTL_PATH.io_commits_info_5_ftqOffset; \
        force U_IF_NAME.io_commits_info_5_instrSize = RTL_PATH.io_commits_info_5_instrSize; \
        force U_IF_NAME.io_commits_info_5_fpWen = RTL_PATH.io_commits_info_5_fpWen; \
        force U_IF_NAME.io_commits_info_5_rfWen = RTL_PATH.io_commits_info_5_rfWen; \
        force U_IF_NAME.io_commits_info_5_needFlush = RTL_PATH.io_commits_info_5_needFlush; \
        force U_IF_NAME.io_commits_info_5_traceBlockInPipe_itype = RTL_PATH.io_commits_info_5_traceBlockInPipe_itype; \
        force U_IF_NAME.io_commits_info_5_traceBlockInPipe_iretire = RTL_PATH.io_commits_info_5_traceBlockInPipe_iretire; \
        force U_IF_NAME.io_commits_info_5_traceBlockInPipe_ilastsize = RTL_PATH.io_commits_info_5_traceBlockInPipe_ilastsize; \
        force U_IF_NAME.io_commits_info_5_debug_pc = RTL_PATH.io_commits_info_5_debug_pc; \
        force U_IF_NAME.io_commits_info_5_debug_instr = RTL_PATH.io_commits_info_5_debug_instr; \
        force U_IF_NAME.io_commits_info_5_debug_ldest = RTL_PATH.io_commits_info_5_debug_ldest; \
        force U_IF_NAME.io_commits_info_5_debug_pdest = RTL_PATH.io_commits_info_5_debug_pdest; \
        force U_IF_NAME.io_commits_info_5_debug_otherPdest_0 = RTL_PATH.io_commits_info_5_debug_otherPdest_0; \
        force U_IF_NAME.io_commits_info_5_debug_otherPdest_1 = RTL_PATH.io_commits_info_5_debug_otherPdest_1; \
        force U_IF_NAME.io_commits_info_5_debug_otherPdest_2 = RTL_PATH.io_commits_info_5_debug_otherPdest_2; \
        force U_IF_NAME.io_commits_info_5_debug_otherPdest_3 = RTL_PATH.io_commits_info_5_debug_otherPdest_3; \
        force U_IF_NAME.io_commits_info_5_debug_otherPdest_4 = RTL_PATH.io_commits_info_5_debug_otherPdest_4; \
        force U_IF_NAME.io_commits_info_5_debug_otherPdest_5 = RTL_PATH.io_commits_info_5_debug_otherPdest_5; \
        force U_IF_NAME.io_commits_info_5_debug_otherPdest_6 = RTL_PATH.io_commits_info_5_debug_otherPdest_6; \
        force U_IF_NAME.io_commits_info_5_debug_fuType = RTL_PATH.io_commits_info_5_debug_fuType; \
        force U_IF_NAME.io_commits_info_5_dirtyFs = RTL_PATH.io_commits_info_5_dirtyFs; \
        force U_IF_NAME.io_commits_info_5_dirtyVs = RTL_PATH.io_commits_info_5_dirtyVs; \
        force U_IF_NAME.io_commits_info_6_walk_v = RTL_PATH.io_commits_info_6_walk_v; \
        force U_IF_NAME.io_commits_info_6_commit_v = RTL_PATH.io_commits_info_6_commit_v; \
        force U_IF_NAME.io_commits_info_6_commit_w = RTL_PATH.io_commits_info_6_commit_w; \
        force U_IF_NAME.io_commits_info_6_realDestSize = RTL_PATH.io_commits_info_6_realDestSize; \
        force U_IF_NAME.io_commits_info_6_interrupt_safe = RTL_PATH.io_commits_info_6_interrupt_safe; \
        force U_IF_NAME.io_commits_info_6_wflags = RTL_PATH.io_commits_info_6_wflags; \
        force U_IF_NAME.io_commits_info_6_fflags = RTL_PATH.io_commits_info_6_fflags; \
        force U_IF_NAME.io_commits_info_6_vxsat = RTL_PATH.io_commits_info_6_vxsat; \
        force U_IF_NAME.io_commits_info_6_isRVC = RTL_PATH.io_commits_info_6_isRVC; \
        force U_IF_NAME.io_commits_info_6_isVset = RTL_PATH.io_commits_info_6_isVset; \
        force U_IF_NAME.io_commits_info_6_isHls = RTL_PATH.io_commits_info_6_isHls; \
        force U_IF_NAME.io_commits_info_6_isVls = RTL_PATH.io_commits_info_6_isVls; \
        force U_IF_NAME.io_commits_info_6_vls = RTL_PATH.io_commits_info_6_vls; \
        force U_IF_NAME.io_commits_info_6_mmio = RTL_PATH.io_commits_info_6_mmio; \
        force U_IF_NAME.io_commits_info_6_commitType = RTL_PATH.io_commits_info_6_commitType; \
        force U_IF_NAME.io_commits_info_6_ftqIdx_flag = RTL_PATH.io_commits_info_6_ftqIdx_flag; \
        force U_IF_NAME.io_commits_info_6_ftqIdx_value = RTL_PATH.io_commits_info_6_ftqIdx_value; \
        force U_IF_NAME.io_commits_info_6_ftqOffset = RTL_PATH.io_commits_info_6_ftqOffset; \
        force U_IF_NAME.io_commits_info_6_instrSize = RTL_PATH.io_commits_info_6_instrSize; \
        force U_IF_NAME.io_commits_info_6_fpWen = RTL_PATH.io_commits_info_6_fpWen; \
        force U_IF_NAME.io_commits_info_6_rfWen = RTL_PATH.io_commits_info_6_rfWen; \
        force U_IF_NAME.io_commits_info_6_needFlush = RTL_PATH.io_commits_info_6_needFlush; \
        force U_IF_NAME.io_commits_info_6_traceBlockInPipe_itype = RTL_PATH.io_commits_info_6_traceBlockInPipe_itype; \
        force U_IF_NAME.io_commits_info_6_traceBlockInPipe_iretire = RTL_PATH.io_commits_info_6_traceBlockInPipe_iretire; \
        force U_IF_NAME.io_commits_info_6_traceBlockInPipe_ilastsize = RTL_PATH.io_commits_info_6_traceBlockInPipe_ilastsize; \
        force U_IF_NAME.io_commits_info_6_debug_pc = RTL_PATH.io_commits_info_6_debug_pc; \
        force U_IF_NAME.io_commits_info_6_debug_instr = RTL_PATH.io_commits_info_6_debug_instr; \
        force U_IF_NAME.io_commits_info_6_debug_ldest = RTL_PATH.io_commits_info_6_debug_ldest; \
        force U_IF_NAME.io_commits_info_6_debug_pdest = RTL_PATH.io_commits_info_6_debug_pdest; \
        force U_IF_NAME.io_commits_info_6_debug_otherPdest_0 = RTL_PATH.io_commits_info_6_debug_otherPdest_0; \
        force U_IF_NAME.io_commits_info_6_debug_otherPdest_1 = RTL_PATH.io_commits_info_6_debug_otherPdest_1; \
        force U_IF_NAME.io_commits_info_6_debug_otherPdest_2 = RTL_PATH.io_commits_info_6_debug_otherPdest_2; \
        force U_IF_NAME.io_commits_info_6_debug_otherPdest_3 = RTL_PATH.io_commits_info_6_debug_otherPdest_3; \
        force U_IF_NAME.io_commits_info_6_debug_otherPdest_4 = RTL_PATH.io_commits_info_6_debug_otherPdest_4; \
        force U_IF_NAME.io_commits_info_6_debug_otherPdest_5 = RTL_PATH.io_commits_info_6_debug_otherPdest_5; \
        force U_IF_NAME.io_commits_info_6_debug_otherPdest_6 = RTL_PATH.io_commits_info_6_debug_otherPdest_6; \
        force U_IF_NAME.io_commits_info_6_debug_fuType = RTL_PATH.io_commits_info_6_debug_fuType; \
        force U_IF_NAME.io_commits_info_6_dirtyFs = RTL_PATH.io_commits_info_6_dirtyFs; \
        force U_IF_NAME.io_commits_info_6_dirtyVs = RTL_PATH.io_commits_info_6_dirtyVs; \
        force U_IF_NAME.io_commits_info_7_walk_v = RTL_PATH.io_commits_info_7_walk_v; \
        force U_IF_NAME.io_commits_info_7_commit_v = RTL_PATH.io_commits_info_7_commit_v; \
        force U_IF_NAME.io_commits_info_7_commit_w = RTL_PATH.io_commits_info_7_commit_w; \
        force U_IF_NAME.io_commits_info_7_realDestSize = RTL_PATH.io_commits_info_7_realDestSize; \
        force U_IF_NAME.io_commits_info_7_interrupt_safe = RTL_PATH.io_commits_info_7_interrupt_safe; \
        force U_IF_NAME.io_commits_info_7_wflags = RTL_PATH.io_commits_info_7_wflags; \
        force U_IF_NAME.io_commits_info_7_fflags = RTL_PATH.io_commits_info_7_fflags; \
        force U_IF_NAME.io_commits_info_7_vxsat = RTL_PATH.io_commits_info_7_vxsat; \
        force U_IF_NAME.io_commits_info_7_isRVC = RTL_PATH.io_commits_info_7_isRVC; \
        force U_IF_NAME.io_commits_info_7_isVset = RTL_PATH.io_commits_info_7_isVset; \
        force U_IF_NAME.io_commits_info_7_isHls = RTL_PATH.io_commits_info_7_isHls; \
        force U_IF_NAME.io_commits_info_7_isVls = RTL_PATH.io_commits_info_7_isVls; \
        force U_IF_NAME.io_commits_info_7_vls = RTL_PATH.io_commits_info_7_vls; \
        force U_IF_NAME.io_commits_info_7_mmio = RTL_PATH.io_commits_info_7_mmio; \
        force U_IF_NAME.io_commits_info_7_commitType = RTL_PATH.io_commits_info_7_commitType; \
        force U_IF_NAME.io_commits_info_7_ftqIdx_flag = RTL_PATH.io_commits_info_7_ftqIdx_flag; \
        force U_IF_NAME.io_commits_info_7_ftqIdx_value = RTL_PATH.io_commits_info_7_ftqIdx_value; \
        force U_IF_NAME.io_commits_info_7_ftqOffset = RTL_PATH.io_commits_info_7_ftqOffset; \
        force U_IF_NAME.io_commits_info_7_instrSize = RTL_PATH.io_commits_info_7_instrSize; \
        force U_IF_NAME.io_commits_info_7_fpWen = RTL_PATH.io_commits_info_7_fpWen; \
        force U_IF_NAME.io_commits_info_7_rfWen = RTL_PATH.io_commits_info_7_rfWen; \
        force U_IF_NAME.io_commits_info_7_needFlush = RTL_PATH.io_commits_info_7_needFlush; \
        force U_IF_NAME.io_commits_info_7_traceBlockInPipe_itype = RTL_PATH.io_commits_info_7_traceBlockInPipe_itype; \
        force U_IF_NAME.io_commits_info_7_traceBlockInPipe_iretire = RTL_PATH.io_commits_info_7_traceBlockInPipe_iretire; \
        force U_IF_NAME.io_commits_info_7_traceBlockInPipe_ilastsize = RTL_PATH.io_commits_info_7_traceBlockInPipe_ilastsize; \
        force U_IF_NAME.io_commits_info_7_debug_pc = RTL_PATH.io_commits_info_7_debug_pc; \
        force U_IF_NAME.io_commits_info_7_debug_instr = RTL_PATH.io_commits_info_7_debug_instr; \
        force U_IF_NAME.io_commits_info_7_debug_ldest = RTL_PATH.io_commits_info_7_debug_ldest; \
        force U_IF_NAME.io_commits_info_7_debug_pdest = RTL_PATH.io_commits_info_7_debug_pdest; \
        force U_IF_NAME.io_commits_info_7_debug_otherPdest_0 = RTL_PATH.io_commits_info_7_debug_otherPdest_0; \
        force U_IF_NAME.io_commits_info_7_debug_otherPdest_1 = RTL_PATH.io_commits_info_7_debug_otherPdest_1; \
        force U_IF_NAME.io_commits_info_7_debug_otherPdest_2 = RTL_PATH.io_commits_info_7_debug_otherPdest_2; \
        force U_IF_NAME.io_commits_info_7_debug_otherPdest_3 = RTL_PATH.io_commits_info_7_debug_otherPdest_3; \
        force U_IF_NAME.io_commits_info_7_debug_otherPdest_4 = RTL_PATH.io_commits_info_7_debug_otherPdest_4; \
        force U_IF_NAME.io_commits_info_7_debug_otherPdest_5 = RTL_PATH.io_commits_info_7_debug_otherPdest_5; \
        force U_IF_NAME.io_commits_info_7_debug_otherPdest_6 = RTL_PATH.io_commits_info_7_debug_otherPdest_6; \
        force U_IF_NAME.io_commits_info_7_debug_fuType = RTL_PATH.io_commits_info_7_debug_fuType; \
        force U_IF_NAME.io_commits_info_7_dirtyFs = RTL_PATH.io_commits_info_7_dirtyFs; \
        force U_IF_NAME.io_commits_info_7_dirtyVs = RTL_PATH.io_commits_info_7_dirtyVs; \
        force U_IF_NAME.io_commits_robIdx_0_flag = RTL_PATH.io_commits_robIdx_0_flag; \
        force U_IF_NAME.io_commits_robIdx_0_value = RTL_PATH.io_commits_robIdx_0_value; \
        force U_IF_NAME.io_commits_robIdx_1_flag = RTL_PATH.io_commits_robIdx_1_flag; \
        force U_IF_NAME.io_commits_robIdx_1_value = RTL_PATH.io_commits_robIdx_1_value; \
        force U_IF_NAME.io_commits_robIdx_2_flag = RTL_PATH.io_commits_robIdx_2_flag; \
        force U_IF_NAME.io_commits_robIdx_2_value = RTL_PATH.io_commits_robIdx_2_value; \
        force U_IF_NAME.io_commits_robIdx_3_flag = RTL_PATH.io_commits_robIdx_3_flag; \
        force U_IF_NAME.io_commits_robIdx_3_value = RTL_PATH.io_commits_robIdx_3_value; \
        force U_IF_NAME.io_commits_robIdx_4_flag = RTL_PATH.io_commits_robIdx_4_flag; \
        force U_IF_NAME.io_commits_robIdx_4_value = RTL_PATH.io_commits_robIdx_4_value; \
        force U_IF_NAME.io_commits_robIdx_5_flag = RTL_PATH.io_commits_robIdx_5_flag; \
        force U_IF_NAME.io_commits_robIdx_5_value = RTL_PATH.io_commits_robIdx_5_value; \
        force U_IF_NAME.io_commits_robIdx_6_flag = RTL_PATH.io_commits_robIdx_6_flag; \
        force U_IF_NAME.io_commits_robIdx_6_value = RTL_PATH.io_commits_robIdx_6_value; \
        force U_IF_NAME.io_commits_robIdx_7_flag = RTL_PATH.io_commits_robIdx_7_flag; \
        force U_IF_NAME.io_commits_robIdx_7_value = RTL_PATH.io_commits_robIdx_7_value; \
        force RTL_PATH.io_trace_blockCommit = U_IF_NAME.io_trace_blockCommit; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_0_valid = RTL_PATH.io_trace_traceCommitInfo_blocks_0_valid; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value = RTL_PATH.io_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_0_bits_ftqOffset = RTL_PATH.io_trace_traceCommitInfo_blocks_0_bits_ftqOffset; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype = RTL_PATH.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire = RTL_PATH.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize = RTL_PATH.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_1_valid = RTL_PATH.io_trace_traceCommitInfo_blocks_1_valid; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value = RTL_PATH.io_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_1_bits_ftqOffset = RTL_PATH.io_trace_traceCommitInfo_blocks_1_bits_ftqOffset; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype = RTL_PATH.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire = RTL_PATH.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize = RTL_PATH.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_2_valid = RTL_PATH.io_trace_traceCommitInfo_blocks_2_valid; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value = RTL_PATH.io_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_2_bits_ftqOffset = RTL_PATH.io_trace_traceCommitInfo_blocks_2_bits_ftqOffset; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype = RTL_PATH.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire = RTL_PATH.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize = RTL_PATH.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_3_valid = RTL_PATH.io_trace_traceCommitInfo_blocks_3_valid; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value = RTL_PATH.io_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_3_bits_ftqOffset = RTL_PATH.io_trace_traceCommitInfo_blocks_3_bits_ftqOffset; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype = RTL_PATH.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire = RTL_PATH.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize = RTL_PATH.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_4_valid = RTL_PATH.io_trace_traceCommitInfo_blocks_4_valid; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value = RTL_PATH.io_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_4_bits_ftqOffset = RTL_PATH.io_trace_traceCommitInfo_blocks_4_bits_ftqOffset; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype = RTL_PATH.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire = RTL_PATH.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize = RTL_PATH.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_5_valid = RTL_PATH.io_trace_traceCommitInfo_blocks_5_valid; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value = RTL_PATH.io_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_5_bits_ftqOffset = RTL_PATH.io_trace_traceCommitInfo_blocks_5_bits_ftqOffset; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype = RTL_PATH.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire = RTL_PATH.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize = RTL_PATH.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_6_valid = RTL_PATH.io_trace_traceCommitInfo_blocks_6_valid; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value = RTL_PATH.io_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_6_bits_ftqOffset = RTL_PATH.io_trace_traceCommitInfo_blocks_6_bits_ftqOffset; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype = RTL_PATH.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire = RTL_PATH.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize = RTL_PATH.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_7_valid = RTL_PATH.io_trace_traceCommitInfo_blocks_7_valid; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value = RTL_PATH.io_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_7_bits_ftqOffset = RTL_PATH.io_trace_traceCommitInfo_blocks_7_bits_ftqOffset; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype = RTL_PATH.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire = RTL_PATH.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize = RTL_PATH.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize; \
        force U_IF_NAME.io_rabCommits_isCommit = RTL_PATH.io_rabCommits_isCommit; \
        force U_IF_NAME.io_rabCommits_commitValid_0 = RTL_PATH.io_rabCommits_commitValid_0; \
        force U_IF_NAME.io_rabCommits_commitValid_1 = RTL_PATH.io_rabCommits_commitValid_1; \
        force U_IF_NAME.io_rabCommits_commitValid_2 = RTL_PATH.io_rabCommits_commitValid_2; \
        force U_IF_NAME.io_rabCommits_commitValid_3 = RTL_PATH.io_rabCommits_commitValid_3; \
        force U_IF_NAME.io_rabCommits_commitValid_4 = RTL_PATH.io_rabCommits_commitValid_4; \
        force U_IF_NAME.io_rabCommits_commitValid_5 = RTL_PATH.io_rabCommits_commitValid_5; \
        force U_IF_NAME.io_rabCommits_isWalk = RTL_PATH.io_rabCommits_isWalk; \
        force U_IF_NAME.io_rabCommits_walkValid_0 = RTL_PATH.io_rabCommits_walkValid_0; \
        force U_IF_NAME.io_rabCommits_walkValid_1 = RTL_PATH.io_rabCommits_walkValid_1; \
        force U_IF_NAME.io_rabCommits_walkValid_2 = RTL_PATH.io_rabCommits_walkValid_2; \
        force U_IF_NAME.io_rabCommits_walkValid_3 = RTL_PATH.io_rabCommits_walkValid_3; \
        force U_IF_NAME.io_rabCommits_walkValid_4 = RTL_PATH.io_rabCommits_walkValid_4; \
        force U_IF_NAME.io_rabCommits_walkValid_5 = RTL_PATH.io_rabCommits_walkValid_5; \
        force U_IF_NAME.io_rabCommits_info_0_ldest = RTL_PATH.io_rabCommits_info_0_ldest; \
        force U_IF_NAME.io_rabCommits_info_0_pdest = RTL_PATH.io_rabCommits_info_0_pdest; \
        force U_IF_NAME.io_rabCommits_info_0_rfWen = RTL_PATH.io_rabCommits_info_0_rfWen; \
        force U_IF_NAME.io_rabCommits_info_0_fpWen = RTL_PATH.io_rabCommits_info_0_fpWen; \
        force U_IF_NAME.io_rabCommits_info_0_vecWen = RTL_PATH.io_rabCommits_info_0_vecWen; \
        force U_IF_NAME.io_rabCommits_info_0_v0Wen = RTL_PATH.io_rabCommits_info_0_v0Wen; \
        force U_IF_NAME.io_rabCommits_info_0_vlWen = RTL_PATH.io_rabCommits_info_0_vlWen; \
        force U_IF_NAME.io_rabCommits_info_0_isMove = RTL_PATH.io_rabCommits_info_0_isMove; \
        force U_IF_NAME.io_rabCommits_info_1_ldest = RTL_PATH.io_rabCommits_info_1_ldest; \
        force U_IF_NAME.io_rabCommits_info_1_pdest = RTL_PATH.io_rabCommits_info_1_pdest; \
        force U_IF_NAME.io_rabCommits_info_1_rfWen = RTL_PATH.io_rabCommits_info_1_rfWen; \
        force U_IF_NAME.io_rabCommits_info_1_fpWen = RTL_PATH.io_rabCommits_info_1_fpWen; \
        force U_IF_NAME.io_rabCommits_info_1_vecWen = RTL_PATH.io_rabCommits_info_1_vecWen; \
        force U_IF_NAME.io_rabCommits_info_1_v0Wen = RTL_PATH.io_rabCommits_info_1_v0Wen; \
        force U_IF_NAME.io_rabCommits_info_1_vlWen = RTL_PATH.io_rabCommits_info_1_vlWen; \
        force U_IF_NAME.io_rabCommits_info_1_isMove = RTL_PATH.io_rabCommits_info_1_isMove; \
        force U_IF_NAME.io_rabCommits_info_2_ldest = RTL_PATH.io_rabCommits_info_2_ldest; \
        force U_IF_NAME.io_rabCommits_info_2_pdest = RTL_PATH.io_rabCommits_info_2_pdest; \
        force U_IF_NAME.io_rabCommits_info_2_rfWen = RTL_PATH.io_rabCommits_info_2_rfWen; \
        force U_IF_NAME.io_rabCommits_info_2_fpWen = RTL_PATH.io_rabCommits_info_2_fpWen; \
        force U_IF_NAME.io_rabCommits_info_2_vecWen = RTL_PATH.io_rabCommits_info_2_vecWen; \
        force U_IF_NAME.io_rabCommits_info_2_v0Wen = RTL_PATH.io_rabCommits_info_2_v0Wen; \
        force U_IF_NAME.io_rabCommits_info_2_vlWen = RTL_PATH.io_rabCommits_info_2_vlWen; \
        force U_IF_NAME.io_rabCommits_info_2_isMove = RTL_PATH.io_rabCommits_info_2_isMove; \
        force U_IF_NAME.io_rabCommits_info_3_ldest = RTL_PATH.io_rabCommits_info_3_ldest; \
        force U_IF_NAME.io_rabCommits_info_3_pdest = RTL_PATH.io_rabCommits_info_3_pdest; \
        force U_IF_NAME.io_rabCommits_info_3_rfWen = RTL_PATH.io_rabCommits_info_3_rfWen; \
        force U_IF_NAME.io_rabCommits_info_3_fpWen = RTL_PATH.io_rabCommits_info_3_fpWen; \
        force U_IF_NAME.io_rabCommits_info_3_vecWen = RTL_PATH.io_rabCommits_info_3_vecWen; \
        force U_IF_NAME.io_rabCommits_info_3_v0Wen = RTL_PATH.io_rabCommits_info_3_v0Wen; \
        force U_IF_NAME.io_rabCommits_info_3_vlWen = RTL_PATH.io_rabCommits_info_3_vlWen; \
        force U_IF_NAME.io_rabCommits_info_3_isMove = RTL_PATH.io_rabCommits_info_3_isMove; \
        force U_IF_NAME.io_rabCommits_info_4_ldest = RTL_PATH.io_rabCommits_info_4_ldest; \
        force U_IF_NAME.io_rabCommits_info_4_pdest = RTL_PATH.io_rabCommits_info_4_pdest; \
        force U_IF_NAME.io_rabCommits_info_4_rfWen = RTL_PATH.io_rabCommits_info_4_rfWen; \
        force U_IF_NAME.io_rabCommits_info_4_fpWen = RTL_PATH.io_rabCommits_info_4_fpWen; \
        force U_IF_NAME.io_rabCommits_info_4_vecWen = RTL_PATH.io_rabCommits_info_4_vecWen; \
        force U_IF_NAME.io_rabCommits_info_4_v0Wen = RTL_PATH.io_rabCommits_info_4_v0Wen; \
        force U_IF_NAME.io_rabCommits_info_4_vlWen = RTL_PATH.io_rabCommits_info_4_vlWen; \
        force U_IF_NAME.io_rabCommits_info_4_isMove = RTL_PATH.io_rabCommits_info_4_isMove; \
        force U_IF_NAME.io_rabCommits_info_5_ldest = RTL_PATH.io_rabCommits_info_5_ldest; \
        force U_IF_NAME.io_rabCommits_info_5_pdest = RTL_PATH.io_rabCommits_info_5_pdest; \
        force U_IF_NAME.io_rabCommits_info_5_rfWen = RTL_PATH.io_rabCommits_info_5_rfWen; \
        force U_IF_NAME.io_rabCommits_info_5_fpWen = RTL_PATH.io_rabCommits_info_5_fpWen; \
        force U_IF_NAME.io_rabCommits_info_5_vecWen = RTL_PATH.io_rabCommits_info_5_vecWen; \
        force U_IF_NAME.io_rabCommits_info_5_v0Wen = RTL_PATH.io_rabCommits_info_5_v0Wen; \
        force U_IF_NAME.io_rabCommits_info_5_vlWen = RTL_PATH.io_rabCommits_info_5_vlWen; \
        force U_IF_NAME.io_rabCommits_info_5_isMove = RTL_PATH.io_rabCommits_info_5_isMove; \
        force U_IF_NAME.io_diffCommits_commitValid_0 = RTL_PATH.io_diffCommits_commitValid_0; \
        force U_IF_NAME.io_diffCommits_commitValid_1 = RTL_PATH.io_diffCommits_commitValid_1; \
        force U_IF_NAME.io_diffCommits_commitValid_2 = RTL_PATH.io_diffCommits_commitValid_2; \
        force U_IF_NAME.io_diffCommits_commitValid_3 = RTL_PATH.io_diffCommits_commitValid_3; \
        force U_IF_NAME.io_diffCommits_commitValid_4 = RTL_PATH.io_diffCommits_commitValid_4; \
        force U_IF_NAME.io_diffCommits_commitValid_5 = RTL_PATH.io_diffCommits_commitValid_5; \
        force U_IF_NAME.io_diffCommits_commitValid_6 = RTL_PATH.io_diffCommits_commitValid_6; \
        force U_IF_NAME.io_diffCommits_commitValid_7 = RTL_PATH.io_diffCommits_commitValid_7; \
        force U_IF_NAME.io_diffCommits_commitValid_8 = RTL_PATH.io_diffCommits_commitValid_8; \
        force U_IF_NAME.io_diffCommits_commitValid_9 = RTL_PATH.io_diffCommits_commitValid_9; \
        force U_IF_NAME.io_diffCommits_commitValid_10 = RTL_PATH.io_diffCommits_commitValid_10; \
        force U_IF_NAME.io_diffCommits_commitValid_11 = RTL_PATH.io_diffCommits_commitValid_11; \
        force U_IF_NAME.io_diffCommits_commitValid_12 = RTL_PATH.io_diffCommits_commitValid_12; \
        force U_IF_NAME.io_diffCommits_commitValid_13 = RTL_PATH.io_diffCommits_commitValid_13; \
        force U_IF_NAME.io_diffCommits_commitValid_14 = RTL_PATH.io_diffCommits_commitValid_14; \
        force U_IF_NAME.io_diffCommits_commitValid_15 = RTL_PATH.io_diffCommits_commitValid_15; \
        force U_IF_NAME.io_diffCommits_commitValid_16 = RTL_PATH.io_diffCommits_commitValid_16; \
        force U_IF_NAME.io_diffCommits_commitValid_17 = RTL_PATH.io_diffCommits_commitValid_17; \
        force U_IF_NAME.io_diffCommits_commitValid_18 = RTL_PATH.io_diffCommits_commitValid_18; \
        force U_IF_NAME.io_diffCommits_commitValid_19 = RTL_PATH.io_diffCommits_commitValid_19; \
        force U_IF_NAME.io_diffCommits_commitValid_20 = RTL_PATH.io_diffCommits_commitValid_20; \
        force U_IF_NAME.io_diffCommits_commitValid_21 = RTL_PATH.io_diffCommits_commitValid_21; \
        force U_IF_NAME.io_diffCommits_commitValid_22 = RTL_PATH.io_diffCommits_commitValid_22; \
        force U_IF_NAME.io_diffCommits_commitValid_23 = RTL_PATH.io_diffCommits_commitValid_23; \
        force U_IF_NAME.io_diffCommits_commitValid_24 = RTL_PATH.io_diffCommits_commitValid_24; \
        force U_IF_NAME.io_diffCommits_commitValid_25 = RTL_PATH.io_diffCommits_commitValid_25; \
        force U_IF_NAME.io_diffCommits_commitValid_26 = RTL_PATH.io_diffCommits_commitValid_26; \
        force U_IF_NAME.io_diffCommits_commitValid_27 = RTL_PATH.io_diffCommits_commitValid_27; \
        force U_IF_NAME.io_diffCommits_commitValid_28 = RTL_PATH.io_diffCommits_commitValid_28; \
        force U_IF_NAME.io_diffCommits_commitValid_29 = RTL_PATH.io_diffCommits_commitValid_29; \
        force U_IF_NAME.io_diffCommits_commitValid_30 = RTL_PATH.io_diffCommits_commitValid_30; \
        force U_IF_NAME.io_diffCommits_commitValid_31 = RTL_PATH.io_diffCommits_commitValid_31; \
        force U_IF_NAME.io_diffCommits_commitValid_32 = RTL_PATH.io_diffCommits_commitValid_32; \
        force U_IF_NAME.io_diffCommits_commitValid_33 = RTL_PATH.io_diffCommits_commitValid_33; \
        force U_IF_NAME.io_diffCommits_commitValid_34 = RTL_PATH.io_diffCommits_commitValid_34; \
        force U_IF_NAME.io_diffCommits_commitValid_35 = RTL_PATH.io_diffCommits_commitValid_35; \
        force U_IF_NAME.io_diffCommits_commitValid_36 = RTL_PATH.io_diffCommits_commitValid_36; \
        force U_IF_NAME.io_diffCommits_commitValid_37 = RTL_PATH.io_diffCommits_commitValid_37; \
        force U_IF_NAME.io_diffCommits_commitValid_38 = RTL_PATH.io_diffCommits_commitValid_38; \
        force U_IF_NAME.io_diffCommits_commitValid_39 = RTL_PATH.io_diffCommits_commitValid_39; \
        force U_IF_NAME.io_diffCommits_commitValid_40 = RTL_PATH.io_diffCommits_commitValid_40; \
        force U_IF_NAME.io_diffCommits_commitValid_41 = RTL_PATH.io_diffCommits_commitValid_41; \
        force U_IF_NAME.io_diffCommits_commitValid_42 = RTL_PATH.io_diffCommits_commitValid_42; \
        force U_IF_NAME.io_diffCommits_commitValid_43 = RTL_PATH.io_diffCommits_commitValid_43; \
        force U_IF_NAME.io_diffCommits_commitValid_44 = RTL_PATH.io_diffCommits_commitValid_44; \
        force U_IF_NAME.io_diffCommits_commitValid_45 = RTL_PATH.io_diffCommits_commitValid_45; \
        force U_IF_NAME.io_diffCommits_commitValid_46 = RTL_PATH.io_diffCommits_commitValid_46; \
        force U_IF_NAME.io_diffCommits_commitValid_47 = RTL_PATH.io_diffCommits_commitValid_47; \
        force U_IF_NAME.io_diffCommits_commitValid_48 = RTL_PATH.io_diffCommits_commitValid_48; \
        force U_IF_NAME.io_diffCommits_commitValid_49 = RTL_PATH.io_diffCommits_commitValid_49; \
        force U_IF_NAME.io_diffCommits_commitValid_50 = RTL_PATH.io_diffCommits_commitValid_50; \
        force U_IF_NAME.io_diffCommits_commitValid_51 = RTL_PATH.io_diffCommits_commitValid_51; \
        force U_IF_NAME.io_diffCommits_commitValid_52 = RTL_PATH.io_diffCommits_commitValid_52; \
        force U_IF_NAME.io_diffCommits_commitValid_53 = RTL_PATH.io_diffCommits_commitValid_53; \
        force U_IF_NAME.io_diffCommits_commitValid_54 = RTL_PATH.io_diffCommits_commitValid_54; \
        force U_IF_NAME.io_diffCommits_commitValid_55 = RTL_PATH.io_diffCommits_commitValid_55; \
        force U_IF_NAME.io_diffCommits_commitValid_56 = RTL_PATH.io_diffCommits_commitValid_56; \
        force U_IF_NAME.io_diffCommits_commitValid_57 = RTL_PATH.io_diffCommits_commitValid_57; \
        force U_IF_NAME.io_diffCommits_commitValid_58 = RTL_PATH.io_diffCommits_commitValid_58; \
        force U_IF_NAME.io_diffCommits_commitValid_59 = RTL_PATH.io_diffCommits_commitValid_59; \
        force U_IF_NAME.io_diffCommits_commitValid_60 = RTL_PATH.io_diffCommits_commitValid_60; \
        force U_IF_NAME.io_diffCommits_commitValid_61 = RTL_PATH.io_diffCommits_commitValid_61; \
        force U_IF_NAME.io_diffCommits_commitValid_62 = RTL_PATH.io_diffCommits_commitValid_62; \
        force U_IF_NAME.io_diffCommits_commitValid_63 = RTL_PATH.io_diffCommits_commitValid_63; \
        force U_IF_NAME.io_diffCommits_commitValid_64 = RTL_PATH.io_diffCommits_commitValid_64; \
        force U_IF_NAME.io_diffCommits_commitValid_65 = RTL_PATH.io_diffCommits_commitValid_65; \
        force U_IF_NAME.io_diffCommits_commitValid_66 = RTL_PATH.io_diffCommits_commitValid_66; \
        force U_IF_NAME.io_diffCommits_commitValid_67 = RTL_PATH.io_diffCommits_commitValid_67; \
        force U_IF_NAME.io_diffCommits_commitValid_68 = RTL_PATH.io_diffCommits_commitValid_68; \
        force U_IF_NAME.io_diffCommits_commitValid_69 = RTL_PATH.io_diffCommits_commitValid_69; \
        force U_IF_NAME.io_diffCommits_commitValid_70 = RTL_PATH.io_diffCommits_commitValid_70; \
        force U_IF_NAME.io_diffCommits_commitValid_71 = RTL_PATH.io_diffCommits_commitValid_71; \
        force U_IF_NAME.io_diffCommits_commitValid_72 = RTL_PATH.io_diffCommits_commitValid_72; \
        force U_IF_NAME.io_diffCommits_commitValid_73 = RTL_PATH.io_diffCommits_commitValid_73; \
        force U_IF_NAME.io_diffCommits_commitValid_74 = RTL_PATH.io_diffCommits_commitValid_74; \
        force U_IF_NAME.io_diffCommits_commitValid_75 = RTL_PATH.io_diffCommits_commitValid_75; \
        force U_IF_NAME.io_diffCommits_commitValid_76 = RTL_PATH.io_diffCommits_commitValid_76; \
        force U_IF_NAME.io_diffCommits_commitValid_77 = RTL_PATH.io_diffCommits_commitValid_77; \
        force U_IF_NAME.io_diffCommits_commitValid_78 = RTL_PATH.io_diffCommits_commitValid_78; \
        force U_IF_NAME.io_diffCommits_commitValid_79 = RTL_PATH.io_diffCommits_commitValid_79; \
        force U_IF_NAME.io_diffCommits_commitValid_80 = RTL_PATH.io_diffCommits_commitValid_80; \
        force U_IF_NAME.io_diffCommits_commitValid_81 = RTL_PATH.io_diffCommits_commitValid_81; \
        force U_IF_NAME.io_diffCommits_commitValid_82 = RTL_PATH.io_diffCommits_commitValid_82; \
        force U_IF_NAME.io_diffCommits_commitValid_83 = RTL_PATH.io_diffCommits_commitValid_83; \
        force U_IF_NAME.io_diffCommits_commitValid_84 = RTL_PATH.io_diffCommits_commitValid_84; \
        force U_IF_NAME.io_diffCommits_commitValid_85 = RTL_PATH.io_diffCommits_commitValid_85; \
        force U_IF_NAME.io_diffCommits_commitValid_86 = RTL_PATH.io_diffCommits_commitValid_86; \
        force U_IF_NAME.io_diffCommits_commitValid_87 = RTL_PATH.io_diffCommits_commitValid_87; \
        force U_IF_NAME.io_diffCommits_commitValid_88 = RTL_PATH.io_diffCommits_commitValid_88; \
        force U_IF_NAME.io_diffCommits_commitValid_89 = RTL_PATH.io_diffCommits_commitValid_89; \
        force U_IF_NAME.io_diffCommits_commitValid_90 = RTL_PATH.io_diffCommits_commitValid_90; \
        force U_IF_NAME.io_diffCommits_commitValid_91 = RTL_PATH.io_diffCommits_commitValid_91; \
        force U_IF_NAME.io_diffCommits_commitValid_92 = RTL_PATH.io_diffCommits_commitValid_92; \
        force U_IF_NAME.io_diffCommits_commitValid_93 = RTL_PATH.io_diffCommits_commitValid_93; \
        force U_IF_NAME.io_diffCommits_commitValid_94 = RTL_PATH.io_diffCommits_commitValid_94; \
        force U_IF_NAME.io_diffCommits_commitValid_95 = RTL_PATH.io_diffCommits_commitValid_95; \
        force U_IF_NAME.io_diffCommits_commitValid_96 = RTL_PATH.io_diffCommits_commitValid_96; \
        force U_IF_NAME.io_diffCommits_commitValid_97 = RTL_PATH.io_diffCommits_commitValid_97; \
        force U_IF_NAME.io_diffCommits_commitValid_98 = RTL_PATH.io_diffCommits_commitValid_98; \
        force U_IF_NAME.io_diffCommits_commitValid_99 = RTL_PATH.io_diffCommits_commitValid_99; \
        force U_IF_NAME.io_diffCommits_commitValid_100 = RTL_PATH.io_diffCommits_commitValid_100; \
        force U_IF_NAME.io_diffCommits_commitValid_101 = RTL_PATH.io_diffCommits_commitValid_101; \
        force U_IF_NAME.io_diffCommits_commitValid_102 = RTL_PATH.io_diffCommits_commitValid_102; \
        force U_IF_NAME.io_diffCommits_commitValid_103 = RTL_PATH.io_diffCommits_commitValid_103; \
        force U_IF_NAME.io_diffCommits_commitValid_104 = RTL_PATH.io_diffCommits_commitValid_104; \
        force U_IF_NAME.io_diffCommits_commitValid_105 = RTL_PATH.io_diffCommits_commitValid_105; \
        force U_IF_NAME.io_diffCommits_commitValid_106 = RTL_PATH.io_diffCommits_commitValid_106; \
        force U_IF_NAME.io_diffCommits_commitValid_107 = RTL_PATH.io_diffCommits_commitValid_107; \
        force U_IF_NAME.io_diffCommits_commitValid_108 = RTL_PATH.io_diffCommits_commitValid_108; \
        force U_IF_NAME.io_diffCommits_commitValid_109 = RTL_PATH.io_diffCommits_commitValid_109; \
        force U_IF_NAME.io_diffCommits_commitValid_110 = RTL_PATH.io_diffCommits_commitValid_110; \
        force U_IF_NAME.io_diffCommits_commitValid_111 = RTL_PATH.io_diffCommits_commitValid_111; \
        force U_IF_NAME.io_diffCommits_commitValid_112 = RTL_PATH.io_diffCommits_commitValid_112; \
        force U_IF_NAME.io_diffCommits_commitValid_113 = RTL_PATH.io_diffCommits_commitValid_113; \
        force U_IF_NAME.io_diffCommits_commitValid_114 = RTL_PATH.io_diffCommits_commitValid_114; \
        force U_IF_NAME.io_diffCommits_commitValid_115 = RTL_PATH.io_diffCommits_commitValid_115; \
        force U_IF_NAME.io_diffCommits_commitValid_116 = RTL_PATH.io_diffCommits_commitValid_116; \
        force U_IF_NAME.io_diffCommits_commitValid_117 = RTL_PATH.io_diffCommits_commitValid_117; \
        force U_IF_NAME.io_diffCommits_commitValid_118 = RTL_PATH.io_diffCommits_commitValid_118; \
        force U_IF_NAME.io_diffCommits_commitValid_119 = RTL_PATH.io_diffCommits_commitValid_119; \
        force U_IF_NAME.io_diffCommits_commitValid_120 = RTL_PATH.io_diffCommits_commitValid_120; \
        force U_IF_NAME.io_diffCommits_commitValid_121 = RTL_PATH.io_diffCommits_commitValid_121; \
        force U_IF_NAME.io_diffCommits_commitValid_122 = RTL_PATH.io_diffCommits_commitValid_122; \
        force U_IF_NAME.io_diffCommits_commitValid_123 = RTL_PATH.io_diffCommits_commitValid_123; \
        force U_IF_NAME.io_diffCommits_commitValid_124 = RTL_PATH.io_diffCommits_commitValid_124; \
        force U_IF_NAME.io_diffCommits_commitValid_125 = RTL_PATH.io_diffCommits_commitValid_125; \
        force U_IF_NAME.io_diffCommits_commitValid_126 = RTL_PATH.io_diffCommits_commitValid_126; \
        force U_IF_NAME.io_diffCommits_commitValid_127 = RTL_PATH.io_diffCommits_commitValid_127; \
        force U_IF_NAME.io_diffCommits_commitValid_128 = RTL_PATH.io_diffCommits_commitValid_128; \
        force U_IF_NAME.io_diffCommits_commitValid_129 = RTL_PATH.io_diffCommits_commitValid_129; \
        force U_IF_NAME.io_diffCommits_commitValid_130 = RTL_PATH.io_diffCommits_commitValid_130; \
        force U_IF_NAME.io_diffCommits_commitValid_131 = RTL_PATH.io_diffCommits_commitValid_131; \
        force U_IF_NAME.io_diffCommits_commitValid_132 = RTL_PATH.io_diffCommits_commitValid_132; \
        force U_IF_NAME.io_diffCommits_commitValid_133 = RTL_PATH.io_diffCommits_commitValid_133; \
        force U_IF_NAME.io_diffCommits_commitValid_134 = RTL_PATH.io_diffCommits_commitValid_134; \
        force U_IF_NAME.io_diffCommits_commitValid_135 = RTL_PATH.io_diffCommits_commitValid_135; \
        force U_IF_NAME.io_diffCommits_commitValid_136 = RTL_PATH.io_diffCommits_commitValid_136; \
        force U_IF_NAME.io_diffCommits_commitValid_137 = RTL_PATH.io_diffCommits_commitValid_137; \
        force U_IF_NAME.io_diffCommits_commitValid_138 = RTL_PATH.io_diffCommits_commitValid_138; \
        force U_IF_NAME.io_diffCommits_commitValid_139 = RTL_PATH.io_diffCommits_commitValid_139; \
        force U_IF_NAME.io_diffCommits_commitValid_140 = RTL_PATH.io_diffCommits_commitValid_140; \
        force U_IF_NAME.io_diffCommits_commitValid_141 = RTL_PATH.io_diffCommits_commitValid_141; \
        force U_IF_NAME.io_diffCommits_commitValid_142 = RTL_PATH.io_diffCommits_commitValid_142; \
        force U_IF_NAME.io_diffCommits_commitValid_143 = RTL_PATH.io_diffCommits_commitValid_143; \
        force U_IF_NAME.io_diffCommits_commitValid_144 = RTL_PATH.io_diffCommits_commitValid_144; \
        force U_IF_NAME.io_diffCommits_commitValid_145 = RTL_PATH.io_diffCommits_commitValid_145; \
        force U_IF_NAME.io_diffCommits_commitValid_146 = RTL_PATH.io_diffCommits_commitValid_146; \
        force U_IF_NAME.io_diffCommits_commitValid_147 = RTL_PATH.io_diffCommits_commitValid_147; \
        force U_IF_NAME.io_diffCommits_commitValid_148 = RTL_PATH.io_diffCommits_commitValid_148; \
        force U_IF_NAME.io_diffCommits_commitValid_149 = RTL_PATH.io_diffCommits_commitValid_149; \
        force U_IF_NAME.io_diffCommits_commitValid_150 = RTL_PATH.io_diffCommits_commitValid_150; \
        force U_IF_NAME.io_diffCommits_commitValid_151 = RTL_PATH.io_diffCommits_commitValid_151; \
        force U_IF_NAME.io_diffCommits_commitValid_152 = RTL_PATH.io_diffCommits_commitValid_152; \
        force U_IF_NAME.io_diffCommits_commitValid_153 = RTL_PATH.io_diffCommits_commitValid_153; \
        force U_IF_NAME.io_diffCommits_commitValid_154 = RTL_PATH.io_diffCommits_commitValid_154; \
        force U_IF_NAME.io_diffCommits_commitValid_155 = RTL_PATH.io_diffCommits_commitValid_155; \
        force U_IF_NAME.io_diffCommits_commitValid_156 = RTL_PATH.io_diffCommits_commitValid_156; \
        force U_IF_NAME.io_diffCommits_commitValid_157 = RTL_PATH.io_diffCommits_commitValid_157; \
        force U_IF_NAME.io_diffCommits_commitValid_158 = RTL_PATH.io_diffCommits_commitValid_158; \
        force U_IF_NAME.io_diffCommits_commitValid_159 = RTL_PATH.io_diffCommits_commitValid_159; \
        force U_IF_NAME.io_diffCommits_commitValid_160 = RTL_PATH.io_diffCommits_commitValid_160; \
        force U_IF_NAME.io_diffCommits_commitValid_161 = RTL_PATH.io_diffCommits_commitValid_161; \
        force U_IF_NAME.io_diffCommits_commitValid_162 = RTL_PATH.io_diffCommits_commitValid_162; \
        force U_IF_NAME.io_diffCommits_commitValid_163 = RTL_PATH.io_diffCommits_commitValid_163; \
        force U_IF_NAME.io_diffCommits_commitValid_164 = RTL_PATH.io_diffCommits_commitValid_164; \
        force U_IF_NAME.io_diffCommits_commitValid_165 = RTL_PATH.io_diffCommits_commitValid_165; \
        force U_IF_NAME.io_diffCommits_commitValid_166 = RTL_PATH.io_diffCommits_commitValid_166; \
        force U_IF_NAME.io_diffCommits_commitValid_167 = RTL_PATH.io_diffCommits_commitValid_167; \
        force U_IF_NAME.io_diffCommits_commitValid_168 = RTL_PATH.io_diffCommits_commitValid_168; \
        force U_IF_NAME.io_diffCommits_commitValid_169 = RTL_PATH.io_diffCommits_commitValid_169; \
        force U_IF_NAME.io_diffCommits_commitValid_170 = RTL_PATH.io_diffCommits_commitValid_170; \
        force U_IF_NAME.io_diffCommits_commitValid_171 = RTL_PATH.io_diffCommits_commitValid_171; \
        force U_IF_NAME.io_diffCommits_commitValid_172 = RTL_PATH.io_diffCommits_commitValid_172; \
        force U_IF_NAME.io_diffCommits_commitValid_173 = RTL_PATH.io_diffCommits_commitValid_173; \
        force U_IF_NAME.io_diffCommits_commitValid_174 = RTL_PATH.io_diffCommits_commitValid_174; \
        force U_IF_NAME.io_diffCommits_commitValid_175 = RTL_PATH.io_diffCommits_commitValid_175; \
        force U_IF_NAME.io_diffCommits_commitValid_176 = RTL_PATH.io_diffCommits_commitValid_176; \
        force U_IF_NAME.io_diffCommits_commitValid_177 = RTL_PATH.io_diffCommits_commitValid_177; \
        force U_IF_NAME.io_diffCommits_commitValid_178 = RTL_PATH.io_diffCommits_commitValid_178; \
        force U_IF_NAME.io_diffCommits_commitValid_179 = RTL_PATH.io_diffCommits_commitValid_179; \
        force U_IF_NAME.io_diffCommits_commitValid_180 = RTL_PATH.io_diffCommits_commitValid_180; \
        force U_IF_NAME.io_diffCommits_commitValid_181 = RTL_PATH.io_diffCommits_commitValid_181; \
        force U_IF_NAME.io_diffCommits_commitValid_182 = RTL_PATH.io_diffCommits_commitValid_182; \
        force U_IF_NAME.io_diffCommits_commitValid_183 = RTL_PATH.io_diffCommits_commitValid_183; \
        force U_IF_NAME.io_diffCommits_commitValid_184 = RTL_PATH.io_diffCommits_commitValid_184; \
        force U_IF_NAME.io_diffCommits_commitValid_185 = RTL_PATH.io_diffCommits_commitValid_185; \
        force U_IF_NAME.io_diffCommits_commitValid_186 = RTL_PATH.io_diffCommits_commitValid_186; \
        force U_IF_NAME.io_diffCommits_commitValid_187 = RTL_PATH.io_diffCommits_commitValid_187; \
        force U_IF_NAME.io_diffCommits_commitValid_188 = RTL_PATH.io_diffCommits_commitValid_188; \
        force U_IF_NAME.io_diffCommits_commitValid_189 = RTL_PATH.io_diffCommits_commitValid_189; \
        force U_IF_NAME.io_diffCommits_commitValid_190 = RTL_PATH.io_diffCommits_commitValid_190; \
        force U_IF_NAME.io_diffCommits_commitValid_191 = RTL_PATH.io_diffCommits_commitValid_191; \
        force U_IF_NAME.io_diffCommits_commitValid_192 = RTL_PATH.io_diffCommits_commitValid_192; \
        force U_IF_NAME.io_diffCommits_commitValid_193 = RTL_PATH.io_diffCommits_commitValid_193; \
        force U_IF_NAME.io_diffCommits_commitValid_194 = RTL_PATH.io_diffCommits_commitValid_194; \
        force U_IF_NAME.io_diffCommits_commitValid_195 = RTL_PATH.io_diffCommits_commitValid_195; \
        force U_IF_NAME.io_diffCommits_commitValid_196 = RTL_PATH.io_diffCommits_commitValid_196; \
        force U_IF_NAME.io_diffCommits_commitValid_197 = RTL_PATH.io_diffCommits_commitValid_197; \
        force U_IF_NAME.io_diffCommits_commitValid_198 = RTL_PATH.io_diffCommits_commitValid_198; \
        force U_IF_NAME.io_diffCommits_commitValid_199 = RTL_PATH.io_diffCommits_commitValid_199; \
        force U_IF_NAME.io_diffCommits_commitValid_200 = RTL_PATH.io_diffCommits_commitValid_200; \
        force U_IF_NAME.io_diffCommits_commitValid_201 = RTL_PATH.io_diffCommits_commitValid_201; \
        force U_IF_NAME.io_diffCommits_commitValid_202 = RTL_PATH.io_diffCommits_commitValid_202; \
        force U_IF_NAME.io_diffCommits_commitValid_203 = RTL_PATH.io_diffCommits_commitValid_203; \
        force U_IF_NAME.io_diffCommits_commitValid_204 = RTL_PATH.io_diffCommits_commitValid_204; \
        force U_IF_NAME.io_diffCommits_commitValid_205 = RTL_PATH.io_diffCommits_commitValid_205; \
        force U_IF_NAME.io_diffCommits_commitValid_206 = RTL_PATH.io_diffCommits_commitValid_206; \
        force U_IF_NAME.io_diffCommits_commitValid_207 = RTL_PATH.io_diffCommits_commitValid_207; \
        force U_IF_NAME.io_diffCommits_commitValid_208 = RTL_PATH.io_diffCommits_commitValid_208; \
        force U_IF_NAME.io_diffCommits_commitValid_209 = RTL_PATH.io_diffCommits_commitValid_209; \
        force U_IF_NAME.io_diffCommits_commitValid_210 = RTL_PATH.io_diffCommits_commitValid_210; \
        force U_IF_NAME.io_diffCommits_commitValid_211 = RTL_PATH.io_diffCommits_commitValid_211; \
        force U_IF_NAME.io_diffCommits_commitValid_212 = RTL_PATH.io_diffCommits_commitValid_212; \
        force U_IF_NAME.io_diffCommits_commitValid_213 = RTL_PATH.io_diffCommits_commitValid_213; \
        force U_IF_NAME.io_diffCommits_commitValid_214 = RTL_PATH.io_diffCommits_commitValid_214; \
        force U_IF_NAME.io_diffCommits_commitValid_215 = RTL_PATH.io_diffCommits_commitValid_215; \
        force U_IF_NAME.io_diffCommits_commitValid_216 = RTL_PATH.io_diffCommits_commitValid_216; \
        force U_IF_NAME.io_diffCommits_commitValid_217 = RTL_PATH.io_diffCommits_commitValid_217; \
        force U_IF_NAME.io_diffCommits_commitValid_218 = RTL_PATH.io_diffCommits_commitValid_218; \
        force U_IF_NAME.io_diffCommits_commitValid_219 = RTL_PATH.io_diffCommits_commitValid_219; \
        force U_IF_NAME.io_diffCommits_commitValid_220 = RTL_PATH.io_diffCommits_commitValid_220; \
        force U_IF_NAME.io_diffCommits_commitValid_221 = RTL_PATH.io_diffCommits_commitValid_221; \
        force U_IF_NAME.io_diffCommits_commitValid_222 = RTL_PATH.io_diffCommits_commitValid_222; \
        force U_IF_NAME.io_diffCommits_commitValid_223 = RTL_PATH.io_diffCommits_commitValid_223; \
        force U_IF_NAME.io_diffCommits_commitValid_224 = RTL_PATH.io_diffCommits_commitValid_224; \
        force U_IF_NAME.io_diffCommits_commitValid_225 = RTL_PATH.io_diffCommits_commitValid_225; \
        force U_IF_NAME.io_diffCommits_commitValid_226 = RTL_PATH.io_diffCommits_commitValid_226; \
        force U_IF_NAME.io_diffCommits_commitValid_227 = RTL_PATH.io_diffCommits_commitValid_227; \
        force U_IF_NAME.io_diffCommits_commitValid_228 = RTL_PATH.io_diffCommits_commitValid_228; \
        force U_IF_NAME.io_diffCommits_commitValid_229 = RTL_PATH.io_diffCommits_commitValid_229; \
        force U_IF_NAME.io_diffCommits_commitValid_230 = RTL_PATH.io_diffCommits_commitValid_230; \
        force U_IF_NAME.io_diffCommits_commitValid_231 = RTL_PATH.io_diffCommits_commitValid_231; \
        force U_IF_NAME.io_diffCommits_commitValid_232 = RTL_PATH.io_diffCommits_commitValid_232; \
        force U_IF_NAME.io_diffCommits_commitValid_233 = RTL_PATH.io_diffCommits_commitValid_233; \
        force U_IF_NAME.io_diffCommits_commitValid_234 = RTL_PATH.io_diffCommits_commitValid_234; \
        force U_IF_NAME.io_diffCommits_commitValid_235 = RTL_PATH.io_diffCommits_commitValid_235; \
        force U_IF_NAME.io_diffCommits_commitValid_236 = RTL_PATH.io_diffCommits_commitValid_236; \
        force U_IF_NAME.io_diffCommits_commitValid_237 = RTL_PATH.io_diffCommits_commitValid_237; \
        force U_IF_NAME.io_diffCommits_commitValid_238 = RTL_PATH.io_diffCommits_commitValid_238; \
        force U_IF_NAME.io_diffCommits_commitValid_239 = RTL_PATH.io_diffCommits_commitValid_239; \
        force U_IF_NAME.io_diffCommits_commitValid_240 = RTL_PATH.io_diffCommits_commitValid_240; \
        force U_IF_NAME.io_diffCommits_commitValid_241 = RTL_PATH.io_diffCommits_commitValid_241; \
        force U_IF_NAME.io_diffCommits_commitValid_242 = RTL_PATH.io_diffCommits_commitValid_242; \
        force U_IF_NAME.io_diffCommits_commitValid_243 = RTL_PATH.io_diffCommits_commitValid_243; \
        force U_IF_NAME.io_diffCommits_commitValid_244 = RTL_PATH.io_diffCommits_commitValid_244; \
        force U_IF_NAME.io_diffCommits_commitValid_245 = RTL_PATH.io_diffCommits_commitValid_245; \
        force U_IF_NAME.io_diffCommits_commitValid_246 = RTL_PATH.io_diffCommits_commitValid_246; \
        force U_IF_NAME.io_diffCommits_commitValid_247 = RTL_PATH.io_diffCommits_commitValid_247; \
        force U_IF_NAME.io_diffCommits_commitValid_248 = RTL_PATH.io_diffCommits_commitValid_248; \
        force U_IF_NAME.io_diffCommits_commitValid_249 = RTL_PATH.io_diffCommits_commitValid_249; \
        force U_IF_NAME.io_diffCommits_commitValid_250 = RTL_PATH.io_diffCommits_commitValid_250; \
        force U_IF_NAME.io_diffCommits_commitValid_251 = RTL_PATH.io_diffCommits_commitValid_251; \
        force U_IF_NAME.io_diffCommits_commitValid_252 = RTL_PATH.io_diffCommits_commitValid_252; \
        force U_IF_NAME.io_diffCommits_commitValid_253 = RTL_PATH.io_diffCommits_commitValid_253; \
        force U_IF_NAME.io_diffCommits_commitValid_254 = RTL_PATH.io_diffCommits_commitValid_254; \
        force U_IF_NAME.io_diffCommits_info_0_ldest = RTL_PATH.io_diffCommits_info_0_ldest; \
        force U_IF_NAME.io_diffCommits_info_0_pdest = RTL_PATH.io_diffCommits_info_0_pdest; \
        force U_IF_NAME.io_diffCommits_info_0_rfWen = RTL_PATH.io_diffCommits_info_0_rfWen; \
        force U_IF_NAME.io_diffCommits_info_0_fpWen = RTL_PATH.io_diffCommits_info_0_fpWen; \
        force U_IF_NAME.io_diffCommits_info_0_vecWen = RTL_PATH.io_diffCommits_info_0_vecWen; \
        force U_IF_NAME.io_diffCommits_info_0_v0Wen = RTL_PATH.io_diffCommits_info_0_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_0_vlWen = RTL_PATH.io_diffCommits_info_0_vlWen; \
        force U_IF_NAME.io_diffCommits_info_1_ldest = RTL_PATH.io_diffCommits_info_1_ldest; \
        force U_IF_NAME.io_diffCommits_info_1_pdest = RTL_PATH.io_diffCommits_info_1_pdest; \
        force U_IF_NAME.io_diffCommits_info_1_rfWen = RTL_PATH.io_diffCommits_info_1_rfWen; \
        force U_IF_NAME.io_diffCommits_info_1_fpWen = RTL_PATH.io_diffCommits_info_1_fpWen; \
        force U_IF_NAME.io_diffCommits_info_1_vecWen = RTL_PATH.io_diffCommits_info_1_vecWen; \
        force U_IF_NAME.io_diffCommits_info_1_v0Wen = RTL_PATH.io_diffCommits_info_1_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_1_vlWen = RTL_PATH.io_diffCommits_info_1_vlWen; \
        force U_IF_NAME.io_diffCommits_info_2_ldest = RTL_PATH.io_diffCommits_info_2_ldest; \
        force U_IF_NAME.io_diffCommits_info_2_pdest = RTL_PATH.io_diffCommits_info_2_pdest; \
        force U_IF_NAME.io_diffCommits_info_2_rfWen = RTL_PATH.io_diffCommits_info_2_rfWen; \
        force U_IF_NAME.io_diffCommits_info_2_fpWen = RTL_PATH.io_diffCommits_info_2_fpWen; \
        force U_IF_NAME.io_diffCommits_info_2_vecWen = RTL_PATH.io_diffCommits_info_2_vecWen; \
        force U_IF_NAME.io_diffCommits_info_2_v0Wen = RTL_PATH.io_diffCommits_info_2_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_2_vlWen = RTL_PATH.io_diffCommits_info_2_vlWen; \
        force U_IF_NAME.io_diffCommits_info_3_ldest = RTL_PATH.io_diffCommits_info_3_ldest; \
        force U_IF_NAME.io_diffCommits_info_3_pdest = RTL_PATH.io_diffCommits_info_3_pdest; \
        force U_IF_NAME.io_diffCommits_info_3_rfWen = RTL_PATH.io_diffCommits_info_3_rfWen; \
        force U_IF_NAME.io_diffCommits_info_3_fpWen = RTL_PATH.io_diffCommits_info_3_fpWen; \
        force U_IF_NAME.io_diffCommits_info_3_vecWen = RTL_PATH.io_diffCommits_info_3_vecWen; \
        force U_IF_NAME.io_diffCommits_info_3_v0Wen = RTL_PATH.io_diffCommits_info_3_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_3_vlWen = RTL_PATH.io_diffCommits_info_3_vlWen; \
        force U_IF_NAME.io_diffCommits_info_4_ldest = RTL_PATH.io_diffCommits_info_4_ldest; \
        force U_IF_NAME.io_diffCommits_info_4_pdest = RTL_PATH.io_diffCommits_info_4_pdest; \
        force U_IF_NAME.io_diffCommits_info_4_rfWen = RTL_PATH.io_diffCommits_info_4_rfWen; \
        force U_IF_NAME.io_diffCommits_info_4_fpWen = RTL_PATH.io_diffCommits_info_4_fpWen; \
        force U_IF_NAME.io_diffCommits_info_4_vecWen = RTL_PATH.io_diffCommits_info_4_vecWen; \
        force U_IF_NAME.io_diffCommits_info_4_v0Wen = RTL_PATH.io_diffCommits_info_4_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_4_vlWen = RTL_PATH.io_diffCommits_info_4_vlWen; \
        force U_IF_NAME.io_diffCommits_info_5_ldest = RTL_PATH.io_diffCommits_info_5_ldest; \
        force U_IF_NAME.io_diffCommits_info_5_pdest = RTL_PATH.io_diffCommits_info_5_pdest; \
        force U_IF_NAME.io_diffCommits_info_5_rfWen = RTL_PATH.io_diffCommits_info_5_rfWen; \
        force U_IF_NAME.io_diffCommits_info_5_fpWen = RTL_PATH.io_diffCommits_info_5_fpWen; \
        force U_IF_NAME.io_diffCommits_info_5_vecWen = RTL_PATH.io_diffCommits_info_5_vecWen; \
        force U_IF_NAME.io_diffCommits_info_5_v0Wen = RTL_PATH.io_diffCommits_info_5_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_5_vlWen = RTL_PATH.io_diffCommits_info_5_vlWen; \
        force U_IF_NAME.io_diffCommits_info_6_ldest = RTL_PATH.io_diffCommits_info_6_ldest; \
        force U_IF_NAME.io_diffCommits_info_6_pdest = RTL_PATH.io_diffCommits_info_6_pdest; \
        force U_IF_NAME.io_diffCommits_info_6_rfWen = RTL_PATH.io_diffCommits_info_6_rfWen; \
        force U_IF_NAME.io_diffCommits_info_6_fpWen = RTL_PATH.io_diffCommits_info_6_fpWen; \
        force U_IF_NAME.io_diffCommits_info_6_vecWen = RTL_PATH.io_diffCommits_info_6_vecWen; \
        force U_IF_NAME.io_diffCommits_info_6_v0Wen = RTL_PATH.io_diffCommits_info_6_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_6_vlWen = RTL_PATH.io_diffCommits_info_6_vlWen; \
        force U_IF_NAME.io_diffCommits_info_7_ldest = RTL_PATH.io_diffCommits_info_7_ldest; \
        force U_IF_NAME.io_diffCommits_info_7_pdest = RTL_PATH.io_diffCommits_info_7_pdest; \
        force U_IF_NAME.io_diffCommits_info_7_rfWen = RTL_PATH.io_diffCommits_info_7_rfWen; \
        force U_IF_NAME.io_diffCommits_info_7_fpWen = RTL_PATH.io_diffCommits_info_7_fpWen; \
        force U_IF_NAME.io_diffCommits_info_7_vecWen = RTL_PATH.io_diffCommits_info_7_vecWen; \
        force U_IF_NAME.io_diffCommits_info_7_v0Wen = RTL_PATH.io_diffCommits_info_7_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_7_vlWen = RTL_PATH.io_diffCommits_info_7_vlWen; \
        force U_IF_NAME.io_diffCommits_info_8_ldest = RTL_PATH.io_diffCommits_info_8_ldest; \
        force U_IF_NAME.io_diffCommits_info_8_pdest = RTL_PATH.io_diffCommits_info_8_pdest; \
        force U_IF_NAME.io_diffCommits_info_8_rfWen = RTL_PATH.io_diffCommits_info_8_rfWen; \
        force U_IF_NAME.io_diffCommits_info_8_fpWen = RTL_PATH.io_diffCommits_info_8_fpWen; \
        force U_IF_NAME.io_diffCommits_info_8_vecWen = RTL_PATH.io_diffCommits_info_8_vecWen; \
        force U_IF_NAME.io_diffCommits_info_8_v0Wen = RTL_PATH.io_diffCommits_info_8_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_8_vlWen = RTL_PATH.io_diffCommits_info_8_vlWen; \
        force U_IF_NAME.io_diffCommits_info_9_ldest = RTL_PATH.io_diffCommits_info_9_ldest; \
        force U_IF_NAME.io_diffCommits_info_9_pdest = RTL_PATH.io_diffCommits_info_9_pdest; \
        force U_IF_NAME.io_diffCommits_info_9_rfWen = RTL_PATH.io_diffCommits_info_9_rfWen; \
        force U_IF_NAME.io_diffCommits_info_9_fpWen = RTL_PATH.io_diffCommits_info_9_fpWen; \
        force U_IF_NAME.io_diffCommits_info_9_vecWen = RTL_PATH.io_diffCommits_info_9_vecWen; \
        force U_IF_NAME.io_diffCommits_info_9_v0Wen = RTL_PATH.io_diffCommits_info_9_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_9_vlWen = RTL_PATH.io_diffCommits_info_9_vlWen; \
        force U_IF_NAME.io_diffCommits_info_10_ldest = RTL_PATH.io_diffCommits_info_10_ldest; \
        force U_IF_NAME.io_diffCommits_info_10_pdest = RTL_PATH.io_diffCommits_info_10_pdest; \
        force U_IF_NAME.io_diffCommits_info_10_rfWen = RTL_PATH.io_diffCommits_info_10_rfWen; \
        force U_IF_NAME.io_diffCommits_info_10_fpWen = RTL_PATH.io_diffCommits_info_10_fpWen; \
        force U_IF_NAME.io_diffCommits_info_10_vecWen = RTL_PATH.io_diffCommits_info_10_vecWen; \
        force U_IF_NAME.io_diffCommits_info_10_v0Wen = RTL_PATH.io_diffCommits_info_10_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_10_vlWen = RTL_PATH.io_diffCommits_info_10_vlWen; \
        force U_IF_NAME.io_diffCommits_info_11_ldest = RTL_PATH.io_diffCommits_info_11_ldest; \
        force U_IF_NAME.io_diffCommits_info_11_pdest = RTL_PATH.io_diffCommits_info_11_pdest; \
        force U_IF_NAME.io_diffCommits_info_11_rfWen = RTL_PATH.io_diffCommits_info_11_rfWen; \
        force U_IF_NAME.io_diffCommits_info_11_fpWen = RTL_PATH.io_diffCommits_info_11_fpWen; \
        force U_IF_NAME.io_diffCommits_info_11_vecWen = RTL_PATH.io_diffCommits_info_11_vecWen; \
        force U_IF_NAME.io_diffCommits_info_11_v0Wen = RTL_PATH.io_diffCommits_info_11_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_11_vlWen = RTL_PATH.io_diffCommits_info_11_vlWen; \
        force U_IF_NAME.io_diffCommits_info_12_ldest = RTL_PATH.io_diffCommits_info_12_ldest; \
        force U_IF_NAME.io_diffCommits_info_12_pdest = RTL_PATH.io_diffCommits_info_12_pdest; \
        force U_IF_NAME.io_diffCommits_info_12_rfWen = RTL_PATH.io_diffCommits_info_12_rfWen; \
        force U_IF_NAME.io_diffCommits_info_12_fpWen = RTL_PATH.io_diffCommits_info_12_fpWen; \
        force U_IF_NAME.io_diffCommits_info_12_vecWen = RTL_PATH.io_diffCommits_info_12_vecWen; \
        force U_IF_NAME.io_diffCommits_info_12_v0Wen = RTL_PATH.io_diffCommits_info_12_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_12_vlWen = RTL_PATH.io_diffCommits_info_12_vlWen; \
        force U_IF_NAME.io_diffCommits_info_13_ldest = RTL_PATH.io_diffCommits_info_13_ldest; \
        force U_IF_NAME.io_diffCommits_info_13_pdest = RTL_PATH.io_diffCommits_info_13_pdest; \
        force U_IF_NAME.io_diffCommits_info_13_rfWen = RTL_PATH.io_diffCommits_info_13_rfWen; \
        force U_IF_NAME.io_diffCommits_info_13_fpWen = RTL_PATH.io_diffCommits_info_13_fpWen; \
        force U_IF_NAME.io_diffCommits_info_13_vecWen = RTL_PATH.io_diffCommits_info_13_vecWen; \
        force U_IF_NAME.io_diffCommits_info_13_v0Wen = RTL_PATH.io_diffCommits_info_13_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_13_vlWen = RTL_PATH.io_diffCommits_info_13_vlWen; \
        force U_IF_NAME.io_diffCommits_info_14_ldest = RTL_PATH.io_diffCommits_info_14_ldest; \
        force U_IF_NAME.io_diffCommits_info_14_pdest = RTL_PATH.io_diffCommits_info_14_pdest; \
        force U_IF_NAME.io_diffCommits_info_14_rfWen = RTL_PATH.io_diffCommits_info_14_rfWen; \
        force U_IF_NAME.io_diffCommits_info_14_fpWen = RTL_PATH.io_diffCommits_info_14_fpWen; \
        force U_IF_NAME.io_diffCommits_info_14_vecWen = RTL_PATH.io_diffCommits_info_14_vecWen; \
        force U_IF_NAME.io_diffCommits_info_14_v0Wen = RTL_PATH.io_diffCommits_info_14_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_14_vlWen = RTL_PATH.io_diffCommits_info_14_vlWen; \
        force U_IF_NAME.io_diffCommits_info_15_ldest = RTL_PATH.io_diffCommits_info_15_ldest; \
        force U_IF_NAME.io_diffCommits_info_15_pdest = RTL_PATH.io_diffCommits_info_15_pdest; \
        force U_IF_NAME.io_diffCommits_info_15_rfWen = RTL_PATH.io_diffCommits_info_15_rfWen; \
        force U_IF_NAME.io_diffCommits_info_15_fpWen = RTL_PATH.io_diffCommits_info_15_fpWen; \
        force U_IF_NAME.io_diffCommits_info_15_vecWen = RTL_PATH.io_diffCommits_info_15_vecWen; \
        force U_IF_NAME.io_diffCommits_info_15_v0Wen = RTL_PATH.io_diffCommits_info_15_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_15_vlWen = RTL_PATH.io_diffCommits_info_15_vlWen; \
        force U_IF_NAME.io_diffCommits_info_16_ldest = RTL_PATH.io_diffCommits_info_16_ldest; \
        force U_IF_NAME.io_diffCommits_info_16_pdest = RTL_PATH.io_diffCommits_info_16_pdest; \
        force U_IF_NAME.io_diffCommits_info_16_rfWen = RTL_PATH.io_diffCommits_info_16_rfWen; \
        force U_IF_NAME.io_diffCommits_info_16_fpWen = RTL_PATH.io_diffCommits_info_16_fpWen; \
        force U_IF_NAME.io_diffCommits_info_16_vecWen = RTL_PATH.io_diffCommits_info_16_vecWen; \
        force U_IF_NAME.io_diffCommits_info_16_v0Wen = RTL_PATH.io_diffCommits_info_16_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_16_vlWen = RTL_PATH.io_diffCommits_info_16_vlWen; \
        force U_IF_NAME.io_diffCommits_info_17_ldest = RTL_PATH.io_diffCommits_info_17_ldest; \
        force U_IF_NAME.io_diffCommits_info_17_pdest = RTL_PATH.io_diffCommits_info_17_pdest; \
        force U_IF_NAME.io_diffCommits_info_17_rfWen = RTL_PATH.io_diffCommits_info_17_rfWen; \
        force U_IF_NAME.io_diffCommits_info_17_fpWen = RTL_PATH.io_diffCommits_info_17_fpWen; \
        force U_IF_NAME.io_diffCommits_info_17_vecWen = RTL_PATH.io_diffCommits_info_17_vecWen; \
        force U_IF_NAME.io_diffCommits_info_17_v0Wen = RTL_PATH.io_diffCommits_info_17_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_17_vlWen = RTL_PATH.io_diffCommits_info_17_vlWen; \
        force U_IF_NAME.io_diffCommits_info_18_ldest = RTL_PATH.io_diffCommits_info_18_ldest; \
        force U_IF_NAME.io_diffCommits_info_18_pdest = RTL_PATH.io_diffCommits_info_18_pdest; \
        force U_IF_NAME.io_diffCommits_info_18_rfWen = RTL_PATH.io_diffCommits_info_18_rfWen; \
        force U_IF_NAME.io_diffCommits_info_18_fpWen = RTL_PATH.io_diffCommits_info_18_fpWen; \
        force U_IF_NAME.io_diffCommits_info_18_vecWen = RTL_PATH.io_diffCommits_info_18_vecWen; \
        force U_IF_NAME.io_diffCommits_info_18_v0Wen = RTL_PATH.io_diffCommits_info_18_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_18_vlWen = RTL_PATH.io_diffCommits_info_18_vlWen; \
        force U_IF_NAME.io_diffCommits_info_19_ldest = RTL_PATH.io_diffCommits_info_19_ldest; \
        force U_IF_NAME.io_diffCommits_info_19_pdest = RTL_PATH.io_diffCommits_info_19_pdest; \
        force U_IF_NAME.io_diffCommits_info_19_rfWen = RTL_PATH.io_diffCommits_info_19_rfWen; \
        force U_IF_NAME.io_diffCommits_info_19_fpWen = RTL_PATH.io_diffCommits_info_19_fpWen; \
        force U_IF_NAME.io_diffCommits_info_19_vecWen = RTL_PATH.io_diffCommits_info_19_vecWen; \
        force U_IF_NAME.io_diffCommits_info_19_v0Wen = RTL_PATH.io_diffCommits_info_19_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_19_vlWen = RTL_PATH.io_diffCommits_info_19_vlWen; \
        force U_IF_NAME.io_diffCommits_info_20_ldest = RTL_PATH.io_diffCommits_info_20_ldest; \
        force U_IF_NAME.io_diffCommits_info_20_pdest = RTL_PATH.io_diffCommits_info_20_pdest; \
        force U_IF_NAME.io_diffCommits_info_20_rfWen = RTL_PATH.io_diffCommits_info_20_rfWen; \
        force U_IF_NAME.io_diffCommits_info_20_fpWen = RTL_PATH.io_diffCommits_info_20_fpWen; \
        force U_IF_NAME.io_diffCommits_info_20_vecWen = RTL_PATH.io_diffCommits_info_20_vecWen; \
        force U_IF_NAME.io_diffCommits_info_20_v0Wen = RTL_PATH.io_diffCommits_info_20_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_20_vlWen = RTL_PATH.io_diffCommits_info_20_vlWen; \
        force U_IF_NAME.io_diffCommits_info_21_ldest = RTL_PATH.io_diffCommits_info_21_ldest; \
        force U_IF_NAME.io_diffCommits_info_21_pdest = RTL_PATH.io_diffCommits_info_21_pdest; \
        force U_IF_NAME.io_diffCommits_info_21_rfWen = RTL_PATH.io_diffCommits_info_21_rfWen; \
        force U_IF_NAME.io_diffCommits_info_21_fpWen = RTL_PATH.io_diffCommits_info_21_fpWen; \
        force U_IF_NAME.io_diffCommits_info_21_vecWen = RTL_PATH.io_diffCommits_info_21_vecWen; \
        force U_IF_NAME.io_diffCommits_info_21_v0Wen = RTL_PATH.io_diffCommits_info_21_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_21_vlWen = RTL_PATH.io_diffCommits_info_21_vlWen; \
        force U_IF_NAME.io_diffCommits_info_22_ldest = RTL_PATH.io_diffCommits_info_22_ldest; \
        force U_IF_NAME.io_diffCommits_info_22_pdest = RTL_PATH.io_diffCommits_info_22_pdest; \
        force U_IF_NAME.io_diffCommits_info_22_rfWen = RTL_PATH.io_diffCommits_info_22_rfWen; \
        force U_IF_NAME.io_diffCommits_info_22_fpWen = RTL_PATH.io_diffCommits_info_22_fpWen; \
        force U_IF_NAME.io_diffCommits_info_22_vecWen = RTL_PATH.io_diffCommits_info_22_vecWen; \
        force U_IF_NAME.io_diffCommits_info_22_v0Wen = RTL_PATH.io_diffCommits_info_22_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_22_vlWen = RTL_PATH.io_diffCommits_info_22_vlWen; \
        force U_IF_NAME.io_diffCommits_info_23_ldest = RTL_PATH.io_diffCommits_info_23_ldest; \
        force U_IF_NAME.io_diffCommits_info_23_pdest = RTL_PATH.io_diffCommits_info_23_pdest; \
        force U_IF_NAME.io_diffCommits_info_23_rfWen = RTL_PATH.io_diffCommits_info_23_rfWen; \
        force U_IF_NAME.io_diffCommits_info_23_fpWen = RTL_PATH.io_diffCommits_info_23_fpWen; \
        force U_IF_NAME.io_diffCommits_info_23_vecWen = RTL_PATH.io_diffCommits_info_23_vecWen; \
        force U_IF_NAME.io_diffCommits_info_23_v0Wen = RTL_PATH.io_diffCommits_info_23_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_23_vlWen = RTL_PATH.io_diffCommits_info_23_vlWen; \
        force U_IF_NAME.io_diffCommits_info_24_ldest = RTL_PATH.io_diffCommits_info_24_ldest; \
        force U_IF_NAME.io_diffCommits_info_24_pdest = RTL_PATH.io_diffCommits_info_24_pdest; \
        force U_IF_NAME.io_diffCommits_info_24_rfWen = RTL_PATH.io_diffCommits_info_24_rfWen; \
        force U_IF_NAME.io_diffCommits_info_24_fpWen = RTL_PATH.io_diffCommits_info_24_fpWen; \
        force U_IF_NAME.io_diffCommits_info_24_vecWen = RTL_PATH.io_diffCommits_info_24_vecWen; \
        force U_IF_NAME.io_diffCommits_info_24_v0Wen = RTL_PATH.io_diffCommits_info_24_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_24_vlWen = RTL_PATH.io_diffCommits_info_24_vlWen; \
        force U_IF_NAME.io_diffCommits_info_25_ldest = RTL_PATH.io_diffCommits_info_25_ldest; \
        force U_IF_NAME.io_diffCommits_info_25_pdest = RTL_PATH.io_diffCommits_info_25_pdest; \
        force U_IF_NAME.io_diffCommits_info_25_rfWen = RTL_PATH.io_diffCommits_info_25_rfWen; \
        force U_IF_NAME.io_diffCommits_info_25_fpWen = RTL_PATH.io_diffCommits_info_25_fpWen; \
        force U_IF_NAME.io_diffCommits_info_25_vecWen = RTL_PATH.io_diffCommits_info_25_vecWen; \
        force U_IF_NAME.io_diffCommits_info_25_v0Wen = RTL_PATH.io_diffCommits_info_25_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_25_vlWen = RTL_PATH.io_diffCommits_info_25_vlWen; \
        force U_IF_NAME.io_diffCommits_info_26_ldest = RTL_PATH.io_diffCommits_info_26_ldest; \
        force U_IF_NAME.io_diffCommits_info_26_pdest = RTL_PATH.io_diffCommits_info_26_pdest; \
        force U_IF_NAME.io_diffCommits_info_26_rfWen = RTL_PATH.io_diffCommits_info_26_rfWen; \
        force U_IF_NAME.io_diffCommits_info_26_fpWen = RTL_PATH.io_diffCommits_info_26_fpWen; \
        force U_IF_NAME.io_diffCommits_info_26_vecWen = RTL_PATH.io_diffCommits_info_26_vecWen; \
        force U_IF_NAME.io_diffCommits_info_26_v0Wen = RTL_PATH.io_diffCommits_info_26_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_26_vlWen = RTL_PATH.io_diffCommits_info_26_vlWen; \
        force U_IF_NAME.io_diffCommits_info_27_ldest = RTL_PATH.io_diffCommits_info_27_ldest; \
        force U_IF_NAME.io_diffCommits_info_27_pdest = RTL_PATH.io_diffCommits_info_27_pdest; \
        force U_IF_NAME.io_diffCommits_info_27_rfWen = RTL_PATH.io_diffCommits_info_27_rfWen; \
        force U_IF_NAME.io_diffCommits_info_27_fpWen = RTL_PATH.io_diffCommits_info_27_fpWen; \
        force U_IF_NAME.io_diffCommits_info_27_vecWen = RTL_PATH.io_diffCommits_info_27_vecWen; \
        force U_IF_NAME.io_diffCommits_info_27_v0Wen = RTL_PATH.io_diffCommits_info_27_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_27_vlWen = RTL_PATH.io_diffCommits_info_27_vlWen; \
        force U_IF_NAME.io_diffCommits_info_28_ldest = RTL_PATH.io_diffCommits_info_28_ldest; \
        force U_IF_NAME.io_diffCommits_info_28_pdest = RTL_PATH.io_diffCommits_info_28_pdest; \
        force U_IF_NAME.io_diffCommits_info_28_rfWen = RTL_PATH.io_diffCommits_info_28_rfWen; \
        force U_IF_NAME.io_diffCommits_info_28_fpWen = RTL_PATH.io_diffCommits_info_28_fpWen; \
        force U_IF_NAME.io_diffCommits_info_28_vecWen = RTL_PATH.io_diffCommits_info_28_vecWen; \
        force U_IF_NAME.io_diffCommits_info_28_v0Wen = RTL_PATH.io_diffCommits_info_28_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_28_vlWen = RTL_PATH.io_diffCommits_info_28_vlWen; \
        force U_IF_NAME.io_diffCommits_info_29_ldest = RTL_PATH.io_diffCommits_info_29_ldest; \
        force U_IF_NAME.io_diffCommits_info_29_pdest = RTL_PATH.io_diffCommits_info_29_pdest; \
        force U_IF_NAME.io_diffCommits_info_29_rfWen = RTL_PATH.io_diffCommits_info_29_rfWen; \
        force U_IF_NAME.io_diffCommits_info_29_fpWen = RTL_PATH.io_diffCommits_info_29_fpWen; \
        force U_IF_NAME.io_diffCommits_info_29_vecWen = RTL_PATH.io_diffCommits_info_29_vecWen; \
        force U_IF_NAME.io_diffCommits_info_29_v0Wen = RTL_PATH.io_diffCommits_info_29_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_29_vlWen = RTL_PATH.io_diffCommits_info_29_vlWen; \
        force U_IF_NAME.io_diffCommits_info_30_ldest = RTL_PATH.io_diffCommits_info_30_ldest; \
        force U_IF_NAME.io_diffCommits_info_30_pdest = RTL_PATH.io_diffCommits_info_30_pdest; \
        force U_IF_NAME.io_diffCommits_info_30_rfWen = RTL_PATH.io_diffCommits_info_30_rfWen; \
        force U_IF_NAME.io_diffCommits_info_30_fpWen = RTL_PATH.io_diffCommits_info_30_fpWen; \
        force U_IF_NAME.io_diffCommits_info_30_vecWen = RTL_PATH.io_diffCommits_info_30_vecWen; \
        force U_IF_NAME.io_diffCommits_info_30_v0Wen = RTL_PATH.io_diffCommits_info_30_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_30_vlWen = RTL_PATH.io_diffCommits_info_30_vlWen; \
        force U_IF_NAME.io_diffCommits_info_31_ldest = RTL_PATH.io_diffCommits_info_31_ldest; \
        force U_IF_NAME.io_diffCommits_info_31_pdest = RTL_PATH.io_diffCommits_info_31_pdest; \
        force U_IF_NAME.io_diffCommits_info_31_rfWen = RTL_PATH.io_diffCommits_info_31_rfWen; \
        force U_IF_NAME.io_diffCommits_info_31_fpWen = RTL_PATH.io_diffCommits_info_31_fpWen; \
        force U_IF_NAME.io_diffCommits_info_31_vecWen = RTL_PATH.io_diffCommits_info_31_vecWen; \
        force U_IF_NAME.io_diffCommits_info_31_v0Wen = RTL_PATH.io_diffCommits_info_31_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_31_vlWen = RTL_PATH.io_diffCommits_info_31_vlWen; \
        force U_IF_NAME.io_diffCommits_info_32_ldest = RTL_PATH.io_diffCommits_info_32_ldest; \
        force U_IF_NAME.io_diffCommits_info_32_pdest = RTL_PATH.io_diffCommits_info_32_pdest; \
        force U_IF_NAME.io_diffCommits_info_32_rfWen = RTL_PATH.io_diffCommits_info_32_rfWen; \
        force U_IF_NAME.io_diffCommits_info_32_fpWen = RTL_PATH.io_diffCommits_info_32_fpWen; \
        force U_IF_NAME.io_diffCommits_info_32_vecWen = RTL_PATH.io_diffCommits_info_32_vecWen; \
        force U_IF_NAME.io_diffCommits_info_32_v0Wen = RTL_PATH.io_diffCommits_info_32_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_32_vlWen = RTL_PATH.io_diffCommits_info_32_vlWen; \
        force U_IF_NAME.io_diffCommits_info_33_ldest = RTL_PATH.io_diffCommits_info_33_ldest; \
        force U_IF_NAME.io_diffCommits_info_33_pdest = RTL_PATH.io_diffCommits_info_33_pdest; \
        force U_IF_NAME.io_diffCommits_info_33_rfWen = RTL_PATH.io_diffCommits_info_33_rfWen; \
        force U_IF_NAME.io_diffCommits_info_33_fpWen = RTL_PATH.io_diffCommits_info_33_fpWen; \
        force U_IF_NAME.io_diffCommits_info_33_vecWen = RTL_PATH.io_diffCommits_info_33_vecWen; \
        force U_IF_NAME.io_diffCommits_info_33_v0Wen = RTL_PATH.io_diffCommits_info_33_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_33_vlWen = RTL_PATH.io_diffCommits_info_33_vlWen; \
        force U_IF_NAME.io_diffCommits_info_34_ldest = RTL_PATH.io_diffCommits_info_34_ldest; \
        force U_IF_NAME.io_diffCommits_info_34_pdest = RTL_PATH.io_diffCommits_info_34_pdest; \
        force U_IF_NAME.io_diffCommits_info_34_rfWen = RTL_PATH.io_diffCommits_info_34_rfWen; \
        force U_IF_NAME.io_diffCommits_info_34_fpWen = RTL_PATH.io_diffCommits_info_34_fpWen; \
        force U_IF_NAME.io_diffCommits_info_34_vecWen = RTL_PATH.io_diffCommits_info_34_vecWen; \
        force U_IF_NAME.io_diffCommits_info_34_v0Wen = RTL_PATH.io_diffCommits_info_34_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_34_vlWen = RTL_PATH.io_diffCommits_info_34_vlWen; \
        force U_IF_NAME.io_diffCommits_info_35_ldest = RTL_PATH.io_diffCommits_info_35_ldest; \
        force U_IF_NAME.io_diffCommits_info_35_pdest = RTL_PATH.io_diffCommits_info_35_pdest; \
        force U_IF_NAME.io_diffCommits_info_35_rfWen = RTL_PATH.io_diffCommits_info_35_rfWen; \
        force U_IF_NAME.io_diffCommits_info_35_fpWen = RTL_PATH.io_diffCommits_info_35_fpWen; \
        force U_IF_NAME.io_diffCommits_info_35_vecWen = RTL_PATH.io_diffCommits_info_35_vecWen; \
        force U_IF_NAME.io_diffCommits_info_35_v0Wen = RTL_PATH.io_diffCommits_info_35_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_35_vlWen = RTL_PATH.io_diffCommits_info_35_vlWen; \
        force U_IF_NAME.io_diffCommits_info_36_ldest = RTL_PATH.io_diffCommits_info_36_ldest; \
        force U_IF_NAME.io_diffCommits_info_36_pdest = RTL_PATH.io_diffCommits_info_36_pdest; \
        force U_IF_NAME.io_diffCommits_info_36_rfWen = RTL_PATH.io_diffCommits_info_36_rfWen; \
        force U_IF_NAME.io_diffCommits_info_36_fpWen = RTL_PATH.io_diffCommits_info_36_fpWen; \
        force U_IF_NAME.io_diffCommits_info_36_vecWen = RTL_PATH.io_diffCommits_info_36_vecWen; \
        force U_IF_NAME.io_diffCommits_info_36_v0Wen = RTL_PATH.io_diffCommits_info_36_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_36_vlWen = RTL_PATH.io_diffCommits_info_36_vlWen; \
        force U_IF_NAME.io_diffCommits_info_37_ldest = RTL_PATH.io_diffCommits_info_37_ldest; \
        force U_IF_NAME.io_diffCommits_info_37_pdest = RTL_PATH.io_diffCommits_info_37_pdest; \
        force U_IF_NAME.io_diffCommits_info_37_rfWen = RTL_PATH.io_diffCommits_info_37_rfWen; \
        force U_IF_NAME.io_diffCommits_info_37_fpWen = RTL_PATH.io_diffCommits_info_37_fpWen; \
        force U_IF_NAME.io_diffCommits_info_37_vecWen = RTL_PATH.io_diffCommits_info_37_vecWen; \
        force U_IF_NAME.io_diffCommits_info_37_v0Wen = RTL_PATH.io_diffCommits_info_37_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_37_vlWen = RTL_PATH.io_diffCommits_info_37_vlWen; \
        force U_IF_NAME.io_diffCommits_info_38_ldest = RTL_PATH.io_diffCommits_info_38_ldest; \
        force U_IF_NAME.io_diffCommits_info_38_pdest = RTL_PATH.io_diffCommits_info_38_pdest; \
        force U_IF_NAME.io_diffCommits_info_38_rfWen = RTL_PATH.io_diffCommits_info_38_rfWen; \
        force U_IF_NAME.io_diffCommits_info_38_fpWen = RTL_PATH.io_diffCommits_info_38_fpWen; \
        force U_IF_NAME.io_diffCommits_info_38_vecWen = RTL_PATH.io_diffCommits_info_38_vecWen; \
        force U_IF_NAME.io_diffCommits_info_38_v0Wen = RTL_PATH.io_diffCommits_info_38_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_38_vlWen = RTL_PATH.io_diffCommits_info_38_vlWen; \
        force U_IF_NAME.io_diffCommits_info_39_ldest = RTL_PATH.io_diffCommits_info_39_ldest; \
        force U_IF_NAME.io_diffCommits_info_39_pdest = RTL_PATH.io_diffCommits_info_39_pdest; \
        force U_IF_NAME.io_diffCommits_info_39_rfWen = RTL_PATH.io_diffCommits_info_39_rfWen; \
        force U_IF_NAME.io_diffCommits_info_39_fpWen = RTL_PATH.io_diffCommits_info_39_fpWen; \
        force U_IF_NAME.io_diffCommits_info_39_vecWen = RTL_PATH.io_diffCommits_info_39_vecWen; \
        force U_IF_NAME.io_diffCommits_info_39_v0Wen = RTL_PATH.io_diffCommits_info_39_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_39_vlWen = RTL_PATH.io_diffCommits_info_39_vlWen; \
        force U_IF_NAME.io_diffCommits_info_40_ldest = RTL_PATH.io_diffCommits_info_40_ldest; \
        force U_IF_NAME.io_diffCommits_info_40_pdest = RTL_PATH.io_diffCommits_info_40_pdest; \
        force U_IF_NAME.io_diffCommits_info_40_rfWen = RTL_PATH.io_diffCommits_info_40_rfWen; \
        force U_IF_NAME.io_diffCommits_info_40_fpWen = RTL_PATH.io_diffCommits_info_40_fpWen; \
        force U_IF_NAME.io_diffCommits_info_40_vecWen = RTL_PATH.io_diffCommits_info_40_vecWen; \
        force U_IF_NAME.io_diffCommits_info_40_v0Wen = RTL_PATH.io_diffCommits_info_40_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_40_vlWen = RTL_PATH.io_diffCommits_info_40_vlWen; \
        force U_IF_NAME.io_diffCommits_info_41_ldest = RTL_PATH.io_diffCommits_info_41_ldest; \
        force U_IF_NAME.io_diffCommits_info_41_pdest = RTL_PATH.io_diffCommits_info_41_pdest; \
        force U_IF_NAME.io_diffCommits_info_41_rfWen = RTL_PATH.io_diffCommits_info_41_rfWen; \
        force U_IF_NAME.io_diffCommits_info_41_fpWen = RTL_PATH.io_diffCommits_info_41_fpWen; \
        force U_IF_NAME.io_diffCommits_info_41_vecWen = RTL_PATH.io_diffCommits_info_41_vecWen; \
        force U_IF_NAME.io_diffCommits_info_41_v0Wen = RTL_PATH.io_diffCommits_info_41_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_41_vlWen = RTL_PATH.io_diffCommits_info_41_vlWen; \
        force U_IF_NAME.io_diffCommits_info_42_ldest = RTL_PATH.io_diffCommits_info_42_ldest; \
        force U_IF_NAME.io_diffCommits_info_42_pdest = RTL_PATH.io_diffCommits_info_42_pdest; \
        force U_IF_NAME.io_diffCommits_info_42_rfWen = RTL_PATH.io_diffCommits_info_42_rfWen; \
        force U_IF_NAME.io_diffCommits_info_42_fpWen = RTL_PATH.io_diffCommits_info_42_fpWen; \
        force U_IF_NAME.io_diffCommits_info_42_vecWen = RTL_PATH.io_diffCommits_info_42_vecWen; \
        force U_IF_NAME.io_diffCommits_info_42_v0Wen = RTL_PATH.io_diffCommits_info_42_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_42_vlWen = RTL_PATH.io_diffCommits_info_42_vlWen; \
        force U_IF_NAME.io_diffCommits_info_43_ldest = RTL_PATH.io_diffCommits_info_43_ldest; \
        force U_IF_NAME.io_diffCommits_info_43_pdest = RTL_PATH.io_diffCommits_info_43_pdest; \
        force U_IF_NAME.io_diffCommits_info_43_rfWen = RTL_PATH.io_diffCommits_info_43_rfWen; \
        force U_IF_NAME.io_diffCommits_info_43_fpWen = RTL_PATH.io_diffCommits_info_43_fpWen; \
        force U_IF_NAME.io_diffCommits_info_43_vecWen = RTL_PATH.io_diffCommits_info_43_vecWen; \
        force U_IF_NAME.io_diffCommits_info_43_v0Wen = RTL_PATH.io_diffCommits_info_43_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_43_vlWen = RTL_PATH.io_diffCommits_info_43_vlWen; \
        force U_IF_NAME.io_diffCommits_info_44_ldest = RTL_PATH.io_diffCommits_info_44_ldest; \
        force U_IF_NAME.io_diffCommits_info_44_pdest = RTL_PATH.io_diffCommits_info_44_pdest; \
        force U_IF_NAME.io_diffCommits_info_44_rfWen = RTL_PATH.io_diffCommits_info_44_rfWen; \
        force U_IF_NAME.io_diffCommits_info_44_fpWen = RTL_PATH.io_diffCommits_info_44_fpWen; \
        force U_IF_NAME.io_diffCommits_info_44_vecWen = RTL_PATH.io_diffCommits_info_44_vecWen; \
        force U_IF_NAME.io_diffCommits_info_44_v0Wen = RTL_PATH.io_diffCommits_info_44_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_44_vlWen = RTL_PATH.io_diffCommits_info_44_vlWen; \
        force U_IF_NAME.io_diffCommits_info_45_ldest = RTL_PATH.io_diffCommits_info_45_ldest; \
        force U_IF_NAME.io_diffCommits_info_45_pdest = RTL_PATH.io_diffCommits_info_45_pdest; \
        force U_IF_NAME.io_diffCommits_info_45_rfWen = RTL_PATH.io_diffCommits_info_45_rfWen; \
        force U_IF_NAME.io_diffCommits_info_45_fpWen = RTL_PATH.io_diffCommits_info_45_fpWen; \
        force U_IF_NAME.io_diffCommits_info_45_vecWen = RTL_PATH.io_diffCommits_info_45_vecWen; \
        force U_IF_NAME.io_diffCommits_info_45_v0Wen = RTL_PATH.io_diffCommits_info_45_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_45_vlWen = RTL_PATH.io_diffCommits_info_45_vlWen; \
        force U_IF_NAME.io_diffCommits_info_46_ldest = RTL_PATH.io_diffCommits_info_46_ldest; \
        force U_IF_NAME.io_diffCommits_info_46_pdest = RTL_PATH.io_diffCommits_info_46_pdest; \
        force U_IF_NAME.io_diffCommits_info_46_rfWen = RTL_PATH.io_diffCommits_info_46_rfWen; \
        force U_IF_NAME.io_diffCommits_info_46_fpWen = RTL_PATH.io_diffCommits_info_46_fpWen; \
        force U_IF_NAME.io_diffCommits_info_46_vecWen = RTL_PATH.io_diffCommits_info_46_vecWen; \
        force U_IF_NAME.io_diffCommits_info_46_v0Wen = RTL_PATH.io_diffCommits_info_46_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_46_vlWen = RTL_PATH.io_diffCommits_info_46_vlWen; \
        force U_IF_NAME.io_diffCommits_info_47_ldest = RTL_PATH.io_diffCommits_info_47_ldest; \
        force U_IF_NAME.io_diffCommits_info_47_pdest = RTL_PATH.io_diffCommits_info_47_pdest; \
        force U_IF_NAME.io_diffCommits_info_47_rfWen = RTL_PATH.io_diffCommits_info_47_rfWen; \
        force U_IF_NAME.io_diffCommits_info_47_fpWen = RTL_PATH.io_diffCommits_info_47_fpWen; \
        force U_IF_NAME.io_diffCommits_info_47_vecWen = RTL_PATH.io_diffCommits_info_47_vecWen; \
        force U_IF_NAME.io_diffCommits_info_47_v0Wen = RTL_PATH.io_diffCommits_info_47_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_47_vlWen = RTL_PATH.io_diffCommits_info_47_vlWen; \
        force U_IF_NAME.io_diffCommits_info_48_ldest = RTL_PATH.io_diffCommits_info_48_ldest; \
        force U_IF_NAME.io_diffCommits_info_48_pdest = RTL_PATH.io_diffCommits_info_48_pdest; \
        force U_IF_NAME.io_diffCommits_info_48_rfWen = RTL_PATH.io_diffCommits_info_48_rfWen; \
        force U_IF_NAME.io_diffCommits_info_48_fpWen = RTL_PATH.io_diffCommits_info_48_fpWen; \
        force U_IF_NAME.io_diffCommits_info_48_vecWen = RTL_PATH.io_diffCommits_info_48_vecWen; \
        force U_IF_NAME.io_diffCommits_info_48_v0Wen = RTL_PATH.io_diffCommits_info_48_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_48_vlWen = RTL_PATH.io_diffCommits_info_48_vlWen; \
        force U_IF_NAME.io_diffCommits_info_49_ldest = RTL_PATH.io_diffCommits_info_49_ldest; \
        force U_IF_NAME.io_diffCommits_info_49_pdest = RTL_PATH.io_diffCommits_info_49_pdest; \
        force U_IF_NAME.io_diffCommits_info_49_rfWen = RTL_PATH.io_diffCommits_info_49_rfWen; \
        force U_IF_NAME.io_diffCommits_info_49_fpWen = RTL_PATH.io_diffCommits_info_49_fpWen; \
        force U_IF_NAME.io_diffCommits_info_49_vecWen = RTL_PATH.io_diffCommits_info_49_vecWen; \
        force U_IF_NAME.io_diffCommits_info_49_v0Wen = RTL_PATH.io_diffCommits_info_49_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_49_vlWen = RTL_PATH.io_diffCommits_info_49_vlWen; \
        force U_IF_NAME.io_diffCommits_info_50_ldest = RTL_PATH.io_diffCommits_info_50_ldest; \
        force U_IF_NAME.io_diffCommits_info_50_pdest = RTL_PATH.io_diffCommits_info_50_pdest; \
        force U_IF_NAME.io_diffCommits_info_50_rfWen = RTL_PATH.io_diffCommits_info_50_rfWen; \
        force U_IF_NAME.io_diffCommits_info_50_fpWen = RTL_PATH.io_diffCommits_info_50_fpWen; \
        force U_IF_NAME.io_diffCommits_info_50_vecWen = RTL_PATH.io_diffCommits_info_50_vecWen; \
        force U_IF_NAME.io_diffCommits_info_50_v0Wen = RTL_PATH.io_diffCommits_info_50_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_50_vlWen = RTL_PATH.io_diffCommits_info_50_vlWen; \
        force U_IF_NAME.io_diffCommits_info_51_ldest = RTL_PATH.io_diffCommits_info_51_ldest; \
        force U_IF_NAME.io_diffCommits_info_51_pdest = RTL_PATH.io_diffCommits_info_51_pdest; \
        force U_IF_NAME.io_diffCommits_info_51_rfWen = RTL_PATH.io_diffCommits_info_51_rfWen; \
        force U_IF_NAME.io_diffCommits_info_51_fpWen = RTL_PATH.io_diffCommits_info_51_fpWen; \
        force U_IF_NAME.io_diffCommits_info_51_vecWen = RTL_PATH.io_diffCommits_info_51_vecWen; \
        force U_IF_NAME.io_diffCommits_info_51_v0Wen = RTL_PATH.io_diffCommits_info_51_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_51_vlWen = RTL_PATH.io_diffCommits_info_51_vlWen; \
        force U_IF_NAME.io_diffCommits_info_52_ldest = RTL_PATH.io_diffCommits_info_52_ldest; \
        force U_IF_NAME.io_diffCommits_info_52_pdest = RTL_PATH.io_diffCommits_info_52_pdest; \
        force U_IF_NAME.io_diffCommits_info_52_rfWen = RTL_PATH.io_diffCommits_info_52_rfWen; \
        force U_IF_NAME.io_diffCommits_info_52_fpWen = RTL_PATH.io_diffCommits_info_52_fpWen; \
        force U_IF_NAME.io_diffCommits_info_52_vecWen = RTL_PATH.io_diffCommits_info_52_vecWen; \
        force U_IF_NAME.io_diffCommits_info_52_v0Wen = RTL_PATH.io_diffCommits_info_52_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_52_vlWen = RTL_PATH.io_diffCommits_info_52_vlWen; \
        force U_IF_NAME.io_diffCommits_info_53_ldest = RTL_PATH.io_diffCommits_info_53_ldest; \
        force U_IF_NAME.io_diffCommits_info_53_pdest = RTL_PATH.io_diffCommits_info_53_pdest; \
        force U_IF_NAME.io_diffCommits_info_53_rfWen = RTL_PATH.io_diffCommits_info_53_rfWen; \
        force U_IF_NAME.io_diffCommits_info_53_fpWen = RTL_PATH.io_diffCommits_info_53_fpWen; \
        force U_IF_NAME.io_diffCommits_info_53_vecWen = RTL_PATH.io_diffCommits_info_53_vecWen; \
        force U_IF_NAME.io_diffCommits_info_53_v0Wen = RTL_PATH.io_diffCommits_info_53_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_53_vlWen = RTL_PATH.io_diffCommits_info_53_vlWen; \
        force U_IF_NAME.io_diffCommits_info_54_ldest = RTL_PATH.io_diffCommits_info_54_ldest; \
        force U_IF_NAME.io_diffCommits_info_54_pdest = RTL_PATH.io_diffCommits_info_54_pdest; \
        force U_IF_NAME.io_diffCommits_info_54_rfWen = RTL_PATH.io_diffCommits_info_54_rfWen; \
        force U_IF_NAME.io_diffCommits_info_54_fpWen = RTL_PATH.io_diffCommits_info_54_fpWen; \
        force U_IF_NAME.io_diffCommits_info_54_vecWen = RTL_PATH.io_diffCommits_info_54_vecWen; \
        force U_IF_NAME.io_diffCommits_info_54_v0Wen = RTL_PATH.io_diffCommits_info_54_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_54_vlWen = RTL_PATH.io_diffCommits_info_54_vlWen; \
        force U_IF_NAME.io_diffCommits_info_55_ldest = RTL_PATH.io_diffCommits_info_55_ldest; \
        force U_IF_NAME.io_diffCommits_info_55_pdest = RTL_PATH.io_diffCommits_info_55_pdest; \
        force U_IF_NAME.io_diffCommits_info_55_rfWen = RTL_PATH.io_diffCommits_info_55_rfWen; \
        force U_IF_NAME.io_diffCommits_info_55_fpWen = RTL_PATH.io_diffCommits_info_55_fpWen; \
        force U_IF_NAME.io_diffCommits_info_55_vecWen = RTL_PATH.io_diffCommits_info_55_vecWen; \
        force U_IF_NAME.io_diffCommits_info_55_v0Wen = RTL_PATH.io_diffCommits_info_55_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_55_vlWen = RTL_PATH.io_diffCommits_info_55_vlWen; \
        force U_IF_NAME.io_diffCommits_info_56_ldest = RTL_PATH.io_diffCommits_info_56_ldest; \
        force U_IF_NAME.io_diffCommits_info_56_pdest = RTL_PATH.io_diffCommits_info_56_pdest; \
        force U_IF_NAME.io_diffCommits_info_56_rfWen = RTL_PATH.io_diffCommits_info_56_rfWen; \
        force U_IF_NAME.io_diffCommits_info_56_fpWen = RTL_PATH.io_diffCommits_info_56_fpWen; \
        force U_IF_NAME.io_diffCommits_info_56_vecWen = RTL_PATH.io_diffCommits_info_56_vecWen; \
        force U_IF_NAME.io_diffCommits_info_56_v0Wen = RTL_PATH.io_diffCommits_info_56_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_56_vlWen = RTL_PATH.io_diffCommits_info_56_vlWen; \
        force U_IF_NAME.io_diffCommits_info_57_ldest = RTL_PATH.io_diffCommits_info_57_ldest; \
        force U_IF_NAME.io_diffCommits_info_57_pdest = RTL_PATH.io_diffCommits_info_57_pdest; \
        force U_IF_NAME.io_diffCommits_info_57_rfWen = RTL_PATH.io_diffCommits_info_57_rfWen; \
        force U_IF_NAME.io_diffCommits_info_57_fpWen = RTL_PATH.io_diffCommits_info_57_fpWen; \
        force U_IF_NAME.io_diffCommits_info_57_vecWen = RTL_PATH.io_diffCommits_info_57_vecWen; \
        force U_IF_NAME.io_diffCommits_info_57_v0Wen = RTL_PATH.io_diffCommits_info_57_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_57_vlWen = RTL_PATH.io_diffCommits_info_57_vlWen; \
        force U_IF_NAME.io_diffCommits_info_58_ldest = RTL_PATH.io_diffCommits_info_58_ldest; \
        force U_IF_NAME.io_diffCommits_info_58_pdest = RTL_PATH.io_diffCommits_info_58_pdest; \
        force U_IF_NAME.io_diffCommits_info_58_rfWen = RTL_PATH.io_diffCommits_info_58_rfWen; \
        force U_IF_NAME.io_diffCommits_info_58_fpWen = RTL_PATH.io_diffCommits_info_58_fpWen; \
        force U_IF_NAME.io_diffCommits_info_58_vecWen = RTL_PATH.io_diffCommits_info_58_vecWen; \
        force U_IF_NAME.io_diffCommits_info_58_v0Wen = RTL_PATH.io_diffCommits_info_58_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_58_vlWen = RTL_PATH.io_diffCommits_info_58_vlWen; \
        force U_IF_NAME.io_diffCommits_info_59_ldest = RTL_PATH.io_diffCommits_info_59_ldest; \
        force U_IF_NAME.io_diffCommits_info_59_pdest = RTL_PATH.io_diffCommits_info_59_pdest; \
        force U_IF_NAME.io_diffCommits_info_59_rfWen = RTL_PATH.io_diffCommits_info_59_rfWen; \
        force U_IF_NAME.io_diffCommits_info_59_fpWen = RTL_PATH.io_diffCommits_info_59_fpWen; \
        force U_IF_NAME.io_diffCommits_info_59_vecWen = RTL_PATH.io_diffCommits_info_59_vecWen; \
        force U_IF_NAME.io_diffCommits_info_59_v0Wen = RTL_PATH.io_diffCommits_info_59_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_59_vlWen = RTL_PATH.io_diffCommits_info_59_vlWen; \
        force U_IF_NAME.io_diffCommits_info_60_ldest = RTL_PATH.io_diffCommits_info_60_ldest; \
        force U_IF_NAME.io_diffCommits_info_60_pdest = RTL_PATH.io_diffCommits_info_60_pdest; \
        force U_IF_NAME.io_diffCommits_info_60_rfWen = RTL_PATH.io_diffCommits_info_60_rfWen; \
        force U_IF_NAME.io_diffCommits_info_60_fpWen = RTL_PATH.io_diffCommits_info_60_fpWen; \
        force U_IF_NAME.io_diffCommits_info_60_vecWen = RTL_PATH.io_diffCommits_info_60_vecWen; \
        force U_IF_NAME.io_diffCommits_info_60_v0Wen = RTL_PATH.io_diffCommits_info_60_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_60_vlWen = RTL_PATH.io_diffCommits_info_60_vlWen; \
        force U_IF_NAME.io_diffCommits_info_61_ldest = RTL_PATH.io_diffCommits_info_61_ldest; \
        force U_IF_NAME.io_diffCommits_info_61_pdest = RTL_PATH.io_diffCommits_info_61_pdest; \
        force U_IF_NAME.io_diffCommits_info_61_rfWen = RTL_PATH.io_diffCommits_info_61_rfWen; \
        force U_IF_NAME.io_diffCommits_info_61_fpWen = RTL_PATH.io_diffCommits_info_61_fpWen; \
        force U_IF_NAME.io_diffCommits_info_61_vecWen = RTL_PATH.io_diffCommits_info_61_vecWen; \
        force U_IF_NAME.io_diffCommits_info_61_v0Wen = RTL_PATH.io_diffCommits_info_61_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_61_vlWen = RTL_PATH.io_diffCommits_info_61_vlWen; \
        force U_IF_NAME.io_diffCommits_info_62_ldest = RTL_PATH.io_diffCommits_info_62_ldest; \
        force U_IF_NAME.io_diffCommits_info_62_pdest = RTL_PATH.io_diffCommits_info_62_pdest; \
        force U_IF_NAME.io_diffCommits_info_62_rfWen = RTL_PATH.io_diffCommits_info_62_rfWen; \
        force U_IF_NAME.io_diffCommits_info_62_fpWen = RTL_PATH.io_diffCommits_info_62_fpWen; \
        force U_IF_NAME.io_diffCommits_info_62_vecWen = RTL_PATH.io_diffCommits_info_62_vecWen; \
        force U_IF_NAME.io_diffCommits_info_62_v0Wen = RTL_PATH.io_diffCommits_info_62_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_62_vlWen = RTL_PATH.io_diffCommits_info_62_vlWen; \
        force U_IF_NAME.io_diffCommits_info_63_ldest = RTL_PATH.io_diffCommits_info_63_ldest; \
        force U_IF_NAME.io_diffCommits_info_63_pdest = RTL_PATH.io_diffCommits_info_63_pdest; \
        force U_IF_NAME.io_diffCommits_info_63_rfWen = RTL_PATH.io_diffCommits_info_63_rfWen; \
        force U_IF_NAME.io_diffCommits_info_63_fpWen = RTL_PATH.io_diffCommits_info_63_fpWen; \
        force U_IF_NAME.io_diffCommits_info_63_vecWen = RTL_PATH.io_diffCommits_info_63_vecWen; \
        force U_IF_NAME.io_diffCommits_info_63_v0Wen = RTL_PATH.io_diffCommits_info_63_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_63_vlWen = RTL_PATH.io_diffCommits_info_63_vlWen; \
        force U_IF_NAME.io_diffCommits_info_64_ldest = RTL_PATH.io_diffCommits_info_64_ldest; \
        force U_IF_NAME.io_diffCommits_info_64_pdest = RTL_PATH.io_diffCommits_info_64_pdest; \
        force U_IF_NAME.io_diffCommits_info_64_rfWen = RTL_PATH.io_diffCommits_info_64_rfWen; \
        force U_IF_NAME.io_diffCommits_info_64_fpWen = RTL_PATH.io_diffCommits_info_64_fpWen; \
        force U_IF_NAME.io_diffCommits_info_64_vecWen = RTL_PATH.io_diffCommits_info_64_vecWen; \
        force U_IF_NAME.io_diffCommits_info_64_v0Wen = RTL_PATH.io_diffCommits_info_64_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_64_vlWen = RTL_PATH.io_diffCommits_info_64_vlWen; \
        force U_IF_NAME.io_diffCommits_info_65_ldest = RTL_PATH.io_diffCommits_info_65_ldest; \
        force U_IF_NAME.io_diffCommits_info_65_pdest = RTL_PATH.io_diffCommits_info_65_pdest; \
        force U_IF_NAME.io_diffCommits_info_65_rfWen = RTL_PATH.io_diffCommits_info_65_rfWen; \
        force U_IF_NAME.io_diffCommits_info_65_fpWen = RTL_PATH.io_diffCommits_info_65_fpWen; \
        force U_IF_NAME.io_diffCommits_info_65_vecWen = RTL_PATH.io_diffCommits_info_65_vecWen; \
        force U_IF_NAME.io_diffCommits_info_65_v0Wen = RTL_PATH.io_diffCommits_info_65_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_65_vlWen = RTL_PATH.io_diffCommits_info_65_vlWen; \
        force U_IF_NAME.io_diffCommits_info_66_ldest = RTL_PATH.io_diffCommits_info_66_ldest; \
        force U_IF_NAME.io_diffCommits_info_66_pdest = RTL_PATH.io_diffCommits_info_66_pdest; \
        force U_IF_NAME.io_diffCommits_info_66_rfWen = RTL_PATH.io_diffCommits_info_66_rfWen; \
        force U_IF_NAME.io_diffCommits_info_66_fpWen = RTL_PATH.io_diffCommits_info_66_fpWen; \
        force U_IF_NAME.io_diffCommits_info_66_vecWen = RTL_PATH.io_diffCommits_info_66_vecWen; \
        force U_IF_NAME.io_diffCommits_info_66_v0Wen = RTL_PATH.io_diffCommits_info_66_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_66_vlWen = RTL_PATH.io_diffCommits_info_66_vlWen; \
        force U_IF_NAME.io_diffCommits_info_67_ldest = RTL_PATH.io_diffCommits_info_67_ldest; \
        force U_IF_NAME.io_diffCommits_info_67_pdest = RTL_PATH.io_diffCommits_info_67_pdest; \
        force U_IF_NAME.io_diffCommits_info_67_rfWen = RTL_PATH.io_diffCommits_info_67_rfWen; \
        force U_IF_NAME.io_diffCommits_info_67_fpWen = RTL_PATH.io_diffCommits_info_67_fpWen; \
        force U_IF_NAME.io_diffCommits_info_67_vecWen = RTL_PATH.io_diffCommits_info_67_vecWen; \
        force U_IF_NAME.io_diffCommits_info_67_v0Wen = RTL_PATH.io_diffCommits_info_67_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_67_vlWen = RTL_PATH.io_diffCommits_info_67_vlWen; \
        force U_IF_NAME.io_diffCommits_info_68_ldest = RTL_PATH.io_diffCommits_info_68_ldest; \
        force U_IF_NAME.io_diffCommits_info_68_pdest = RTL_PATH.io_diffCommits_info_68_pdest; \
        force U_IF_NAME.io_diffCommits_info_68_rfWen = RTL_PATH.io_diffCommits_info_68_rfWen; \
        force U_IF_NAME.io_diffCommits_info_68_fpWen = RTL_PATH.io_diffCommits_info_68_fpWen; \
        force U_IF_NAME.io_diffCommits_info_68_vecWen = RTL_PATH.io_diffCommits_info_68_vecWen; \
        force U_IF_NAME.io_diffCommits_info_68_v0Wen = RTL_PATH.io_diffCommits_info_68_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_68_vlWen = RTL_PATH.io_diffCommits_info_68_vlWen; \
        force U_IF_NAME.io_diffCommits_info_69_ldest = RTL_PATH.io_diffCommits_info_69_ldest; \
        force U_IF_NAME.io_diffCommits_info_69_pdest = RTL_PATH.io_diffCommits_info_69_pdest; \
        force U_IF_NAME.io_diffCommits_info_69_rfWen = RTL_PATH.io_diffCommits_info_69_rfWen; \
        force U_IF_NAME.io_diffCommits_info_69_fpWen = RTL_PATH.io_diffCommits_info_69_fpWen; \
        force U_IF_NAME.io_diffCommits_info_69_vecWen = RTL_PATH.io_diffCommits_info_69_vecWen; \
        force U_IF_NAME.io_diffCommits_info_69_v0Wen = RTL_PATH.io_diffCommits_info_69_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_69_vlWen = RTL_PATH.io_diffCommits_info_69_vlWen; \
        force U_IF_NAME.io_diffCommits_info_70_ldest = RTL_PATH.io_diffCommits_info_70_ldest; \
        force U_IF_NAME.io_diffCommits_info_70_pdest = RTL_PATH.io_diffCommits_info_70_pdest; \
        force U_IF_NAME.io_diffCommits_info_70_rfWen = RTL_PATH.io_diffCommits_info_70_rfWen; \
        force U_IF_NAME.io_diffCommits_info_70_fpWen = RTL_PATH.io_diffCommits_info_70_fpWen; \
        force U_IF_NAME.io_diffCommits_info_70_vecWen = RTL_PATH.io_diffCommits_info_70_vecWen; \
        force U_IF_NAME.io_diffCommits_info_70_v0Wen = RTL_PATH.io_diffCommits_info_70_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_70_vlWen = RTL_PATH.io_diffCommits_info_70_vlWen; \
        force U_IF_NAME.io_diffCommits_info_71_ldest = RTL_PATH.io_diffCommits_info_71_ldest; \
        force U_IF_NAME.io_diffCommits_info_71_pdest = RTL_PATH.io_diffCommits_info_71_pdest; \
        force U_IF_NAME.io_diffCommits_info_71_rfWen = RTL_PATH.io_diffCommits_info_71_rfWen; \
        force U_IF_NAME.io_diffCommits_info_71_fpWen = RTL_PATH.io_diffCommits_info_71_fpWen; \
        force U_IF_NAME.io_diffCommits_info_71_vecWen = RTL_PATH.io_diffCommits_info_71_vecWen; \
        force U_IF_NAME.io_diffCommits_info_71_v0Wen = RTL_PATH.io_diffCommits_info_71_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_71_vlWen = RTL_PATH.io_diffCommits_info_71_vlWen; \
        force U_IF_NAME.io_diffCommits_info_72_ldest = RTL_PATH.io_diffCommits_info_72_ldest; \
        force U_IF_NAME.io_diffCommits_info_72_pdest = RTL_PATH.io_diffCommits_info_72_pdest; \
        force U_IF_NAME.io_diffCommits_info_72_rfWen = RTL_PATH.io_diffCommits_info_72_rfWen; \
        force U_IF_NAME.io_diffCommits_info_72_fpWen = RTL_PATH.io_diffCommits_info_72_fpWen; \
        force U_IF_NAME.io_diffCommits_info_72_vecWen = RTL_PATH.io_diffCommits_info_72_vecWen; \
        force U_IF_NAME.io_diffCommits_info_72_v0Wen = RTL_PATH.io_diffCommits_info_72_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_72_vlWen = RTL_PATH.io_diffCommits_info_72_vlWen; \
        force U_IF_NAME.io_diffCommits_info_73_ldest = RTL_PATH.io_diffCommits_info_73_ldest; \
        force U_IF_NAME.io_diffCommits_info_73_pdest = RTL_PATH.io_diffCommits_info_73_pdest; \
        force U_IF_NAME.io_diffCommits_info_73_rfWen = RTL_PATH.io_diffCommits_info_73_rfWen; \
        force U_IF_NAME.io_diffCommits_info_73_fpWen = RTL_PATH.io_diffCommits_info_73_fpWen; \
        force U_IF_NAME.io_diffCommits_info_73_vecWen = RTL_PATH.io_diffCommits_info_73_vecWen; \
        force U_IF_NAME.io_diffCommits_info_73_v0Wen = RTL_PATH.io_diffCommits_info_73_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_73_vlWen = RTL_PATH.io_diffCommits_info_73_vlWen; \
        force U_IF_NAME.io_diffCommits_info_74_ldest = RTL_PATH.io_diffCommits_info_74_ldest; \
        force U_IF_NAME.io_diffCommits_info_74_pdest = RTL_PATH.io_diffCommits_info_74_pdest; \
        force U_IF_NAME.io_diffCommits_info_74_rfWen = RTL_PATH.io_diffCommits_info_74_rfWen; \
        force U_IF_NAME.io_diffCommits_info_74_fpWen = RTL_PATH.io_diffCommits_info_74_fpWen; \
        force U_IF_NAME.io_diffCommits_info_74_vecWen = RTL_PATH.io_diffCommits_info_74_vecWen; \
        force U_IF_NAME.io_diffCommits_info_74_v0Wen = RTL_PATH.io_diffCommits_info_74_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_74_vlWen = RTL_PATH.io_diffCommits_info_74_vlWen; \
        force U_IF_NAME.io_diffCommits_info_75_ldest = RTL_PATH.io_diffCommits_info_75_ldest; \
        force U_IF_NAME.io_diffCommits_info_75_pdest = RTL_PATH.io_diffCommits_info_75_pdest; \
        force U_IF_NAME.io_diffCommits_info_75_rfWen = RTL_PATH.io_diffCommits_info_75_rfWen; \
        force U_IF_NAME.io_diffCommits_info_75_fpWen = RTL_PATH.io_diffCommits_info_75_fpWen; \
        force U_IF_NAME.io_diffCommits_info_75_vecWen = RTL_PATH.io_diffCommits_info_75_vecWen; \
        force U_IF_NAME.io_diffCommits_info_75_v0Wen = RTL_PATH.io_diffCommits_info_75_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_75_vlWen = RTL_PATH.io_diffCommits_info_75_vlWen; \
        force U_IF_NAME.io_diffCommits_info_76_ldest = RTL_PATH.io_diffCommits_info_76_ldest; \
        force U_IF_NAME.io_diffCommits_info_76_pdest = RTL_PATH.io_diffCommits_info_76_pdest; \
        force U_IF_NAME.io_diffCommits_info_76_rfWen = RTL_PATH.io_diffCommits_info_76_rfWen; \
        force U_IF_NAME.io_diffCommits_info_76_fpWen = RTL_PATH.io_diffCommits_info_76_fpWen; \
        force U_IF_NAME.io_diffCommits_info_76_vecWen = RTL_PATH.io_diffCommits_info_76_vecWen; \
        force U_IF_NAME.io_diffCommits_info_76_v0Wen = RTL_PATH.io_diffCommits_info_76_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_76_vlWen = RTL_PATH.io_diffCommits_info_76_vlWen; \
        force U_IF_NAME.io_diffCommits_info_77_ldest = RTL_PATH.io_diffCommits_info_77_ldest; \
        force U_IF_NAME.io_diffCommits_info_77_pdest = RTL_PATH.io_diffCommits_info_77_pdest; \
        force U_IF_NAME.io_diffCommits_info_77_rfWen = RTL_PATH.io_diffCommits_info_77_rfWen; \
        force U_IF_NAME.io_diffCommits_info_77_fpWen = RTL_PATH.io_diffCommits_info_77_fpWen; \
        force U_IF_NAME.io_diffCommits_info_77_vecWen = RTL_PATH.io_diffCommits_info_77_vecWen; \
        force U_IF_NAME.io_diffCommits_info_77_v0Wen = RTL_PATH.io_diffCommits_info_77_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_77_vlWen = RTL_PATH.io_diffCommits_info_77_vlWen; \
        force U_IF_NAME.io_diffCommits_info_78_ldest = RTL_PATH.io_diffCommits_info_78_ldest; \
        force U_IF_NAME.io_diffCommits_info_78_pdest = RTL_PATH.io_diffCommits_info_78_pdest; \
        force U_IF_NAME.io_diffCommits_info_78_rfWen = RTL_PATH.io_diffCommits_info_78_rfWen; \
        force U_IF_NAME.io_diffCommits_info_78_fpWen = RTL_PATH.io_diffCommits_info_78_fpWen; \
        force U_IF_NAME.io_diffCommits_info_78_vecWen = RTL_PATH.io_diffCommits_info_78_vecWen; \
        force U_IF_NAME.io_diffCommits_info_78_v0Wen = RTL_PATH.io_diffCommits_info_78_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_78_vlWen = RTL_PATH.io_diffCommits_info_78_vlWen; \
        force U_IF_NAME.io_diffCommits_info_79_ldest = RTL_PATH.io_diffCommits_info_79_ldest; \
        force U_IF_NAME.io_diffCommits_info_79_pdest = RTL_PATH.io_diffCommits_info_79_pdest; \
        force U_IF_NAME.io_diffCommits_info_79_rfWen = RTL_PATH.io_diffCommits_info_79_rfWen; \
        force U_IF_NAME.io_diffCommits_info_79_fpWen = RTL_PATH.io_diffCommits_info_79_fpWen; \
        force U_IF_NAME.io_diffCommits_info_79_vecWen = RTL_PATH.io_diffCommits_info_79_vecWen; \
        force U_IF_NAME.io_diffCommits_info_79_v0Wen = RTL_PATH.io_diffCommits_info_79_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_79_vlWen = RTL_PATH.io_diffCommits_info_79_vlWen; \
        force U_IF_NAME.io_diffCommits_info_80_ldest = RTL_PATH.io_diffCommits_info_80_ldest; \
        force U_IF_NAME.io_diffCommits_info_80_pdest = RTL_PATH.io_diffCommits_info_80_pdest; \
        force U_IF_NAME.io_diffCommits_info_80_rfWen = RTL_PATH.io_diffCommits_info_80_rfWen; \
        force U_IF_NAME.io_diffCommits_info_80_fpWen = RTL_PATH.io_diffCommits_info_80_fpWen; \
        force U_IF_NAME.io_diffCommits_info_80_vecWen = RTL_PATH.io_diffCommits_info_80_vecWen; \
        force U_IF_NAME.io_diffCommits_info_80_v0Wen = RTL_PATH.io_diffCommits_info_80_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_80_vlWen = RTL_PATH.io_diffCommits_info_80_vlWen; \
        force U_IF_NAME.io_diffCommits_info_81_ldest = RTL_PATH.io_diffCommits_info_81_ldest; \
        force U_IF_NAME.io_diffCommits_info_81_pdest = RTL_PATH.io_diffCommits_info_81_pdest; \
        force U_IF_NAME.io_diffCommits_info_81_rfWen = RTL_PATH.io_diffCommits_info_81_rfWen; \
        force U_IF_NAME.io_diffCommits_info_81_fpWen = RTL_PATH.io_diffCommits_info_81_fpWen; \
        force U_IF_NAME.io_diffCommits_info_81_vecWen = RTL_PATH.io_diffCommits_info_81_vecWen; \
        force U_IF_NAME.io_diffCommits_info_81_v0Wen = RTL_PATH.io_diffCommits_info_81_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_81_vlWen = RTL_PATH.io_diffCommits_info_81_vlWen; \
        force U_IF_NAME.io_diffCommits_info_82_ldest = RTL_PATH.io_diffCommits_info_82_ldest; \
        force U_IF_NAME.io_diffCommits_info_82_pdest = RTL_PATH.io_diffCommits_info_82_pdest; \
        force U_IF_NAME.io_diffCommits_info_82_rfWen = RTL_PATH.io_diffCommits_info_82_rfWen; \
        force U_IF_NAME.io_diffCommits_info_82_fpWen = RTL_PATH.io_diffCommits_info_82_fpWen; \
        force U_IF_NAME.io_diffCommits_info_82_vecWen = RTL_PATH.io_diffCommits_info_82_vecWen; \
        force U_IF_NAME.io_diffCommits_info_82_v0Wen = RTL_PATH.io_diffCommits_info_82_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_82_vlWen = RTL_PATH.io_diffCommits_info_82_vlWen; \
        force U_IF_NAME.io_diffCommits_info_83_ldest = RTL_PATH.io_diffCommits_info_83_ldest; \
        force U_IF_NAME.io_diffCommits_info_83_pdest = RTL_PATH.io_diffCommits_info_83_pdest; \
        force U_IF_NAME.io_diffCommits_info_83_rfWen = RTL_PATH.io_diffCommits_info_83_rfWen; \
        force U_IF_NAME.io_diffCommits_info_83_fpWen = RTL_PATH.io_diffCommits_info_83_fpWen; \
        force U_IF_NAME.io_diffCommits_info_83_vecWen = RTL_PATH.io_diffCommits_info_83_vecWen; \
        force U_IF_NAME.io_diffCommits_info_83_v0Wen = RTL_PATH.io_diffCommits_info_83_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_83_vlWen = RTL_PATH.io_diffCommits_info_83_vlWen; \
        force U_IF_NAME.io_diffCommits_info_84_ldest = RTL_PATH.io_diffCommits_info_84_ldest; \
        force U_IF_NAME.io_diffCommits_info_84_pdest = RTL_PATH.io_diffCommits_info_84_pdest; \
        force U_IF_NAME.io_diffCommits_info_84_rfWen = RTL_PATH.io_diffCommits_info_84_rfWen; \
        force U_IF_NAME.io_diffCommits_info_84_fpWen = RTL_PATH.io_diffCommits_info_84_fpWen; \
        force U_IF_NAME.io_diffCommits_info_84_vecWen = RTL_PATH.io_diffCommits_info_84_vecWen; \
        force U_IF_NAME.io_diffCommits_info_84_v0Wen = RTL_PATH.io_diffCommits_info_84_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_84_vlWen = RTL_PATH.io_diffCommits_info_84_vlWen; \
        force U_IF_NAME.io_diffCommits_info_85_ldest = RTL_PATH.io_diffCommits_info_85_ldest; \
        force U_IF_NAME.io_diffCommits_info_85_pdest = RTL_PATH.io_diffCommits_info_85_pdest; \
        force U_IF_NAME.io_diffCommits_info_85_rfWen = RTL_PATH.io_diffCommits_info_85_rfWen; \
        force U_IF_NAME.io_diffCommits_info_85_fpWen = RTL_PATH.io_diffCommits_info_85_fpWen; \
        force U_IF_NAME.io_diffCommits_info_85_vecWen = RTL_PATH.io_diffCommits_info_85_vecWen; \
        force U_IF_NAME.io_diffCommits_info_85_v0Wen = RTL_PATH.io_diffCommits_info_85_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_85_vlWen = RTL_PATH.io_diffCommits_info_85_vlWen; \
        force U_IF_NAME.io_diffCommits_info_86_ldest = RTL_PATH.io_diffCommits_info_86_ldest; \
        force U_IF_NAME.io_diffCommits_info_86_pdest = RTL_PATH.io_diffCommits_info_86_pdest; \
        force U_IF_NAME.io_diffCommits_info_86_rfWen = RTL_PATH.io_diffCommits_info_86_rfWen; \
        force U_IF_NAME.io_diffCommits_info_86_fpWen = RTL_PATH.io_diffCommits_info_86_fpWen; \
        force U_IF_NAME.io_diffCommits_info_86_vecWen = RTL_PATH.io_diffCommits_info_86_vecWen; \
        force U_IF_NAME.io_diffCommits_info_86_v0Wen = RTL_PATH.io_diffCommits_info_86_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_86_vlWen = RTL_PATH.io_diffCommits_info_86_vlWen; \
        force U_IF_NAME.io_diffCommits_info_87_ldest = RTL_PATH.io_diffCommits_info_87_ldest; \
        force U_IF_NAME.io_diffCommits_info_87_pdest = RTL_PATH.io_diffCommits_info_87_pdest; \
        force U_IF_NAME.io_diffCommits_info_87_rfWen = RTL_PATH.io_diffCommits_info_87_rfWen; \
        force U_IF_NAME.io_diffCommits_info_87_fpWen = RTL_PATH.io_diffCommits_info_87_fpWen; \
        force U_IF_NAME.io_diffCommits_info_87_vecWen = RTL_PATH.io_diffCommits_info_87_vecWen; \
        force U_IF_NAME.io_diffCommits_info_87_v0Wen = RTL_PATH.io_diffCommits_info_87_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_87_vlWen = RTL_PATH.io_diffCommits_info_87_vlWen; \
        force U_IF_NAME.io_diffCommits_info_88_ldest = RTL_PATH.io_diffCommits_info_88_ldest; \
        force U_IF_NAME.io_diffCommits_info_88_pdest = RTL_PATH.io_diffCommits_info_88_pdest; \
        force U_IF_NAME.io_diffCommits_info_88_rfWen = RTL_PATH.io_diffCommits_info_88_rfWen; \
        force U_IF_NAME.io_diffCommits_info_88_fpWen = RTL_PATH.io_diffCommits_info_88_fpWen; \
        force U_IF_NAME.io_diffCommits_info_88_vecWen = RTL_PATH.io_diffCommits_info_88_vecWen; \
        force U_IF_NAME.io_diffCommits_info_88_v0Wen = RTL_PATH.io_diffCommits_info_88_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_88_vlWen = RTL_PATH.io_diffCommits_info_88_vlWen; \
        force U_IF_NAME.io_diffCommits_info_89_ldest = RTL_PATH.io_diffCommits_info_89_ldest; \
        force U_IF_NAME.io_diffCommits_info_89_pdest = RTL_PATH.io_diffCommits_info_89_pdest; \
        force U_IF_NAME.io_diffCommits_info_89_rfWen = RTL_PATH.io_diffCommits_info_89_rfWen; \
        force U_IF_NAME.io_diffCommits_info_89_fpWen = RTL_PATH.io_diffCommits_info_89_fpWen; \
        force U_IF_NAME.io_diffCommits_info_89_vecWen = RTL_PATH.io_diffCommits_info_89_vecWen; \
        force U_IF_NAME.io_diffCommits_info_89_v0Wen = RTL_PATH.io_diffCommits_info_89_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_89_vlWen = RTL_PATH.io_diffCommits_info_89_vlWen; \
        force U_IF_NAME.io_diffCommits_info_90_ldest = RTL_PATH.io_diffCommits_info_90_ldest; \
        force U_IF_NAME.io_diffCommits_info_90_pdest = RTL_PATH.io_diffCommits_info_90_pdest; \
        force U_IF_NAME.io_diffCommits_info_90_rfWen = RTL_PATH.io_diffCommits_info_90_rfWen; \
        force U_IF_NAME.io_diffCommits_info_90_fpWen = RTL_PATH.io_diffCommits_info_90_fpWen; \
        force U_IF_NAME.io_diffCommits_info_90_vecWen = RTL_PATH.io_diffCommits_info_90_vecWen; \
        force U_IF_NAME.io_diffCommits_info_90_v0Wen = RTL_PATH.io_diffCommits_info_90_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_90_vlWen = RTL_PATH.io_diffCommits_info_90_vlWen; \
        force U_IF_NAME.io_diffCommits_info_91_ldest = RTL_PATH.io_diffCommits_info_91_ldest; \
        force U_IF_NAME.io_diffCommits_info_91_pdest = RTL_PATH.io_diffCommits_info_91_pdest; \
        force U_IF_NAME.io_diffCommits_info_91_rfWen = RTL_PATH.io_diffCommits_info_91_rfWen; \
        force U_IF_NAME.io_diffCommits_info_91_fpWen = RTL_PATH.io_diffCommits_info_91_fpWen; \
        force U_IF_NAME.io_diffCommits_info_91_vecWen = RTL_PATH.io_diffCommits_info_91_vecWen; \
        force U_IF_NAME.io_diffCommits_info_91_v0Wen = RTL_PATH.io_diffCommits_info_91_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_91_vlWen = RTL_PATH.io_diffCommits_info_91_vlWen; \
        force U_IF_NAME.io_diffCommits_info_92_ldest = RTL_PATH.io_diffCommits_info_92_ldest; \
        force U_IF_NAME.io_diffCommits_info_92_pdest = RTL_PATH.io_diffCommits_info_92_pdest; \
        force U_IF_NAME.io_diffCommits_info_92_rfWen = RTL_PATH.io_diffCommits_info_92_rfWen; \
        force U_IF_NAME.io_diffCommits_info_92_fpWen = RTL_PATH.io_diffCommits_info_92_fpWen; \
        force U_IF_NAME.io_diffCommits_info_92_vecWen = RTL_PATH.io_diffCommits_info_92_vecWen; \
        force U_IF_NAME.io_diffCommits_info_92_v0Wen = RTL_PATH.io_diffCommits_info_92_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_92_vlWen = RTL_PATH.io_diffCommits_info_92_vlWen; \
        force U_IF_NAME.io_diffCommits_info_93_ldest = RTL_PATH.io_diffCommits_info_93_ldest; \
        force U_IF_NAME.io_diffCommits_info_93_pdest = RTL_PATH.io_diffCommits_info_93_pdest; \
        force U_IF_NAME.io_diffCommits_info_93_rfWen = RTL_PATH.io_diffCommits_info_93_rfWen; \
        force U_IF_NAME.io_diffCommits_info_93_fpWen = RTL_PATH.io_diffCommits_info_93_fpWen; \
        force U_IF_NAME.io_diffCommits_info_93_vecWen = RTL_PATH.io_diffCommits_info_93_vecWen; \
        force U_IF_NAME.io_diffCommits_info_93_v0Wen = RTL_PATH.io_diffCommits_info_93_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_93_vlWen = RTL_PATH.io_diffCommits_info_93_vlWen; \
        force U_IF_NAME.io_diffCommits_info_94_ldest = RTL_PATH.io_diffCommits_info_94_ldest; \
        force U_IF_NAME.io_diffCommits_info_94_pdest = RTL_PATH.io_diffCommits_info_94_pdest; \
        force U_IF_NAME.io_diffCommits_info_94_rfWen = RTL_PATH.io_diffCommits_info_94_rfWen; \
        force U_IF_NAME.io_diffCommits_info_94_fpWen = RTL_PATH.io_diffCommits_info_94_fpWen; \
        force U_IF_NAME.io_diffCommits_info_94_vecWen = RTL_PATH.io_diffCommits_info_94_vecWen; \
        force U_IF_NAME.io_diffCommits_info_94_v0Wen = RTL_PATH.io_diffCommits_info_94_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_94_vlWen = RTL_PATH.io_diffCommits_info_94_vlWen; \
        force U_IF_NAME.io_diffCommits_info_95_ldest = RTL_PATH.io_diffCommits_info_95_ldest; \
        force U_IF_NAME.io_diffCommits_info_95_pdest = RTL_PATH.io_diffCommits_info_95_pdest; \
        force U_IF_NAME.io_diffCommits_info_95_rfWen = RTL_PATH.io_diffCommits_info_95_rfWen; \
        force U_IF_NAME.io_diffCommits_info_95_fpWen = RTL_PATH.io_diffCommits_info_95_fpWen; \
        force U_IF_NAME.io_diffCommits_info_95_vecWen = RTL_PATH.io_diffCommits_info_95_vecWen; \
        force U_IF_NAME.io_diffCommits_info_95_v0Wen = RTL_PATH.io_diffCommits_info_95_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_95_vlWen = RTL_PATH.io_diffCommits_info_95_vlWen; \
        force U_IF_NAME.io_diffCommits_info_96_ldest = RTL_PATH.io_diffCommits_info_96_ldest; \
        force U_IF_NAME.io_diffCommits_info_96_pdest = RTL_PATH.io_diffCommits_info_96_pdest; \
        force U_IF_NAME.io_diffCommits_info_96_rfWen = RTL_PATH.io_diffCommits_info_96_rfWen; \
        force U_IF_NAME.io_diffCommits_info_96_fpWen = RTL_PATH.io_diffCommits_info_96_fpWen; \
        force U_IF_NAME.io_diffCommits_info_96_vecWen = RTL_PATH.io_diffCommits_info_96_vecWen; \
        force U_IF_NAME.io_diffCommits_info_96_v0Wen = RTL_PATH.io_diffCommits_info_96_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_96_vlWen = RTL_PATH.io_diffCommits_info_96_vlWen; \
        force U_IF_NAME.io_diffCommits_info_97_ldest = RTL_PATH.io_diffCommits_info_97_ldest; \
        force U_IF_NAME.io_diffCommits_info_97_pdest = RTL_PATH.io_diffCommits_info_97_pdest; \
        force U_IF_NAME.io_diffCommits_info_97_rfWen = RTL_PATH.io_diffCommits_info_97_rfWen; \
        force U_IF_NAME.io_diffCommits_info_97_fpWen = RTL_PATH.io_diffCommits_info_97_fpWen; \
        force U_IF_NAME.io_diffCommits_info_97_vecWen = RTL_PATH.io_diffCommits_info_97_vecWen; \
        force U_IF_NAME.io_diffCommits_info_97_v0Wen = RTL_PATH.io_diffCommits_info_97_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_97_vlWen = RTL_PATH.io_diffCommits_info_97_vlWen; \
        force U_IF_NAME.io_diffCommits_info_98_ldest = RTL_PATH.io_diffCommits_info_98_ldest; \
        force U_IF_NAME.io_diffCommits_info_98_pdest = RTL_PATH.io_diffCommits_info_98_pdest; \
        force U_IF_NAME.io_diffCommits_info_98_rfWen = RTL_PATH.io_diffCommits_info_98_rfWen; \
        force U_IF_NAME.io_diffCommits_info_98_fpWen = RTL_PATH.io_diffCommits_info_98_fpWen; \
        force U_IF_NAME.io_diffCommits_info_98_vecWen = RTL_PATH.io_diffCommits_info_98_vecWen; \
        force U_IF_NAME.io_diffCommits_info_98_v0Wen = RTL_PATH.io_diffCommits_info_98_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_98_vlWen = RTL_PATH.io_diffCommits_info_98_vlWen; \
        force U_IF_NAME.io_diffCommits_info_99_ldest = RTL_PATH.io_diffCommits_info_99_ldest; \
        force U_IF_NAME.io_diffCommits_info_99_pdest = RTL_PATH.io_diffCommits_info_99_pdest; \
        force U_IF_NAME.io_diffCommits_info_99_rfWen = RTL_PATH.io_diffCommits_info_99_rfWen; \
        force U_IF_NAME.io_diffCommits_info_99_fpWen = RTL_PATH.io_diffCommits_info_99_fpWen; \
        force U_IF_NAME.io_diffCommits_info_99_vecWen = RTL_PATH.io_diffCommits_info_99_vecWen; \
        force U_IF_NAME.io_diffCommits_info_99_v0Wen = RTL_PATH.io_diffCommits_info_99_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_99_vlWen = RTL_PATH.io_diffCommits_info_99_vlWen; \
        force U_IF_NAME.io_diffCommits_info_100_ldest = RTL_PATH.io_diffCommits_info_100_ldest; \
        force U_IF_NAME.io_diffCommits_info_100_pdest = RTL_PATH.io_diffCommits_info_100_pdest; \
        force U_IF_NAME.io_diffCommits_info_100_rfWen = RTL_PATH.io_diffCommits_info_100_rfWen; \
        force U_IF_NAME.io_diffCommits_info_100_fpWen = RTL_PATH.io_diffCommits_info_100_fpWen; \
        force U_IF_NAME.io_diffCommits_info_100_vecWen = RTL_PATH.io_diffCommits_info_100_vecWen; \
        force U_IF_NAME.io_diffCommits_info_100_v0Wen = RTL_PATH.io_diffCommits_info_100_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_100_vlWen = RTL_PATH.io_diffCommits_info_100_vlWen; \
        force U_IF_NAME.io_diffCommits_info_101_ldest = RTL_PATH.io_diffCommits_info_101_ldest; \
        force U_IF_NAME.io_diffCommits_info_101_pdest = RTL_PATH.io_diffCommits_info_101_pdest; \
        force U_IF_NAME.io_diffCommits_info_101_rfWen = RTL_PATH.io_diffCommits_info_101_rfWen; \
        force U_IF_NAME.io_diffCommits_info_101_fpWen = RTL_PATH.io_diffCommits_info_101_fpWen; \
        force U_IF_NAME.io_diffCommits_info_101_vecWen = RTL_PATH.io_diffCommits_info_101_vecWen; \
        force U_IF_NAME.io_diffCommits_info_101_v0Wen = RTL_PATH.io_diffCommits_info_101_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_101_vlWen = RTL_PATH.io_diffCommits_info_101_vlWen; \
        force U_IF_NAME.io_diffCommits_info_102_ldest = RTL_PATH.io_diffCommits_info_102_ldest; \
        force U_IF_NAME.io_diffCommits_info_102_pdest = RTL_PATH.io_diffCommits_info_102_pdest; \
        force U_IF_NAME.io_diffCommits_info_102_rfWen = RTL_PATH.io_diffCommits_info_102_rfWen; \
        force U_IF_NAME.io_diffCommits_info_102_fpWen = RTL_PATH.io_diffCommits_info_102_fpWen; \
        force U_IF_NAME.io_diffCommits_info_102_vecWen = RTL_PATH.io_diffCommits_info_102_vecWen; \
        force U_IF_NAME.io_diffCommits_info_102_v0Wen = RTL_PATH.io_diffCommits_info_102_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_102_vlWen = RTL_PATH.io_diffCommits_info_102_vlWen; \
        force U_IF_NAME.io_diffCommits_info_103_ldest = RTL_PATH.io_diffCommits_info_103_ldest; \
        force U_IF_NAME.io_diffCommits_info_103_pdest = RTL_PATH.io_diffCommits_info_103_pdest; \
        force U_IF_NAME.io_diffCommits_info_103_rfWen = RTL_PATH.io_diffCommits_info_103_rfWen; \
        force U_IF_NAME.io_diffCommits_info_103_fpWen = RTL_PATH.io_diffCommits_info_103_fpWen; \
        force U_IF_NAME.io_diffCommits_info_103_vecWen = RTL_PATH.io_diffCommits_info_103_vecWen; \
        force U_IF_NAME.io_diffCommits_info_103_v0Wen = RTL_PATH.io_diffCommits_info_103_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_103_vlWen = RTL_PATH.io_diffCommits_info_103_vlWen; \
        force U_IF_NAME.io_diffCommits_info_104_ldest = RTL_PATH.io_diffCommits_info_104_ldest; \
        force U_IF_NAME.io_diffCommits_info_104_pdest = RTL_PATH.io_diffCommits_info_104_pdest; \
        force U_IF_NAME.io_diffCommits_info_104_rfWen = RTL_PATH.io_diffCommits_info_104_rfWen; \
        force U_IF_NAME.io_diffCommits_info_104_fpWen = RTL_PATH.io_diffCommits_info_104_fpWen; \
        force U_IF_NAME.io_diffCommits_info_104_vecWen = RTL_PATH.io_diffCommits_info_104_vecWen; \
        force U_IF_NAME.io_diffCommits_info_104_v0Wen = RTL_PATH.io_diffCommits_info_104_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_104_vlWen = RTL_PATH.io_diffCommits_info_104_vlWen; \
        force U_IF_NAME.io_diffCommits_info_105_ldest = RTL_PATH.io_diffCommits_info_105_ldest; \
        force U_IF_NAME.io_diffCommits_info_105_pdest = RTL_PATH.io_diffCommits_info_105_pdest; \
        force U_IF_NAME.io_diffCommits_info_105_rfWen = RTL_PATH.io_diffCommits_info_105_rfWen; \
        force U_IF_NAME.io_diffCommits_info_105_fpWen = RTL_PATH.io_diffCommits_info_105_fpWen; \
        force U_IF_NAME.io_diffCommits_info_105_vecWen = RTL_PATH.io_diffCommits_info_105_vecWen; \
        force U_IF_NAME.io_diffCommits_info_105_v0Wen = RTL_PATH.io_diffCommits_info_105_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_105_vlWen = RTL_PATH.io_diffCommits_info_105_vlWen; \
        force U_IF_NAME.io_diffCommits_info_106_ldest = RTL_PATH.io_diffCommits_info_106_ldest; \
        force U_IF_NAME.io_diffCommits_info_106_pdest = RTL_PATH.io_diffCommits_info_106_pdest; \
        force U_IF_NAME.io_diffCommits_info_106_rfWen = RTL_PATH.io_diffCommits_info_106_rfWen; \
        force U_IF_NAME.io_diffCommits_info_106_fpWen = RTL_PATH.io_diffCommits_info_106_fpWen; \
        force U_IF_NAME.io_diffCommits_info_106_vecWen = RTL_PATH.io_diffCommits_info_106_vecWen; \
        force U_IF_NAME.io_diffCommits_info_106_v0Wen = RTL_PATH.io_diffCommits_info_106_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_106_vlWen = RTL_PATH.io_diffCommits_info_106_vlWen; \
        force U_IF_NAME.io_diffCommits_info_107_ldest = RTL_PATH.io_diffCommits_info_107_ldest; \
        force U_IF_NAME.io_diffCommits_info_107_pdest = RTL_PATH.io_diffCommits_info_107_pdest; \
        force U_IF_NAME.io_diffCommits_info_107_rfWen = RTL_PATH.io_diffCommits_info_107_rfWen; \
        force U_IF_NAME.io_diffCommits_info_107_fpWen = RTL_PATH.io_diffCommits_info_107_fpWen; \
        force U_IF_NAME.io_diffCommits_info_107_vecWen = RTL_PATH.io_diffCommits_info_107_vecWen; \
        force U_IF_NAME.io_diffCommits_info_107_v0Wen = RTL_PATH.io_diffCommits_info_107_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_107_vlWen = RTL_PATH.io_diffCommits_info_107_vlWen; \
        force U_IF_NAME.io_diffCommits_info_108_ldest = RTL_PATH.io_diffCommits_info_108_ldest; \
        force U_IF_NAME.io_diffCommits_info_108_pdest = RTL_PATH.io_diffCommits_info_108_pdest; \
        force U_IF_NAME.io_diffCommits_info_108_rfWen = RTL_PATH.io_diffCommits_info_108_rfWen; \
        force U_IF_NAME.io_diffCommits_info_108_fpWen = RTL_PATH.io_diffCommits_info_108_fpWen; \
        force U_IF_NAME.io_diffCommits_info_108_vecWen = RTL_PATH.io_diffCommits_info_108_vecWen; \
        force U_IF_NAME.io_diffCommits_info_108_v0Wen = RTL_PATH.io_diffCommits_info_108_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_108_vlWen = RTL_PATH.io_diffCommits_info_108_vlWen; \
        force U_IF_NAME.io_diffCommits_info_109_ldest = RTL_PATH.io_diffCommits_info_109_ldest; \
        force U_IF_NAME.io_diffCommits_info_109_pdest = RTL_PATH.io_diffCommits_info_109_pdest; \
        force U_IF_NAME.io_diffCommits_info_109_rfWen = RTL_PATH.io_diffCommits_info_109_rfWen; \
        force U_IF_NAME.io_diffCommits_info_109_fpWen = RTL_PATH.io_diffCommits_info_109_fpWen; \
        force U_IF_NAME.io_diffCommits_info_109_vecWen = RTL_PATH.io_diffCommits_info_109_vecWen; \
        force U_IF_NAME.io_diffCommits_info_109_v0Wen = RTL_PATH.io_diffCommits_info_109_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_109_vlWen = RTL_PATH.io_diffCommits_info_109_vlWen; \
        force U_IF_NAME.io_diffCommits_info_110_ldest = RTL_PATH.io_diffCommits_info_110_ldest; \
        force U_IF_NAME.io_diffCommits_info_110_pdest = RTL_PATH.io_diffCommits_info_110_pdest; \
        force U_IF_NAME.io_diffCommits_info_110_rfWen = RTL_PATH.io_diffCommits_info_110_rfWen; \
        force U_IF_NAME.io_diffCommits_info_110_fpWen = RTL_PATH.io_diffCommits_info_110_fpWen; \
        force U_IF_NAME.io_diffCommits_info_110_vecWen = RTL_PATH.io_diffCommits_info_110_vecWen; \
        force U_IF_NAME.io_diffCommits_info_110_v0Wen = RTL_PATH.io_diffCommits_info_110_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_110_vlWen = RTL_PATH.io_diffCommits_info_110_vlWen; \
        force U_IF_NAME.io_diffCommits_info_111_ldest = RTL_PATH.io_diffCommits_info_111_ldest; \
        force U_IF_NAME.io_diffCommits_info_111_pdest = RTL_PATH.io_diffCommits_info_111_pdest; \
        force U_IF_NAME.io_diffCommits_info_111_rfWen = RTL_PATH.io_diffCommits_info_111_rfWen; \
        force U_IF_NAME.io_diffCommits_info_111_fpWen = RTL_PATH.io_diffCommits_info_111_fpWen; \
        force U_IF_NAME.io_diffCommits_info_111_vecWen = RTL_PATH.io_diffCommits_info_111_vecWen; \
        force U_IF_NAME.io_diffCommits_info_111_v0Wen = RTL_PATH.io_diffCommits_info_111_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_111_vlWen = RTL_PATH.io_diffCommits_info_111_vlWen; \
        force U_IF_NAME.io_diffCommits_info_112_ldest = RTL_PATH.io_diffCommits_info_112_ldest; \
        force U_IF_NAME.io_diffCommits_info_112_pdest = RTL_PATH.io_diffCommits_info_112_pdest; \
        force U_IF_NAME.io_diffCommits_info_112_rfWen = RTL_PATH.io_diffCommits_info_112_rfWen; \
        force U_IF_NAME.io_diffCommits_info_112_fpWen = RTL_PATH.io_diffCommits_info_112_fpWen; \
        force U_IF_NAME.io_diffCommits_info_112_vecWen = RTL_PATH.io_diffCommits_info_112_vecWen; \
        force U_IF_NAME.io_diffCommits_info_112_v0Wen = RTL_PATH.io_diffCommits_info_112_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_112_vlWen = RTL_PATH.io_diffCommits_info_112_vlWen; \
        force U_IF_NAME.io_diffCommits_info_113_ldest = RTL_PATH.io_diffCommits_info_113_ldest; \
        force U_IF_NAME.io_diffCommits_info_113_pdest = RTL_PATH.io_diffCommits_info_113_pdest; \
        force U_IF_NAME.io_diffCommits_info_113_rfWen = RTL_PATH.io_diffCommits_info_113_rfWen; \
        force U_IF_NAME.io_diffCommits_info_113_fpWen = RTL_PATH.io_diffCommits_info_113_fpWen; \
        force U_IF_NAME.io_diffCommits_info_113_vecWen = RTL_PATH.io_diffCommits_info_113_vecWen; \
        force U_IF_NAME.io_diffCommits_info_113_v0Wen = RTL_PATH.io_diffCommits_info_113_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_113_vlWen = RTL_PATH.io_diffCommits_info_113_vlWen; \
        force U_IF_NAME.io_diffCommits_info_114_ldest = RTL_PATH.io_diffCommits_info_114_ldest; \
        force U_IF_NAME.io_diffCommits_info_114_pdest = RTL_PATH.io_diffCommits_info_114_pdest; \
        force U_IF_NAME.io_diffCommits_info_114_rfWen = RTL_PATH.io_diffCommits_info_114_rfWen; \
        force U_IF_NAME.io_diffCommits_info_114_fpWen = RTL_PATH.io_diffCommits_info_114_fpWen; \
        force U_IF_NAME.io_diffCommits_info_114_vecWen = RTL_PATH.io_diffCommits_info_114_vecWen; \
        force U_IF_NAME.io_diffCommits_info_114_v0Wen = RTL_PATH.io_diffCommits_info_114_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_114_vlWen = RTL_PATH.io_diffCommits_info_114_vlWen; \
        force U_IF_NAME.io_diffCommits_info_115_ldest = RTL_PATH.io_diffCommits_info_115_ldest; \
        force U_IF_NAME.io_diffCommits_info_115_pdest = RTL_PATH.io_diffCommits_info_115_pdest; \
        force U_IF_NAME.io_diffCommits_info_115_rfWen = RTL_PATH.io_diffCommits_info_115_rfWen; \
        force U_IF_NAME.io_diffCommits_info_115_fpWen = RTL_PATH.io_diffCommits_info_115_fpWen; \
        force U_IF_NAME.io_diffCommits_info_115_vecWen = RTL_PATH.io_diffCommits_info_115_vecWen; \
        force U_IF_NAME.io_diffCommits_info_115_v0Wen = RTL_PATH.io_diffCommits_info_115_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_115_vlWen = RTL_PATH.io_diffCommits_info_115_vlWen; \
        force U_IF_NAME.io_diffCommits_info_116_ldest = RTL_PATH.io_diffCommits_info_116_ldest; \
        force U_IF_NAME.io_diffCommits_info_116_pdest = RTL_PATH.io_diffCommits_info_116_pdest; \
        force U_IF_NAME.io_diffCommits_info_116_rfWen = RTL_PATH.io_diffCommits_info_116_rfWen; \
        force U_IF_NAME.io_diffCommits_info_116_fpWen = RTL_PATH.io_diffCommits_info_116_fpWen; \
        force U_IF_NAME.io_diffCommits_info_116_vecWen = RTL_PATH.io_diffCommits_info_116_vecWen; \
        force U_IF_NAME.io_diffCommits_info_116_v0Wen = RTL_PATH.io_diffCommits_info_116_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_116_vlWen = RTL_PATH.io_diffCommits_info_116_vlWen; \
        force U_IF_NAME.io_diffCommits_info_117_ldest = RTL_PATH.io_diffCommits_info_117_ldest; \
        force U_IF_NAME.io_diffCommits_info_117_pdest = RTL_PATH.io_diffCommits_info_117_pdest; \
        force U_IF_NAME.io_diffCommits_info_117_rfWen = RTL_PATH.io_diffCommits_info_117_rfWen; \
        force U_IF_NAME.io_diffCommits_info_117_fpWen = RTL_PATH.io_diffCommits_info_117_fpWen; \
        force U_IF_NAME.io_diffCommits_info_117_vecWen = RTL_PATH.io_diffCommits_info_117_vecWen; \
        force U_IF_NAME.io_diffCommits_info_117_v0Wen = RTL_PATH.io_diffCommits_info_117_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_117_vlWen = RTL_PATH.io_diffCommits_info_117_vlWen; \
        force U_IF_NAME.io_diffCommits_info_118_ldest = RTL_PATH.io_diffCommits_info_118_ldest; \
        force U_IF_NAME.io_diffCommits_info_118_pdest = RTL_PATH.io_diffCommits_info_118_pdest; \
        force U_IF_NAME.io_diffCommits_info_118_rfWen = RTL_PATH.io_diffCommits_info_118_rfWen; \
        force U_IF_NAME.io_diffCommits_info_118_fpWen = RTL_PATH.io_diffCommits_info_118_fpWen; \
        force U_IF_NAME.io_diffCommits_info_118_vecWen = RTL_PATH.io_diffCommits_info_118_vecWen; \
        force U_IF_NAME.io_diffCommits_info_118_v0Wen = RTL_PATH.io_diffCommits_info_118_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_118_vlWen = RTL_PATH.io_diffCommits_info_118_vlWen; \
        force U_IF_NAME.io_diffCommits_info_119_ldest = RTL_PATH.io_diffCommits_info_119_ldest; \
        force U_IF_NAME.io_diffCommits_info_119_pdest = RTL_PATH.io_diffCommits_info_119_pdest; \
        force U_IF_NAME.io_diffCommits_info_119_rfWen = RTL_PATH.io_diffCommits_info_119_rfWen; \
        force U_IF_NAME.io_diffCommits_info_119_fpWen = RTL_PATH.io_diffCommits_info_119_fpWen; \
        force U_IF_NAME.io_diffCommits_info_119_vecWen = RTL_PATH.io_diffCommits_info_119_vecWen; \
        force U_IF_NAME.io_diffCommits_info_119_v0Wen = RTL_PATH.io_diffCommits_info_119_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_119_vlWen = RTL_PATH.io_diffCommits_info_119_vlWen; \
        force U_IF_NAME.io_diffCommits_info_120_ldest = RTL_PATH.io_diffCommits_info_120_ldest; \
        force U_IF_NAME.io_diffCommits_info_120_pdest = RTL_PATH.io_diffCommits_info_120_pdest; \
        force U_IF_NAME.io_diffCommits_info_120_rfWen = RTL_PATH.io_diffCommits_info_120_rfWen; \
        force U_IF_NAME.io_diffCommits_info_120_fpWen = RTL_PATH.io_diffCommits_info_120_fpWen; \
        force U_IF_NAME.io_diffCommits_info_120_vecWen = RTL_PATH.io_diffCommits_info_120_vecWen; \
        force U_IF_NAME.io_diffCommits_info_120_v0Wen = RTL_PATH.io_diffCommits_info_120_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_120_vlWen = RTL_PATH.io_diffCommits_info_120_vlWen; \
        force U_IF_NAME.io_diffCommits_info_121_ldest = RTL_PATH.io_diffCommits_info_121_ldest; \
        force U_IF_NAME.io_diffCommits_info_121_pdest = RTL_PATH.io_diffCommits_info_121_pdest; \
        force U_IF_NAME.io_diffCommits_info_121_rfWen = RTL_PATH.io_diffCommits_info_121_rfWen; \
        force U_IF_NAME.io_diffCommits_info_121_fpWen = RTL_PATH.io_diffCommits_info_121_fpWen; \
        force U_IF_NAME.io_diffCommits_info_121_vecWen = RTL_PATH.io_diffCommits_info_121_vecWen; \
        force U_IF_NAME.io_diffCommits_info_121_v0Wen = RTL_PATH.io_diffCommits_info_121_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_121_vlWen = RTL_PATH.io_diffCommits_info_121_vlWen; \
        force U_IF_NAME.io_diffCommits_info_122_ldest = RTL_PATH.io_diffCommits_info_122_ldest; \
        force U_IF_NAME.io_diffCommits_info_122_pdest = RTL_PATH.io_diffCommits_info_122_pdest; \
        force U_IF_NAME.io_diffCommits_info_122_rfWen = RTL_PATH.io_diffCommits_info_122_rfWen; \
        force U_IF_NAME.io_diffCommits_info_122_fpWen = RTL_PATH.io_diffCommits_info_122_fpWen; \
        force U_IF_NAME.io_diffCommits_info_122_vecWen = RTL_PATH.io_diffCommits_info_122_vecWen; \
        force U_IF_NAME.io_diffCommits_info_122_v0Wen = RTL_PATH.io_diffCommits_info_122_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_122_vlWen = RTL_PATH.io_diffCommits_info_122_vlWen; \
        force U_IF_NAME.io_diffCommits_info_123_ldest = RTL_PATH.io_diffCommits_info_123_ldest; \
        force U_IF_NAME.io_diffCommits_info_123_pdest = RTL_PATH.io_diffCommits_info_123_pdest; \
        force U_IF_NAME.io_diffCommits_info_123_rfWen = RTL_PATH.io_diffCommits_info_123_rfWen; \
        force U_IF_NAME.io_diffCommits_info_123_fpWen = RTL_PATH.io_diffCommits_info_123_fpWen; \
        force U_IF_NAME.io_diffCommits_info_123_vecWen = RTL_PATH.io_diffCommits_info_123_vecWen; \
        force U_IF_NAME.io_diffCommits_info_123_v0Wen = RTL_PATH.io_diffCommits_info_123_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_123_vlWen = RTL_PATH.io_diffCommits_info_123_vlWen; \
        force U_IF_NAME.io_diffCommits_info_124_ldest = RTL_PATH.io_diffCommits_info_124_ldest; \
        force U_IF_NAME.io_diffCommits_info_124_pdest = RTL_PATH.io_diffCommits_info_124_pdest; \
        force U_IF_NAME.io_diffCommits_info_124_rfWen = RTL_PATH.io_diffCommits_info_124_rfWen; \
        force U_IF_NAME.io_diffCommits_info_124_fpWen = RTL_PATH.io_diffCommits_info_124_fpWen; \
        force U_IF_NAME.io_diffCommits_info_124_vecWen = RTL_PATH.io_diffCommits_info_124_vecWen; \
        force U_IF_NAME.io_diffCommits_info_124_v0Wen = RTL_PATH.io_diffCommits_info_124_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_124_vlWen = RTL_PATH.io_diffCommits_info_124_vlWen; \
        force U_IF_NAME.io_diffCommits_info_125_ldest = RTL_PATH.io_diffCommits_info_125_ldest; \
        force U_IF_NAME.io_diffCommits_info_125_pdest = RTL_PATH.io_diffCommits_info_125_pdest; \
        force U_IF_NAME.io_diffCommits_info_125_rfWen = RTL_PATH.io_diffCommits_info_125_rfWen; \
        force U_IF_NAME.io_diffCommits_info_125_fpWen = RTL_PATH.io_diffCommits_info_125_fpWen; \
        force U_IF_NAME.io_diffCommits_info_125_vecWen = RTL_PATH.io_diffCommits_info_125_vecWen; \
        force U_IF_NAME.io_diffCommits_info_125_v0Wen = RTL_PATH.io_diffCommits_info_125_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_125_vlWen = RTL_PATH.io_diffCommits_info_125_vlWen; \
        force U_IF_NAME.io_diffCommits_info_126_ldest = RTL_PATH.io_diffCommits_info_126_ldest; \
        force U_IF_NAME.io_diffCommits_info_126_pdest = RTL_PATH.io_diffCommits_info_126_pdest; \
        force U_IF_NAME.io_diffCommits_info_126_rfWen = RTL_PATH.io_diffCommits_info_126_rfWen; \
        force U_IF_NAME.io_diffCommits_info_126_fpWen = RTL_PATH.io_diffCommits_info_126_fpWen; \
        force U_IF_NAME.io_diffCommits_info_126_vecWen = RTL_PATH.io_diffCommits_info_126_vecWen; \
        force U_IF_NAME.io_diffCommits_info_126_v0Wen = RTL_PATH.io_diffCommits_info_126_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_126_vlWen = RTL_PATH.io_diffCommits_info_126_vlWen; \
        force U_IF_NAME.io_diffCommits_info_127_ldest = RTL_PATH.io_diffCommits_info_127_ldest; \
        force U_IF_NAME.io_diffCommits_info_127_pdest = RTL_PATH.io_diffCommits_info_127_pdest; \
        force U_IF_NAME.io_diffCommits_info_127_rfWen = RTL_PATH.io_diffCommits_info_127_rfWen; \
        force U_IF_NAME.io_diffCommits_info_127_fpWen = RTL_PATH.io_diffCommits_info_127_fpWen; \
        force U_IF_NAME.io_diffCommits_info_127_vecWen = RTL_PATH.io_diffCommits_info_127_vecWen; \
        force U_IF_NAME.io_diffCommits_info_127_v0Wen = RTL_PATH.io_diffCommits_info_127_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_127_vlWen = RTL_PATH.io_diffCommits_info_127_vlWen; \
        force U_IF_NAME.io_diffCommits_info_128_ldest = RTL_PATH.io_diffCommits_info_128_ldest; \
        force U_IF_NAME.io_diffCommits_info_128_pdest = RTL_PATH.io_diffCommits_info_128_pdest; \
        force U_IF_NAME.io_diffCommits_info_128_rfWen = RTL_PATH.io_diffCommits_info_128_rfWen; \
        force U_IF_NAME.io_diffCommits_info_128_fpWen = RTL_PATH.io_diffCommits_info_128_fpWen; \
        force U_IF_NAME.io_diffCommits_info_128_vecWen = RTL_PATH.io_diffCommits_info_128_vecWen; \
        force U_IF_NAME.io_diffCommits_info_128_v0Wen = RTL_PATH.io_diffCommits_info_128_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_128_vlWen = RTL_PATH.io_diffCommits_info_128_vlWen; \
        force U_IF_NAME.io_diffCommits_info_129_ldest = RTL_PATH.io_diffCommits_info_129_ldest; \
        force U_IF_NAME.io_diffCommits_info_129_pdest = RTL_PATH.io_diffCommits_info_129_pdest; \
        force U_IF_NAME.io_diffCommits_info_129_rfWen = RTL_PATH.io_diffCommits_info_129_rfWen; \
        force U_IF_NAME.io_diffCommits_info_129_fpWen = RTL_PATH.io_diffCommits_info_129_fpWen; \
        force U_IF_NAME.io_diffCommits_info_129_vecWen = RTL_PATH.io_diffCommits_info_129_vecWen; \
        force U_IF_NAME.io_diffCommits_info_129_v0Wen = RTL_PATH.io_diffCommits_info_129_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_129_vlWen = RTL_PATH.io_diffCommits_info_129_vlWen; \
        force U_IF_NAME.io_diffCommits_info_130_ldest = RTL_PATH.io_diffCommits_info_130_ldest; \
        force U_IF_NAME.io_diffCommits_info_130_pdest = RTL_PATH.io_diffCommits_info_130_pdest; \
        force U_IF_NAME.io_diffCommits_info_130_rfWen = RTL_PATH.io_diffCommits_info_130_rfWen; \
        force U_IF_NAME.io_diffCommits_info_130_fpWen = RTL_PATH.io_diffCommits_info_130_fpWen; \
        force U_IF_NAME.io_diffCommits_info_130_vecWen = RTL_PATH.io_diffCommits_info_130_vecWen; \
        force U_IF_NAME.io_diffCommits_info_130_v0Wen = RTL_PATH.io_diffCommits_info_130_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_130_vlWen = RTL_PATH.io_diffCommits_info_130_vlWen; \
        force U_IF_NAME.io_diffCommits_info_131_ldest = RTL_PATH.io_diffCommits_info_131_ldest; \
        force U_IF_NAME.io_diffCommits_info_131_pdest = RTL_PATH.io_diffCommits_info_131_pdest; \
        force U_IF_NAME.io_diffCommits_info_131_rfWen = RTL_PATH.io_diffCommits_info_131_rfWen; \
        force U_IF_NAME.io_diffCommits_info_131_fpWen = RTL_PATH.io_diffCommits_info_131_fpWen; \
        force U_IF_NAME.io_diffCommits_info_131_vecWen = RTL_PATH.io_diffCommits_info_131_vecWen; \
        force U_IF_NAME.io_diffCommits_info_131_v0Wen = RTL_PATH.io_diffCommits_info_131_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_131_vlWen = RTL_PATH.io_diffCommits_info_131_vlWen; \
        force U_IF_NAME.io_diffCommits_info_132_ldest = RTL_PATH.io_diffCommits_info_132_ldest; \
        force U_IF_NAME.io_diffCommits_info_132_pdest = RTL_PATH.io_diffCommits_info_132_pdest; \
        force U_IF_NAME.io_diffCommits_info_132_rfWen = RTL_PATH.io_diffCommits_info_132_rfWen; \
        force U_IF_NAME.io_diffCommits_info_132_fpWen = RTL_PATH.io_diffCommits_info_132_fpWen; \
        force U_IF_NAME.io_diffCommits_info_132_vecWen = RTL_PATH.io_diffCommits_info_132_vecWen; \
        force U_IF_NAME.io_diffCommits_info_132_v0Wen = RTL_PATH.io_diffCommits_info_132_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_132_vlWen = RTL_PATH.io_diffCommits_info_132_vlWen; \
        force U_IF_NAME.io_diffCommits_info_133_ldest = RTL_PATH.io_diffCommits_info_133_ldest; \
        force U_IF_NAME.io_diffCommits_info_133_pdest = RTL_PATH.io_diffCommits_info_133_pdest; \
        force U_IF_NAME.io_diffCommits_info_133_rfWen = RTL_PATH.io_diffCommits_info_133_rfWen; \
        force U_IF_NAME.io_diffCommits_info_133_fpWen = RTL_PATH.io_diffCommits_info_133_fpWen; \
        force U_IF_NAME.io_diffCommits_info_133_vecWen = RTL_PATH.io_diffCommits_info_133_vecWen; \
        force U_IF_NAME.io_diffCommits_info_133_v0Wen = RTL_PATH.io_diffCommits_info_133_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_133_vlWen = RTL_PATH.io_diffCommits_info_133_vlWen; \
        force U_IF_NAME.io_diffCommits_info_134_ldest = RTL_PATH.io_diffCommits_info_134_ldest; \
        force U_IF_NAME.io_diffCommits_info_134_pdest = RTL_PATH.io_diffCommits_info_134_pdest; \
        force U_IF_NAME.io_diffCommits_info_134_rfWen = RTL_PATH.io_diffCommits_info_134_rfWen; \
        force U_IF_NAME.io_diffCommits_info_134_fpWen = RTL_PATH.io_diffCommits_info_134_fpWen; \
        force U_IF_NAME.io_diffCommits_info_134_vecWen = RTL_PATH.io_diffCommits_info_134_vecWen; \
        force U_IF_NAME.io_diffCommits_info_134_v0Wen = RTL_PATH.io_diffCommits_info_134_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_134_vlWen = RTL_PATH.io_diffCommits_info_134_vlWen; \
        force U_IF_NAME.io_diffCommits_info_135_ldest = RTL_PATH.io_diffCommits_info_135_ldest; \
        force U_IF_NAME.io_diffCommits_info_135_pdest = RTL_PATH.io_diffCommits_info_135_pdest; \
        force U_IF_NAME.io_diffCommits_info_135_rfWen = RTL_PATH.io_diffCommits_info_135_rfWen; \
        force U_IF_NAME.io_diffCommits_info_135_fpWen = RTL_PATH.io_diffCommits_info_135_fpWen; \
        force U_IF_NAME.io_diffCommits_info_135_vecWen = RTL_PATH.io_diffCommits_info_135_vecWen; \
        force U_IF_NAME.io_diffCommits_info_135_v0Wen = RTL_PATH.io_diffCommits_info_135_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_135_vlWen = RTL_PATH.io_diffCommits_info_135_vlWen; \
        force U_IF_NAME.io_diffCommits_info_136_ldest = RTL_PATH.io_diffCommits_info_136_ldest; \
        force U_IF_NAME.io_diffCommits_info_136_pdest = RTL_PATH.io_diffCommits_info_136_pdest; \
        force U_IF_NAME.io_diffCommits_info_136_rfWen = RTL_PATH.io_diffCommits_info_136_rfWen; \
        force U_IF_NAME.io_diffCommits_info_136_fpWen = RTL_PATH.io_diffCommits_info_136_fpWen; \
        force U_IF_NAME.io_diffCommits_info_136_vecWen = RTL_PATH.io_diffCommits_info_136_vecWen; \
        force U_IF_NAME.io_diffCommits_info_136_v0Wen = RTL_PATH.io_diffCommits_info_136_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_136_vlWen = RTL_PATH.io_diffCommits_info_136_vlWen; \
        force U_IF_NAME.io_diffCommits_info_137_ldest = RTL_PATH.io_diffCommits_info_137_ldest; \
        force U_IF_NAME.io_diffCommits_info_137_pdest = RTL_PATH.io_diffCommits_info_137_pdest; \
        force U_IF_NAME.io_diffCommits_info_137_rfWen = RTL_PATH.io_diffCommits_info_137_rfWen; \
        force U_IF_NAME.io_diffCommits_info_137_fpWen = RTL_PATH.io_diffCommits_info_137_fpWen; \
        force U_IF_NAME.io_diffCommits_info_137_vecWen = RTL_PATH.io_diffCommits_info_137_vecWen; \
        force U_IF_NAME.io_diffCommits_info_137_v0Wen = RTL_PATH.io_diffCommits_info_137_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_137_vlWen = RTL_PATH.io_diffCommits_info_137_vlWen; \
        force U_IF_NAME.io_diffCommits_info_138_ldest = RTL_PATH.io_diffCommits_info_138_ldest; \
        force U_IF_NAME.io_diffCommits_info_138_pdest = RTL_PATH.io_diffCommits_info_138_pdest; \
        force U_IF_NAME.io_diffCommits_info_138_rfWen = RTL_PATH.io_diffCommits_info_138_rfWen; \
        force U_IF_NAME.io_diffCommits_info_138_fpWen = RTL_PATH.io_diffCommits_info_138_fpWen; \
        force U_IF_NAME.io_diffCommits_info_138_vecWen = RTL_PATH.io_diffCommits_info_138_vecWen; \
        force U_IF_NAME.io_diffCommits_info_138_v0Wen = RTL_PATH.io_diffCommits_info_138_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_138_vlWen = RTL_PATH.io_diffCommits_info_138_vlWen; \
        force U_IF_NAME.io_diffCommits_info_139_ldest = RTL_PATH.io_diffCommits_info_139_ldest; \
        force U_IF_NAME.io_diffCommits_info_139_pdest = RTL_PATH.io_diffCommits_info_139_pdest; \
        force U_IF_NAME.io_diffCommits_info_139_rfWen = RTL_PATH.io_diffCommits_info_139_rfWen; \
        force U_IF_NAME.io_diffCommits_info_139_fpWen = RTL_PATH.io_diffCommits_info_139_fpWen; \
        force U_IF_NAME.io_diffCommits_info_139_vecWen = RTL_PATH.io_diffCommits_info_139_vecWen; \
        force U_IF_NAME.io_diffCommits_info_139_v0Wen = RTL_PATH.io_diffCommits_info_139_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_139_vlWen = RTL_PATH.io_diffCommits_info_139_vlWen; \
        force U_IF_NAME.io_diffCommits_info_140_ldest = RTL_PATH.io_diffCommits_info_140_ldest; \
        force U_IF_NAME.io_diffCommits_info_140_pdest = RTL_PATH.io_diffCommits_info_140_pdest; \
        force U_IF_NAME.io_diffCommits_info_140_rfWen = RTL_PATH.io_diffCommits_info_140_rfWen; \
        force U_IF_NAME.io_diffCommits_info_140_fpWen = RTL_PATH.io_diffCommits_info_140_fpWen; \
        force U_IF_NAME.io_diffCommits_info_140_vecWen = RTL_PATH.io_diffCommits_info_140_vecWen; \
        force U_IF_NAME.io_diffCommits_info_140_v0Wen = RTL_PATH.io_diffCommits_info_140_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_140_vlWen = RTL_PATH.io_diffCommits_info_140_vlWen; \
        force U_IF_NAME.io_diffCommits_info_141_ldest = RTL_PATH.io_diffCommits_info_141_ldest; \
        force U_IF_NAME.io_diffCommits_info_141_pdest = RTL_PATH.io_diffCommits_info_141_pdest; \
        force U_IF_NAME.io_diffCommits_info_141_rfWen = RTL_PATH.io_diffCommits_info_141_rfWen; \
        force U_IF_NAME.io_diffCommits_info_141_fpWen = RTL_PATH.io_diffCommits_info_141_fpWen; \
        force U_IF_NAME.io_diffCommits_info_141_vecWen = RTL_PATH.io_diffCommits_info_141_vecWen; \
        force U_IF_NAME.io_diffCommits_info_141_v0Wen = RTL_PATH.io_diffCommits_info_141_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_141_vlWen = RTL_PATH.io_diffCommits_info_141_vlWen; \
        force U_IF_NAME.io_diffCommits_info_142_ldest = RTL_PATH.io_diffCommits_info_142_ldest; \
        force U_IF_NAME.io_diffCommits_info_142_pdest = RTL_PATH.io_diffCommits_info_142_pdest; \
        force U_IF_NAME.io_diffCommits_info_142_rfWen = RTL_PATH.io_diffCommits_info_142_rfWen; \
        force U_IF_NAME.io_diffCommits_info_142_fpWen = RTL_PATH.io_diffCommits_info_142_fpWen; \
        force U_IF_NAME.io_diffCommits_info_142_vecWen = RTL_PATH.io_diffCommits_info_142_vecWen; \
        force U_IF_NAME.io_diffCommits_info_142_v0Wen = RTL_PATH.io_diffCommits_info_142_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_142_vlWen = RTL_PATH.io_diffCommits_info_142_vlWen; \
        force U_IF_NAME.io_diffCommits_info_143_ldest = RTL_PATH.io_diffCommits_info_143_ldest; \
        force U_IF_NAME.io_diffCommits_info_143_pdest = RTL_PATH.io_diffCommits_info_143_pdest; \
        force U_IF_NAME.io_diffCommits_info_143_rfWen = RTL_PATH.io_diffCommits_info_143_rfWen; \
        force U_IF_NAME.io_diffCommits_info_143_fpWen = RTL_PATH.io_diffCommits_info_143_fpWen; \
        force U_IF_NAME.io_diffCommits_info_143_vecWen = RTL_PATH.io_diffCommits_info_143_vecWen; \
        force U_IF_NAME.io_diffCommits_info_143_v0Wen = RTL_PATH.io_diffCommits_info_143_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_143_vlWen = RTL_PATH.io_diffCommits_info_143_vlWen; \
        force U_IF_NAME.io_diffCommits_info_144_ldest = RTL_PATH.io_diffCommits_info_144_ldest; \
        force U_IF_NAME.io_diffCommits_info_144_pdest = RTL_PATH.io_diffCommits_info_144_pdest; \
        force U_IF_NAME.io_diffCommits_info_144_rfWen = RTL_PATH.io_diffCommits_info_144_rfWen; \
        force U_IF_NAME.io_diffCommits_info_144_fpWen = RTL_PATH.io_diffCommits_info_144_fpWen; \
        force U_IF_NAME.io_diffCommits_info_144_vecWen = RTL_PATH.io_diffCommits_info_144_vecWen; \
        force U_IF_NAME.io_diffCommits_info_144_v0Wen = RTL_PATH.io_diffCommits_info_144_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_144_vlWen = RTL_PATH.io_diffCommits_info_144_vlWen; \
        force U_IF_NAME.io_diffCommits_info_145_ldest = RTL_PATH.io_diffCommits_info_145_ldest; \
        force U_IF_NAME.io_diffCommits_info_145_pdest = RTL_PATH.io_diffCommits_info_145_pdest; \
        force U_IF_NAME.io_diffCommits_info_145_rfWen = RTL_PATH.io_diffCommits_info_145_rfWen; \
        force U_IF_NAME.io_diffCommits_info_145_fpWen = RTL_PATH.io_diffCommits_info_145_fpWen; \
        force U_IF_NAME.io_diffCommits_info_145_vecWen = RTL_PATH.io_diffCommits_info_145_vecWen; \
        force U_IF_NAME.io_diffCommits_info_145_v0Wen = RTL_PATH.io_diffCommits_info_145_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_145_vlWen = RTL_PATH.io_diffCommits_info_145_vlWen; \
        force U_IF_NAME.io_diffCommits_info_146_ldest = RTL_PATH.io_diffCommits_info_146_ldest; \
        force U_IF_NAME.io_diffCommits_info_146_pdest = RTL_PATH.io_diffCommits_info_146_pdest; \
        force U_IF_NAME.io_diffCommits_info_146_rfWen = RTL_PATH.io_diffCommits_info_146_rfWen; \
        force U_IF_NAME.io_diffCommits_info_146_fpWen = RTL_PATH.io_diffCommits_info_146_fpWen; \
        force U_IF_NAME.io_diffCommits_info_146_vecWen = RTL_PATH.io_diffCommits_info_146_vecWen; \
        force U_IF_NAME.io_diffCommits_info_146_v0Wen = RTL_PATH.io_diffCommits_info_146_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_146_vlWen = RTL_PATH.io_diffCommits_info_146_vlWen; \
        force U_IF_NAME.io_diffCommits_info_147_ldest = RTL_PATH.io_diffCommits_info_147_ldest; \
        force U_IF_NAME.io_diffCommits_info_147_pdest = RTL_PATH.io_diffCommits_info_147_pdest; \
        force U_IF_NAME.io_diffCommits_info_147_rfWen = RTL_PATH.io_diffCommits_info_147_rfWen; \
        force U_IF_NAME.io_diffCommits_info_147_fpWen = RTL_PATH.io_diffCommits_info_147_fpWen; \
        force U_IF_NAME.io_diffCommits_info_147_vecWen = RTL_PATH.io_diffCommits_info_147_vecWen; \
        force U_IF_NAME.io_diffCommits_info_147_v0Wen = RTL_PATH.io_diffCommits_info_147_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_147_vlWen = RTL_PATH.io_diffCommits_info_147_vlWen; \
        force U_IF_NAME.io_diffCommits_info_148_ldest = RTL_PATH.io_diffCommits_info_148_ldest; \
        force U_IF_NAME.io_diffCommits_info_148_pdest = RTL_PATH.io_diffCommits_info_148_pdest; \
        force U_IF_NAME.io_diffCommits_info_148_rfWen = RTL_PATH.io_diffCommits_info_148_rfWen; \
        force U_IF_NAME.io_diffCommits_info_148_fpWen = RTL_PATH.io_diffCommits_info_148_fpWen; \
        force U_IF_NAME.io_diffCommits_info_148_vecWen = RTL_PATH.io_diffCommits_info_148_vecWen; \
        force U_IF_NAME.io_diffCommits_info_148_v0Wen = RTL_PATH.io_diffCommits_info_148_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_148_vlWen = RTL_PATH.io_diffCommits_info_148_vlWen; \
        force U_IF_NAME.io_diffCommits_info_149_ldest = RTL_PATH.io_diffCommits_info_149_ldest; \
        force U_IF_NAME.io_diffCommits_info_149_pdest = RTL_PATH.io_diffCommits_info_149_pdest; \
        force U_IF_NAME.io_diffCommits_info_149_rfWen = RTL_PATH.io_diffCommits_info_149_rfWen; \
        force U_IF_NAME.io_diffCommits_info_149_fpWen = RTL_PATH.io_diffCommits_info_149_fpWen; \
        force U_IF_NAME.io_diffCommits_info_149_vecWen = RTL_PATH.io_diffCommits_info_149_vecWen; \
        force U_IF_NAME.io_diffCommits_info_149_v0Wen = RTL_PATH.io_diffCommits_info_149_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_149_vlWen = RTL_PATH.io_diffCommits_info_149_vlWen; \
        force U_IF_NAME.io_diffCommits_info_150_ldest = RTL_PATH.io_diffCommits_info_150_ldest; \
        force U_IF_NAME.io_diffCommits_info_150_pdest = RTL_PATH.io_diffCommits_info_150_pdest; \
        force U_IF_NAME.io_diffCommits_info_150_rfWen = RTL_PATH.io_diffCommits_info_150_rfWen; \
        force U_IF_NAME.io_diffCommits_info_150_fpWen = RTL_PATH.io_diffCommits_info_150_fpWen; \
        force U_IF_NAME.io_diffCommits_info_150_vecWen = RTL_PATH.io_diffCommits_info_150_vecWen; \
        force U_IF_NAME.io_diffCommits_info_150_v0Wen = RTL_PATH.io_diffCommits_info_150_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_150_vlWen = RTL_PATH.io_diffCommits_info_150_vlWen; \
        force U_IF_NAME.io_diffCommits_info_151_ldest = RTL_PATH.io_diffCommits_info_151_ldest; \
        force U_IF_NAME.io_diffCommits_info_151_pdest = RTL_PATH.io_diffCommits_info_151_pdest; \
        force U_IF_NAME.io_diffCommits_info_151_rfWen = RTL_PATH.io_diffCommits_info_151_rfWen; \
        force U_IF_NAME.io_diffCommits_info_151_fpWen = RTL_PATH.io_diffCommits_info_151_fpWen; \
        force U_IF_NAME.io_diffCommits_info_151_vecWen = RTL_PATH.io_diffCommits_info_151_vecWen; \
        force U_IF_NAME.io_diffCommits_info_151_v0Wen = RTL_PATH.io_diffCommits_info_151_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_151_vlWen = RTL_PATH.io_diffCommits_info_151_vlWen; \
        force U_IF_NAME.io_diffCommits_info_152_ldest = RTL_PATH.io_diffCommits_info_152_ldest; \
        force U_IF_NAME.io_diffCommits_info_152_pdest = RTL_PATH.io_diffCommits_info_152_pdest; \
        force U_IF_NAME.io_diffCommits_info_152_rfWen = RTL_PATH.io_diffCommits_info_152_rfWen; \
        force U_IF_NAME.io_diffCommits_info_152_fpWen = RTL_PATH.io_diffCommits_info_152_fpWen; \
        force U_IF_NAME.io_diffCommits_info_152_vecWen = RTL_PATH.io_diffCommits_info_152_vecWen; \
        force U_IF_NAME.io_diffCommits_info_152_v0Wen = RTL_PATH.io_diffCommits_info_152_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_152_vlWen = RTL_PATH.io_diffCommits_info_152_vlWen; \
        force U_IF_NAME.io_diffCommits_info_153_ldest = RTL_PATH.io_diffCommits_info_153_ldest; \
        force U_IF_NAME.io_diffCommits_info_153_pdest = RTL_PATH.io_diffCommits_info_153_pdest; \
        force U_IF_NAME.io_diffCommits_info_153_rfWen = RTL_PATH.io_diffCommits_info_153_rfWen; \
        force U_IF_NAME.io_diffCommits_info_153_fpWen = RTL_PATH.io_diffCommits_info_153_fpWen; \
        force U_IF_NAME.io_diffCommits_info_153_vecWen = RTL_PATH.io_diffCommits_info_153_vecWen; \
        force U_IF_NAME.io_diffCommits_info_153_v0Wen = RTL_PATH.io_diffCommits_info_153_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_153_vlWen = RTL_PATH.io_diffCommits_info_153_vlWen; \
        force U_IF_NAME.io_diffCommits_info_154_ldest = RTL_PATH.io_diffCommits_info_154_ldest; \
        force U_IF_NAME.io_diffCommits_info_154_pdest = RTL_PATH.io_diffCommits_info_154_pdest; \
        force U_IF_NAME.io_diffCommits_info_154_rfWen = RTL_PATH.io_diffCommits_info_154_rfWen; \
        force U_IF_NAME.io_diffCommits_info_154_fpWen = RTL_PATH.io_diffCommits_info_154_fpWen; \
        force U_IF_NAME.io_diffCommits_info_154_vecWen = RTL_PATH.io_diffCommits_info_154_vecWen; \
        force U_IF_NAME.io_diffCommits_info_154_v0Wen = RTL_PATH.io_diffCommits_info_154_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_154_vlWen = RTL_PATH.io_diffCommits_info_154_vlWen; \
        force U_IF_NAME.io_diffCommits_info_155_ldest = RTL_PATH.io_diffCommits_info_155_ldest; \
        force U_IF_NAME.io_diffCommits_info_155_pdest = RTL_PATH.io_diffCommits_info_155_pdest; \
        force U_IF_NAME.io_diffCommits_info_155_rfWen = RTL_PATH.io_diffCommits_info_155_rfWen; \
        force U_IF_NAME.io_diffCommits_info_155_fpWen = RTL_PATH.io_diffCommits_info_155_fpWen; \
        force U_IF_NAME.io_diffCommits_info_155_vecWen = RTL_PATH.io_diffCommits_info_155_vecWen; \
        force U_IF_NAME.io_diffCommits_info_155_v0Wen = RTL_PATH.io_diffCommits_info_155_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_155_vlWen = RTL_PATH.io_diffCommits_info_155_vlWen; \
        force U_IF_NAME.io_diffCommits_info_156_ldest = RTL_PATH.io_diffCommits_info_156_ldest; \
        force U_IF_NAME.io_diffCommits_info_156_pdest = RTL_PATH.io_diffCommits_info_156_pdest; \
        force U_IF_NAME.io_diffCommits_info_156_rfWen = RTL_PATH.io_diffCommits_info_156_rfWen; \
        force U_IF_NAME.io_diffCommits_info_156_fpWen = RTL_PATH.io_diffCommits_info_156_fpWen; \
        force U_IF_NAME.io_diffCommits_info_156_vecWen = RTL_PATH.io_diffCommits_info_156_vecWen; \
        force U_IF_NAME.io_diffCommits_info_156_v0Wen = RTL_PATH.io_diffCommits_info_156_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_156_vlWen = RTL_PATH.io_diffCommits_info_156_vlWen; \
        force U_IF_NAME.io_diffCommits_info_157_ldest = RTL_PATH.io_diffCommits_info_157_ldest; \
        force U_IF_NAME.io_diffCommits_info_157_pdest = RTL_PATH.io_diffCommits_info_157_pdest; \
        force U_IF_NAME.io_diffCommits_info_157_rfWen = RTL_PATH.io_diffCommits_info_157_rfWen; \
        force U_IF_NAME.io_diffCommits_info_157_fpWen = RTL_PATH.io_diffCommits_info_157_fpWen; \
        force U_IF_NAME.io_diffCommits_info_157_vecWen = RTL_PATH.io_diffCommits_info_157_vecWen; \
        force U_IF_NAME.io_diffCommits_info_157_v0Wen = RTL_PATH.io_diffCommits_info_157_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_157_vlWen = RTL_PATH.io_diffCommits_info_157_vlWen; \
        force U_IF_NAME.io_diffCommits_info_158_ldest = RTL_PATH.io_diffCommits_info_158_ldest; \
        force U_IF_NAME.io_diffCommits_info_158_pdest = RTL_PATH.io_diffCommits_info_158_pdest; \
        force U_IF_NAME.io_diffCommits_info_158_rfWen = RTL_PATH.io_diffCommits_info_158_rfWen; \
        force U_IF_NAME.io_diffCommits_info_158_fpWen = RTL_PATH.io_diffCommits_info_158_fpWen; \
        force U_IF_NAME.io_diffCommits_info_158_vecWen = RTL_PATH.io_diffCommits_info_158_vecWen; \
        force U_IF_NAME.io_diffCommits_info_158_v0Wen = RTL_PATH.io_diffCommits_info_158_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_158_vlWen = RTL_PATH.io_diffCommits_info_158_vlWen; \
        force U_IF_NAME.io_diffCommits_info_159_ldest = RTL_PATH.io_diffCommits_info_159_ldest; \
        force U_IF_NAME.io_diffCommits_info_159_pdest = RTL_PATH.io_diffCommits_info_159_pdest; \
        force U_IF_NAME.io_diffCommits_info_159_rfWen = RTL_PATH.io_diffCommits_info_159_rfWen; \
        force U_IF_NAME.io_diffCommits_info_159_fpWen = RTL_PATH.io_diffCommits_info_159_fpWen; \
        force U_IF_NAME.io_diffCommits_info_159_vecWen = RTL_PATH.io_diffCommits_info_159_vecWen; \
        force U_IF_NAME.io_diffCommits_info_159_v0Wen = RTL_PATH.io_diffCommits_info_159_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_159_vlWen = RTL_PATH.io_diffCommits_info_159_vlWen; \
        force U_IF_NAME.io_diffCommits_info_160_ldest = RTL_PATH.io_diffCommits_info_160_ldest; \
        force U_IF_NAME.io_diffCommits_info_160_pdest = RTL_PATH.io_diffCommits_info_160_pdest; \
        force U_IF_NAME.io_diffCommits_info_160_rfWen = RTL_PATH.io_diffCommits_info_160_rfWen; \
        force U_IF_NAME.io_diffCommits_info_160_fpWen = RTL_PATH.io_diffCommits_info_160_fpWen; \
        force U_IF_NAME.io_diffCommits_info_160_vecWen = RTL_PATH.io_diffCommits_info_160_vecWen; \
        force U_IF_NAME.io_diffCommits_info_160_v0Wen = RTL_PATH.io_diffCommits_info_160_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_160_vlWen = RTL_PATH.io_diffCommits_info_160_vlWen; \
        force U_IF_NAME.io_diffCommits_info_161_ldest = RTL_PATH.io_diffCommits_info_161_ldest; \
        force U_IF_NAME.io_diffCommits_info_161_pdest = RTL_PATH.io_diffCommits_info_161_pdest; \
        force U_IF_NAME.io_diffCommits_info_161_rfWen = RTL_PATH.io_diffCommits_info_161_rfWen; \
        force U_IF_NAME.io_diffCommits_info_161_fpWen = RTL_PATH.io_diffCommits_info_161_fpWen; \
        force U_IF_NAME.io_diffCommits_info_161_vecWen = RTL_PATH.io_diffCommits_info_161_vecWen; \
        force U_IF_NAME.io_diffCommits_info_161_v0Wen = RTL_PATH.io_diffCommits_info_161_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_161_vlWen = RTL_PATH.io_diffCommits_info_161_vlWen; \
        force U_IF_NAME.io_diffCommits_info_162_ldest = RTL_PATH.io_diffCommits_info_162_ldest; \
        force U_IF_NAME.io_diffCommits_info_162_pdest = RTL_PATH.io_diffCommits_info_162_pdest; \
        force U_IF_NAME.io_diffCommits_info_162_rfWen = RTL_PATH.io_diffCommits_info_162_rfWen; \
        force U_IF_NAME.io_diffCommits_info_162_fpWen = RTL_PATH.io_diffCommits_info_162_fpWen; \
        force U_IF_NAME.io_diffCommits_info_162_vecWen = RTL_PATH.io_diffCommits_info_162_vecWen; \
        force U_IF_NAME.io_diffCommits_info_162_v0Wen = RTL_PATH.io_diffCommits_info_162_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_162_vlWen = RTL_PATH.io_diffCommits_info_162_vlWen; \
        force U_IF_NAME.io_diffCommits_info_163_ldest = RTL_PATH.io_diffCommits_info_163_ldest; \
        force U_IF_NAME.io_diffCommits_info_163_pdest = RTL_PATH.io_diffCommits_info_163_pdest; \
        force U_IF_NAME.io_diffCommits_info_163_rfWen = RTL_PATH.io_diffCommits_info_163_rfWen; \
        force U_IF_NAME.io_diffCommits_info_163_fpWen = RTL_PATH.io_diffCommits_info_163_fpWen; \
        force U_IF_NAME.io_diffCommits_info_163_vecWen = RTL_PATH.io_diffCommits_info_163_vecWen; \
        force U_IF_NAME.io_diffCommits_info_163_v0Wen = RTL_PATH.io_diffCommits_info_163_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_163_vlWen = RTL_PATH.io_diffCommits_info_163_vlWen; \
        force U_IF_NAME.io_diffCommits_info_164_ldest = RTL_PATH.io_diffCommits_info_164_ldest; \
        force U_IF_NAME.io_diffCommits_info_164_pdest = RTL_PATH.io_diffCommits_info_164_pdest; \
        force U_IF_NAME.io_diffCommits_info_164_rfWen = RTL_PATH.io_diffCommits_info_164_rfWen; \
        force U_IF_NAME.io_diffCommits_info_164_fpWen = RTL_PATH.io_diffCommits_info_164_fpWen; \
        force U_IF_NAME.io_diffCommits_info_164_vecWen = RTL_PATH.io_diffCommits_info_164_vecWen; \
        force U_IF_NAME.io_diffCommits_info_164_v0Wen = RTL_PATH.io_diffCommits_info_164_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_164_vlWen = RTL_PATH.io_diffCommits_info_164_vlWen; \
        force U_IF_NAME.io_diffCommits_info_165_ldest = RTL_PATH.io_diffCommits_info_165_ldest; \
        force U_IF_NAME.io_diffCommits_info_165_pdest = RTL_PATH.io_diffCommits_info_165_pdest; \
        force U_IF_NAME.io_diffCommits_info_165_rfWen = RTL_PATH.io_diffCommits_info_165_rfWen; \
        force U_IF_NAME.io_diffCommits_info_165_fpWen = RTL_PATH.io_diffCommits_info_165_fpWen; \
        force U_IF_NAME.io_diffCommits_info_165_vecWen = RTL_PATH.io_diffCommits_info_165_vecWen; \
        force U_IF_NAME.io_diffCommits_info_165_v0Wen = RTL_PATH.io_diffCommits_info_165_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_165_vlWen = RTL_PATH.io_diffCommits_info_165_vlWen; \
        force U_IF_NAME.io_diffCommits_info_166_ldest = RTL_PATH.io_diffCommits_info_166_ldest; \
        force U_IF_NAME.io_diffCommits_info_166_pdest = RTL_PATH.io_diffCommits_info_166_pdest; \
        force U_IF_NAME.io_diffCommits_info_166_rfWen = RTL_PATH.io_diffCommits_info_166_rfWen; \
        force U_IF_NAME.io_diffCommits_info_166_fpWen = RTL_PATH.io_diffCommits_info_166_fpWen; \
        force U_IF_NAME.io_diffCommits_info_166_vecWen = RTL_PATH.io_diffCommits_info_166_vecWen; \
        force U_IF_NAME.io_diffCommits_info_166_v0Wen = RTL_PATH.io_diffCommits_info_166_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_166_vlWen = RTL_PATH.io_diffCommits_info_166_vlWen; \
        force U_IF_NAME.io_diffCommits_info_167_ldest = RTL_PATH.io_diffCommits_info_167_ldest; \
        force U_IF_NAME.io_diffCommits_info_167_pdest = RTL_PATH.io_diffCommits_info_167_pdest; \
        force U_IF_NAME.io_diffCommits_info_167_rfWen = RTL_PATH.io_diffCommits_info_167_rfWen; \
        force U_IF_NAME.io_diffCommits_info_167_fpWen = RTL_PATH.io_diffCommits_info_167_fpWen; \
        force U_IF_NAME.io_diffCommits_info_167_vecWen = RTL_PATH.io_diffCommits_info_167_vecWen; \
        force U_IF_NAME.io_diffCommits_info_167_v0Wen = RTL_PATH.io_diffCommits_info_167_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_167_vlWen = RTL_PATH.io_diffCommits_info_167_vlWen; \
        force U_IF_NAME.io_diffCommits_info_168_ldest = RTL_PATH.io_diffCommits_info_168_ldest; \
        force U_IF_NAME.io_diffCommits_info_168_pdest = RTL_PATH.io_diffCommits_info_168_pdest; \
        force U_IF_NAME.io_diffCommits_info_168_rfWen = RTL_PATH.io_diffCommits_info_168_rfWen; \
        force U_IF_NAME.io_diffCommits_info_168_fpWen = RTL_PATH.io_diffCommits_info_168_fpWen; \
        force U_IF_NAME.io_diffCommits_info_168_vecWen = RTL_PATH.io_diffCommits_info_168_vecWen; \
        force U_IF_NAME.io_diffCommits_info_168_v0Wen = RTL_PATH.io_diffCommits_info_168_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_168_vlWen = RTL_PATH.io_diffCommits_info_168_vlWen; \
        force U_IF_NAME.io_diffCommits_info_169_ldest = RTL_PATH.io_diffCommits_info_169_ldest; \
        force U_IF_NAME.io_diffCommits_info_169_pdest = RTL_PATH.io_diffCommits_info_169_pdest; \
        force U_IF_NAME.io_diffCommits_info_169_rfWen = RTL_PATH.io_diffCommits_info_169_rfWen; \
        force U_IF_NAME.io_diffCommits_info_169_fpWen = RTL_PATH.io_diffCommits_info_169_fpWen; \
        force U_IF_NAME.io_diffCommits_info_169_vecWen = RTL_PATH.io_diffCommits_info_169_vecWen; \
        force U_IF_NAME.io_diffCommits_info_169_v0Wen = RTL_PATH.io_diffCommits_info_169_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_169_vlWen = RTL_PATH.io_diffCommits_info_169_vlWen; \
        force U_IF_NAME.io_diffCommits_info_170_ldest = RTL_PATH.io_diffCommits_info_170_ldest; \
        force U_IF_NAME.io_diffCommits_info_170_pdest = RTL_PATH.io_diffCommits_info_170_pdest; \
        force U_IF_NAME.io_diffCommits_info_170_rfWen = RTL_PATH.io_diffCommits_info_170_rfWen; \
        force U_IF_NAME.io_diffCommits_info_170_fpWen = RTL_PATH.io_diffCommits_info_170_fpWen; \
        force U_IF_NAME.io_diffCommits_info_170_vecWen = RTL_PATH.io_diffCommits_info_170_vecWen; \
        force U_IF_NAME.io_diffCommits_info_170_v0Wen = RTL_PATH.io_diffCommits_info_170_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_170_vlWen = RTL_PATH.io_diffCommits_info_170_vlWen; \
        force U_IF_NAME.io_diffCommits_info_171_ldest = RTL_PATH.io_diffCommits_info_171_ldest; \
        force U_IF_NAME.io_diffCommits_info_171_pdest = RTL_PATH.io_diffCommits_info_171_pdest; \
        force U_IF_NAME.io_diffCommits_info_171_rfWen = RTL_PATH.io_diffCommits_info_171_rfWen; \
        force U_IF_NAME.io_diffCommits_info_171_fpWen = RTL_PATH.io_diffCommits_info_171_fpWen; \
        force U_IF_NAME.io_diffCommits_info_171_vecWen = RTL_PATH.io_diffCommits_info_171_vecWen; \
        force U_IF_NAME.io_diffCommits_info_171_v0Wen = RTL_PATH.io_diffCommits_info_171_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_171_vlWen = RTL_PATH.io_diffCommits_info_171_vlWen; \
        force U_IF_NAME.io_diffCommits_info_172_ldest = RTL_PATH.io_diffCommits_info_172_ldest; \
        force U_IF_NAME.io_diffCommits_info_172_pdest = RTL_PATH.io_diffCommits_info_172_pdest; \
        force U_IF_NAME.io_diffCommits_info_172_rfWen = RTL_PATH.io_diffCommits_info_172_rfWen; \
        force U_IF_NAME.io_diffCommits_info_172_fpWen = RTL_PATH.io_diffCommits_info_172_fpWen; \
        force U_IF_NAME.io_diffCommits_info_172_vecWen = RTL_PATH.io_diffCommits_info_172_vecWen; \
        force U_IF_NAME.io_diffCommits_info_172_v0Wen = RTL_PATH.io_diffCommits_info_172_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_172_vlWen = RTL_PATH.io_diffCommits_info_172_vlWen; \
        force U_IF_NAME.io_diffCommits_info_173_ldest = RTL_PATH.io_diffCommits_info_173_ldest; \
        force U_IF_NAME.io_diffCommits_info_173_pdest = RTL_PATH.io_diffCommits_info_173_pdest; \
        force U_IF_NAME.io_diffCommits_info_173_rfWen = RTL_PATH.io_diffCommits_info_173_rfWen; \
        force U_IF_NAME.io_diffCommits_info_173_fpWen = RTL_PATH.io_diffCommits_info_173_fpWen; \
        force U_IF_NAME.io_diffCommits_info_173_vecWen = RTL_PATH.io_diffCommits_info_173_vecWen; \
        force U_IF_NAME.io_diffCommits_info_173_v0Wen = RTL_PATH.io_diffCommits_info_173_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_173_vlWen = RTL_PATH.io_diffCommits_info_173_vlWen; \
        force U_IF_NAME.io_diffCommits_info_174_ldest = RTL_PATH.io_diffCommits_info_174_ldest; \
        force U_IF_NAME.io_diffCommits_info_174_pdest = RTL_PATH.io_diffCommits_info_174_pdest; \
        force U_IF_NAME.io_diffCommits_info_174_rfWen = RTL_PATH.io_diffCommits_info_174_rfWen; \
        force U_IF_NAME.io_diffCommits_info_174_fpWen = RTL_PATH.io_diffCommits_info_174_fpWen; \
        force U_IF_NAME.io_diffCommits_info_174_vecWen = RTL_PATH.io_diffCommits_info_174_vecWen; \
        force U_IF_NAME.io_diffCommits_info_174_v0Wen = RTL_PATH.io_diffCommits_info_174_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_174_vlWen = RTL_PATH.io_diffCommits_info_174_vlWen; \
        force U_IF_NAME.io_diffCommits_info_175_ldest = RTL_PATH.io_diffCommits_info_175_ldest; \
        force U_IF_NAME.io_diffCommits_info_175_pdest = RTL_PATH.io_diffCommits_info_175_pdest; \
        force U_IF_NAME.io_diffCommits_info_175_rfWen = RTL_PATH.io_diffCommits_info_175_rfWen; \
        force U_IF_NAME.io_diffCommits_info_175_fpWen = RTL_PATH.io_diffCommits_info_175_fpWen; \
        force U_IF_NAME.io_diffCommits_info_175_vecWen = RTL_PATH.io_diffCommits_info_175_vecWen; \
        force U_IF_NAME.io_diffCommits_info_175_v0Wen = RTL_PATH.io_diffCommits_info_175_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_175_vlWen = RTL_PATH.io_diffCommits_info_175_vlWen; \
        force U_IF_NAME.io_diffCommits_info_176_ldest = RTL_PATH.io_diffCommits_info_176_ldest; \
        force U_IF_NAME.io_diffCommits_info_176_pdest = RTL_PATH.io_diffCommits_info_176_pdest; \
        force U_IF_NAME.io_diffCommits_info_176_rfWen = RTL_PATH.io_diffCommits_info_176_rfWen; \
        force U_IF_NAME.io_diffCommits_info_176_fpWen = RTL_PATH.io_diffCommits_info_176_fpWen; \
        force U_IF_NAME.io_diffCommits_info_176_vecWen = RTL_PATH.io_diffCommits_info_176_vecWen; \
        force U_IF_NAME.io_diffCommits_info_176_v0Wen = RTL_PATH.io_diffCommits_info_176_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_176_vlWen = RTL_PATH.io_diffCommits_info_176_vlWen; \
        force U_IF_NAME.io_diffCommits_info_177_ldest = RTL_PATH.io_diffCommits_info_177_ldest; \
        force U_IF_NAME.io_diffCommits_info_177_pdest = RTL_PATH.io_diffCommits_info_177_pdest; \
        force U_IF_NAME.io_diffCommits_info_177_rfWen = RTL_PATH.io_diffCommits_info_177_rfWen; \
        force U_IF_NAME.io_diffCommits_info_177_fpWen = RTL_PATH.io_diffCommits_info_177_fpWen; \
        force U_IF_NAME.io_diffCommits_info_177_vecWen = RTL_PATH.io_diffCommits_info_177_vecWen; \
        force U_IF_NAME.io_diffCommits_info_177_v0Wen = RTL_PATH.io_diffCommits_info_177_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_177_vlWen = RTL_PATH.io_diffCommits_info_177_vlWen; \
        force U_IF_NAME.io_diffCommits_info_178_ldest = RTL_PATH.io_diffCommits_info_178_ldest; \
        force U_IF_NAME.io_diffCommits_info_178_pdest = RTL_PATH.io_diffCommits_info_178_pdest; \
        force U_IF_NAME.io_diffCommits_info_178_rfWen = RTL_PATH.io_diffCommits_info_178_rfWen; \
        force U_IF_NAME.io_diffCommits_info_178_fpWen = RTL_PATH.io_diffCommits_info_178_fpWen; \
        force U_IF_NAME.io_diffCommits_info_178_vecWen = RTL_PATH.io_diffCommits_info_178_vecWen; \
        force U_IF_NAME.io_diffCommits_info_178_v0Wen = RTL_PATH.io_diffCommits_info_178_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_178_vlWen = RTL_PATH.io_diffCommits_info_178_vlWen; \
        force U_IF_NAME.io_diffCommits_info_179_ldest = RTL_PATH.io_diffCommits_info_179_ldest; \
        force U_IF_NAME.io_diffCommits_info_179_pdest = RTL_PATH.io_diffCommits_info_179_pdest; \
        force U_IF_NAME.io_diffCommits_info_179_rfWen = RTL_PATH.io_diffCommits_info_179_rfWen; \
        force U_IF_NAME.io_diffCommits_info_179_fpWen = RTL_PATH.io_diffCommits_info_179_fpWen; \
        force U_IF_NAME.io_diffCommits_info_179_vecWen = RTL_PATH.io_diffCommits_info_179_vecWen; \
        force U_IF_NAME.io_diffCommits_info_179_v0Wen = RTL_PATH.io_diffCommits_info_179_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_179_vlWen = RTL_PATH.io_diffCommits_info_179_vlWen; \
        force U_IF_NAME.io_diffCommits_info_180_ldest = RTL_PATH.io_diffCommits_info_180_ldest; \
        force U_IF_NAME.io_diffCommits_info_180_pdest = RTL_PATH.io_diffCommits_info_180_pdest; \
        force U_IF_NAME.io_diffCommits_info_180_rfWen = RTL_PATH.io_diffCommits_info_180_rfWen; \
        force U_IF_NAME.io_diffCommits_info_180_fpWen = RTL_PATH.io_diffCommits_info_180_fpWen; \
        force U_IF_NAME.io_diffCommits_info_180_vecWen = RTL_PATH.io_diffCommits_info_180_vecWen; \
        force U_IF_NAME.io_diffCommits_info_180_v0Wen = RTL_PATH.io_diffCommits_info_180_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_180_vlWen = RTL_PATH.io_diffCommits_info_180_vlWen; \
        force U_IF_NAME.io_diffCommits_info_181_ldest = RTL_PATH.io_diffCommits_info_181_ldest; \
        force U_IF_NAME.io_diffCommits_info_181_pdest = RTL_PATH.io_diffCommits_info_181_pdest; \
        force U_IF_NAME.io_diffCommits_info_181_rfWen = RTL_PATH.io_diffCommits_info_181_rfWen; \
        force U_IF_NAME.io_diffCommits_info_181_fpWen = RTL_PATH.io_diffCommits_info_181_fpWen; \
        force U_IF_NAME.io_diffCommits_info_181_vecWen = RTL_PATH.io_diffCommits_info_181_vecWen; \
        force U_IF_NAME.io_diffCommits_info_181_v0Wen = RTL_PATH.io_diffCommits_info_181_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_181_vlWen = RTL_PATH.io_diffCommits_info_181_vlWen; \
        force U_IF_NAME.io_diffCommits_info_182_ldest = RTL_PATH.io_diffCommits_info_182_ldest; \
        force U_IF_NAME.io_diffCommits_info_182_pdest = RTL_PATH.io_diffCommits_info_182_pdest; \
        force U_IF_NAME.io_diffCommits_info_182_rfWen = RTL_PATH.io_diffCommits_info_182_rfWen; \
        force U_IF_NAME.io_diffCommits_info_182_fpWen = RTL_PATH.io_diffCommits_info_182_fpWen; \
        force U_IF_NAME.io_diffCommits_info_182_vecWen = RTL_PATH.io_diffCommits_info_182_vecWen; \
        force U_IF_NAME.io_diffCommits_info_182_v0Wen = RTL_PATH.io_diffCommits_info_182_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_182_vlWen = RTL_PATH.io_diffCommits_info_182_vlWen; \
        force U_IF_NAME.io_diffCommits_info_183_ldest = RTL_PATH.io_diffCommits_info_183_ldest; \
        force U_IF_NAME.io_diffCommits_info_183_pdest = RTL_PATH.io_diffCommits_info_183_pdest; \
        force U_IF_NAME.io_diffCommits_info_183_rfWen = RTL_PATH.io_diffCommits_info_183_rfWen; \
        force U_IF_NAME.io_diffCommits_info_183_fpWen = RTL_PATH.io_diffCommits_info_183_fpWen; \
        force U_IF_NAME.io_diffCommits_info_183_vecWen = RTL_PATH.io_diffCommits_info_183_vecWen; \
        force U_IF_NAME.io_diffCommits_info_183_v0Wen = RTL_PATH.io_diffCommits_info_183_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_183_vlWen = RTL_PATH.io_diffCommits_info_183_vlWen; \
        force U_IF_NAME.io_diffCommits_info_184_ldest = RTL_PATH.io_diffCommits_info_184_ldest; \
        force U_IF_NAME.io_diffCommits_info_184_pdest = RTL_PATH.io_diffCommits_info_184_pdest; \
        force U_IF_NAME.io_diffCommits_info_184_rfWen = RTL_PATH.io_diffCommits_info_184_rfWen; \
        force U_IF_NAME.io_diffCommits_info_184_fpWen = RTL_PATH.io_diffCommits_info_184_fpWen; \
        force U_IF_NAME.io_diffCommits_info_184_vecWen = RTL_PATH.io_diffCommits_info_184_vecWen; \
        force U_IF_NAME.io_diffCommits_info_184_v0Wen = RTL_PATH.io_diffCommits_info_184_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_184_vlWen = RTL_PATH.io_diffCommits_info_184_vlWen; \
        force U_IF_NAME.io_diffCommits_info_185_ldest = RTL_PATH.io_diffCommits_info_185_ldest; \
        force U_IF_NAME.io_diffCommits_info_185_pdest = RTL_PATH.io_diffCommits_info_185_pdest; \
        force U_IF_NAME.io_diffCommits_info_185_rfWen = RTL_PATH.io_diffCommits_info_185_rfWen; \
        force U_IF_NAME.io_diffCommits_info_185_fpWen = RTL_PATH.io_diffCommits_info_185_fpWen; \
        force U_IF_NAME.io_diffCommits_info_185_vecWen = RTL_PATH.io_diffCommits_info_185_vecWen; \
        force U_IF_NAME.io_diffCommits_info_185_v0Wen = RTL_PATH.io_diffCommits_info_185_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_185_vlWen = RTL_PATH.io_diffCommits_info_185_vlWen; \
        force U_IF_NAME.io_diffCommits_info_186_ldest = RTL_PATH.io_diffCommits_info_186_ldest; \
        force U_IF_NAME.io_diffCommits_info_186_pdest = RTL_PATH.io_diffCommits_info_186_pdest; \
        force U_IF_NAME.io_diffCommits_info_186_rfWen = RTL_PATH.io_diffCommits_info_186_rfWen; \
        force U_IF_NAME.io_diffCommits_info_186_fpWen = RTL_PATH.io_diffCommits_info_186_fpWen; \
        force U_IF_NAME.io_diffCommits_info_186_vecWen = RTL_PATH.io_diffCommits_info_186_vecWen; \
        force U_IF_NAME.io_diffCommits_info_186_v0Wen = RTL_PATH.io_diffCommits_info_186_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_186_vlWen = RTL_PATH.io_diffCommits_info_186_vlWen; \
        force U_IF_NAME.io_diffCommits_info_187_ldest = RTL_PATH.io_diffCommits_info_187_ldest; \
        force U_IF_NAME.io_diffCommits_info_187_pdest = RTL_PATH.io_diffCommits_info_187_pdest; \
        force U_IF_NAME.io_diffCommits_info_187_rfWen = RTL_PATH.io_diffCommits_info_187_rfWen; \
        force U_IF_NAME.io_diffCommits_info_187_fpWen = RTL_PATH.io_diffCommits_info_187_fpWen; \
        force U_IF_NAME.io_diffCommits_info_187_vecWen = RTL_PATH.io_diffCommits_info_187_vecWen; \
        force U_IF_NAME.io_diffCommits_info_187_v0Wen = RTL_PATH.io_diffCommits_info_187_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_187_vlWen = RTL_PATH.io_diffCommits_info_187_vlWen; \
        force U_IF_NAME.io_diffCommits_info_188_ldest = RTL_PATH.io_diffCommits_info_188_ldest; \
        force U_IF_NAME.io_diffCommits_info_188_pdest = RTL_PATH.io_diffCommits_info_188_pdest; \
        force U_IF_NAME.io_diffCommits_info_188_rfWen = RTL_PATH.io_diffCommits_info_188_rfWen; \
        force U_IF_NAME.io_diffCommits_info_188_fpWen = RTL_PATH.io_diffCommits_info_188_fpWen; \
        force U_IF_NAME.io_diffCommits_info_188_vecWen = RTL_PATH.io_diffCommits_info_188_vecWen; \
        force U_IF_NAME.io_diffCommits_info_188_v0Wen = RTL_PATH.io_diffCommits_info_188_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_188_vlWen = RTL_PATH.io_diffCommits_info_188_vlWen; \
        force U_IF_NAME.io_diffCommits_info_189_ldest = RTL_PATH.io_diffCommits_info_189_ldest; \
        force U_IF_NAME.io_diffCommits_info_189_pdest = RTL_PATH.io_diffCommits_info_189_pdest; \
        force U_IF_NAME.io_diffCommits_info_189_rfWen = RTL_PATH.io_diffCommits_info_189_rfWen; \
        force U_IF_NAME.io_diffCommits_info_189_fpWen = RTL_PATH.io_diffCommits_info_189_fpWen; \
        force U_IF_NAME.io_diffCommits_info_189_vecWen = RTL_PATH.io_diffCommits_info_189_vecWen; \
        force U_IF_NAME.io_diffCommits_info_189_v0Wen = RTL_PATH.io_diffCommits_info_189_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_189_vlWen = RTL_PATH.io_diffCommits_info_189_vlWen; \
        force U_IF_NAME.io_diffCommits_info_190_ldest = RTL_PATH.io_diffCommits_info_190_ldest; \
        force U_IF_NAME.io_diffCommits_info_190_pdest = RTL_PATH.io_diffCommits_info_190_pdest; \
        force U_IF_NAME.io_diffCommits_info_190_rfWen = RTL_PATH.io_diffCommits_info_190_rfWen; \
        force U_IF_NAME.io_diffCommits_info_190_fpWen = RTL_PATH.io_diffCommits_info_190_fpWen; \
        force U_IF_NAME.io_diffCommits_info_190_vecWen = RTL_PATH.io_diffCommits_info_190_vecWen; \
        force U_IF_NAME.io_diffCommits_info_190_v0Wen = RTL_PATH.io_diffCommits_info_190_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_190_vlWen = RTL_PATH.io_diffCommits_info_190_vlWen; \
        force U_IF_NAME.io_diffCommits_info_191_ldest = RTL_PATH.io_diffCommits_info_191_ldest; \
        force U_IF_NAME.io_diffCommits_info_191_pdest = RTL_PATH.io_diffCommits_info_191_pdest; \
        force U_IF_NAME.io_diffCommits_info_191_rfWen = RTL_PATH.io_diffCommits_info_191_rfWen; \
        force U_IF_NAME.io_diffCommits_info_191_fpWen = RTL_PATH.io_diffCommits_info_191_fpWen; \
        force U_IF_NAME.io_diffCommits_info_191_vecWen = RTL_PATH.io_diffCommits_info_191_vecWen; \
        force U_IF_NAME.io_diffCommits_info_191_v0Wen = RTL_PATH.io_diffCommits_info_191_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_191_vlWen = RTL_PATH.io_diffCommits_info_191_vlWen; \
        force U_IF_NAME.io_diffCommits_info_192_ldest = RTL_PATH.io_diffCommits_info_192_ldest; \
        force U_IF_NAME.io_diffCommits_info_192_pdest = RTL_PATH.io_diffCommits_info_192_pdest; \
        force U_IF_NAME.io_diffCommits_info_192_rfWen = RTL_PATH.io_diffCommits_info_192_rfWen; \
        force U_IF_NAME.io_diffCommits_info_192_fpWen = RTL_PATH.io_diffCommits_info_192_fpWen; \
        force U_IF_NAME.io_diffCommits_info_192_vecWen = RTL_PATH.io_diffCommits_info_192_vecWen; \
        force U_IF_NAME.io_diffCommits_info_192_v0Wen = RTL_PATH.io_diffCommits_info_192_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_192_vlWen = RTL_PATH.io_diffCommits_info_192_vlWen; \
        force U_IF_NAME.io_diffCommits_info_193_ldest = RTL_PATH.io_diffCommits_info_193_ldest; \
        force U_IF_NAME.io_diffCommits_info_193_pdest = RTL_PATH.io_diffCommits_info_193_pdest; \
        force U_IF_NAME.io_diffCommits_info_193_rfWen = RTL_PATH.io_diffCommits_info_193_rfWen; \
        force U_IF_NAME.io_diffCommits_info_193_fpWen = RTL_PATH.io_diffCommits_info_193_fpWen; \
        force U_IF_NAME.io_diffCommits_info_193_vecWen = RTL_PATH.io_diffCommits_info_193_vecWen; \
        force U_IF_NAME.io_diffCommits_info_193_v0Wen = RTL_PATH.io_diffCommits_info_193_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_193_vlWen = RTL_PATH.io_diffCommits_info_193_vlWen; \
        force U_IF_NAME.io_diffCommits_info_194_ldest = RTL_PATH.io_diffCommits_info_194_ldest; \
        force U_IF_NAME.io_diffCommits_info_194_pdest = RTL_PATH.io_diffCommits_info_194_pdest; \
        force U_IF_NAME.io_diffCommits_info_194_rfWen = RTL_PATH.io_diffCommits_info_194_rfWen; \
        force U_IF_NAME.io_diffCommits_info_194_fpWen = RTL_PATH.io_diffCommits_info_194_fpWen; \
        force U_IF_NAME.io_diffCommits_info_194_vecWen = RTL_PATH.io_diffCommits_info_194_vecWen; \
        force U_IF_NAME.io_diffCommits_info_194_v0Wen = RTL_PATH.io_diffCommits_info_194_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_194_vlWen = RTL_PATH.io_diffCommits_info_194_vlWen; \
        force U_IF_NAME.io_diffCommits_info_195_ldest = RTL_PATH.io_diffCommits_info_195_ldest; \
        force U_IF_NAME.io_diffCommits_info_195_pdest = RTL_PATH.io_diffCommits_info_195_pdest; \
        force U_IF_NAME.io_diffCommits_info_195_rfWen = RTL_PATH.io_diffCommits_info_195_rfWen; \
        force U_IF_NAME.io_diffCommits_info_195_fpWen = RTL_PATH.io_diffCommits_info_195_fpWen; \
        force U_IF_NAME.io_diffCommits_info_195_vecWen = RTL_PATH.io_diffCommits_info_195_vecWen; \
        force U_IF_NAME.io_diffCommits_info_195_v0Wen = RTL_PATH.io_diffCommits_info_195_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_195_vlWen = RTL_PATH.io_diffCommits_info_195_vlWen; \
        force U_IF_NAME.io_diffCommits_info_196_ldest = RTL_PATH.io_diffCommits_info_196_ldest; \
        force U_IF_NAME.io_diffCommits_info_196_pdest = RTL_PATH.io_diffCommits_info_196_pdest; \
        force U_IF_NAME.io_diffCommits_info_196_rfWen = RTL_PATH.io_diffCommits_info_196_rfWen; \
        force U_IF_NAME.io_diffCommits_info_196_fpWen = RTL_PATH.io_diffCommits_info_196_fpWen; \
        force U_IF_NAME.io_diffCommits_info_196_vecWen = RTL_PATH.io_diffCommits_info_196_vecWen; \
        force U_IF_NAME.io_diffCommits_info_196_v0Wen = RTL_PATH.io_diffCommits_info_196_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_196_vlWen = RTL_PATH.io_diffCommits_info_196_vlWen; \
        force U_IF_NAME.io_diffCommits_info_197_ldest = RTL_PATH.io_diffCommits_info_197_ldest; \
        force U_IF_NAME.io_diffCommits_info_197_pdest = RTL_PATH.io_diffCommits_info_197_pdest; \
        force U_IF_NAME.io_diffCommits_info_197_rfWen = RTL_PATH.io_diffCommits_info_197_rfWen; \
        force U_IF_NAME.io_diffCommits_info_197_fpWen = RTL_PATH.io_diffCommits_info_197_fpWen; \
        force U_IF_NAME.io_diffCommits_info_197_vecWen = RTL_PATH.io_diffCommits_info_197_vecWen; \
        force U_IF_NAME.io_diffCommits_info_197_v0Wen = RTL_PATH.io_diffCommits_info_197_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_197_vlWen = RTL_PATH.io_diffCommits_info_197_vlWen; \
        force U_IF_NAME.io_diffCommits_info_198_ldest = RTL_PATH.io_diffCommits_info_198_ldest; \
        force U_IF_NAME.io_diffCommits_info_198_pdest = RTL_PATH.io_diffCommits_info_198_pdest; \
        force U_IF_NAME.io_diffCommits_info_198_rfWen = RTL_PATH.io_diffCommits_info_198_rfWen; \
        force U_IF_NAME.io_diffCommits_info_198_fpWen = RTL_PATH.io_diffCommits_info_198_fpWen; \
        force U_IF_NAME.io_diffCommits_info_198_vecWen = RTL_PATH.io_diffCommits_info_198_vecWen; \
        force U_IF_NAME.io_diffCommits_info_198_v0Wen = RTL_PATH.io_diffCommits_info_198_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_198_vlWen = RTL_PATH.io_diffCommits_info_198_vlWen; \
        force U_IF_NAME.io_diffCommits_info_199_ldest = RTL_PATH.io_diffCommits_info_199_ldest; \
        force U_IF_NAME.io_diffCommits_info_199_pdest = RTL_PATH.io_diffCommits_info_199_pdest; \
        force U_IF_NAME.io_diffCommits_info_199_rfWen = RTL_PATH.io_diffCommits_info_199_rfWen; \
        force U_IF_NAME.io_diffCommits_info_199_fpWen = RTL_PATH.io_diffCommits_info_199_fpWen; \
        force U_IF_NAME.io_diffCommits_info_199_vecWen = RTL_PATH.io_diffCommits_info_199_vecWen; \
        force U_IF_NAME.io_diffCommits_info_199_v0Wen = RTL_PATH.io_diffCommits_info_199_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_199_vlWen = RTL_PATH.io_diffCommits_info_199_vlWen; \
        force U_IF_NAME.io_diffCommits_info_200_ldest = RTL_PATH.io_diffCommits_info_200_ldest; \
        force U_IF_NAME.io_diffCommits_info_200_pdest = RTL_PATH.io_diffCommits_info_200_pdest; \
        force U_IF_NAME.io_diffCommits_info_200_rfWen = RTL_PATH.io_diffCommits_info_200_rfWen; \
        force U_IF_NAME.io_diffCommits_info_200_fpWen = RTL_PATH.io_diffCommits_info_200_fpWen; \
        force U_IF_NAME.io_diffCommits_info_200_vecWen = RTL_PATH.io_diffCommits_info_200_vecWen; \
        force U_IF_NAME.io_diffCommits_info_200_v0Wen = RTL_PATH.io_diffCommits_info_200_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_200_vlWen = RTL_PATH.io_diffCommits_info_200_vlWen; \
        force U_IF_NAME.io_diffCommits_info_201_ldest = RTL_PATH.io_diffCommits_info_201_ldest; \
        force U_IF_NAME.io_diffCommits_info_201_pdest = RTL_PATH.io_diffCommits_info_201_pdest; \
        force U_IF_NAME.io_diffCommits_info_201_rfWen = RTL_PATH.io_diffCommits_info_201_rfWen; \
        force U_IF_NAME.io_diffCommits_info_201_fpWen = RTL_PATH.io_diffCommits_info_201_fpWen; \
        force U_IF_NAME.io_diffCommits_info_201_vecWen = RTL_PATH.io_diffCommits_info_201_vecWen; \
        force U_IF_NAME.io_diffCommits_info_201_v0Wen = RTL_PATH.io_diffCommits_info_201_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_201_vlWen = RTL_PATH.io_diffCommits_info_201_vlWen; \
        force U_IF_NAME.io_diffCommits_info_202_ldest = RTL_PATH.io_diffCommits_info_202_ldest; \
        force U_IF_NAME.io_diffCommits_info_202_pdest = RTL_PATH.io_diffCommits_info_202_pdest; \
        force U_IF_NAME.io_diffCommits_info_202_rfWen = RTL_PATH.io_diffCommits_info_202_rfWen; \
        force U_IF_NAME.io_diffCommits_info_202_fpWen = RTL_PATH.io_diffCommits_info_202_fpWen; \
        force U_IF_NAME.io_diffCommits_info_202_vecWen = RTL_PATH.io_diffCommits_info_202_vecWen; \
        force U_IF_NAME.io_diffCommits_info_202_v0Wen = RTL_PATH.io_diffCommits_info_202_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_202_vlWen = RTL_PATH.io_diffCommits_info_202_vlWen; \
        force U_IF_NAME.io_diffCommits_info_203_ldest = RTL_PATH.io_diffCommits_info_203_ldest; \
        force U_IF_NAME.io_diffCommits_info_203_pdest = RTL_PATH.io_diffCommits_info_203_pdest; \
        force U_IF_NAME.io_diffCommits_info_203_rfWen = RTL_PATH.io_diffCommits_info_203_rfWen; \
        force U_IF_NAME.io_diffCommits_info_203_fpWen = RTL_PATH.io_diffCommits_info_203_fpWen; \
        force U_IF_NAME.io_diffCommits_info_203_vecWen = RTL_PATH.io_diffCommits_info_203_vecWen; \
        force U_IF_NAME.io_diffCommits_info_203_v0Wen = RTL_PATH.io_diffCommits_info_203_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_203_vlWen = RTL_PATH.io_diffCommits_info_203_vlWen; \
        force U_IF_NAME.io_diffCommits_info_204_ldest = RTL_PATH.io_diffCommits_info_204_ldest; \
        force U_IF_NAME.io_diffCommits_info_204_pdest = RTL_PATH.io_diffCommits_info_204_pdest; \
        force U_IF_NAME.io_diffCommits_info_204_rfWen = RTL_PATH.io_diffCommits_info_204_rfWen; \
        force U_IF_NAME.io_diffCommits_info_204_fpWen = RTL_PATH.io_diffCommits_info_204_fpWen; \
        force U_IF_NAME.io_diffCommits_info_204_vecWen = RTL_PATH.io_diffCommits_info_204_vecWen; \
        force U_IF_NAME.io_diffCommits_info_204_v0Wen = RTL_PATH.io_diffCommits_info_204_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_204_vlWen = RTL_PATH.io_diffCommits_info_204_vlWen; \
        force U_IF_NAME.io_diffCommits_info_205_ldest = RTL_PATH.io_diffCommits_info_205_ldest; \
        force U_IF_NAME.io_diffCommits_info_205_pdest = RTL_PATH.io_diffCommits_info_205_pdest; \
        force U_IF_NAME.io_diffCommits_info_205_rfWen = RTL_PATH.io_diffCommits_info_205_rfWen; \
        force U_IF_NAME.io_diffCommits_info_205_fpWen = RTL_PATH.io_diffCommits_info_205_fpWen; \
        force U_IF_NAME.io_diffCommits_info_205_vecWen = RTL_PATH.io_diffCommits_info_205_vecWen; \
        force U_IF_NAME.io_diffCommits_info_205_v0Wen = RTL_PATH.io_diffCommits_info_205_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_205_vlWen = RTL_PATH.io_diffCommits_info_205_vlWen; \
        force U_IF_NAME.io_diffCommits_info_206_ldest = RTL_PATH.io_diffCommits_info_206_ldest; \
        force U_IF_NAME.io_diffCommits_info_206_pdest = RTL_PATH.io_diffCommits_info_206_pdest; \
        force U_IF_NAME.io_diffCommits_info_206_rfWen = RTL_PATH.io_diffCommits_info_206_rfWen; \
        force U_IF_NAME.io_diffCommits_info_206_fpWen = RTL_PATH.io_diffCommits_info_206_fpWen; \
        force U_IF_NAME.io_diffCommits_info_206_vecWen = RTL_PATH.io_diffCommits_info_206_vecWen; \
        force U_IF_NAME.io_diffCommits_info_206_v0Wen = RTL_PATH.io_diffCommits_info_206_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_206_vlWen = RTL_PATH.io_diffCommits_info_206_vlWen; \
        force U_IF_NAME.io_diffCommits_info_207_ldest = RTL_PATH.io_diffCommits_info_207_ldest; \
        force U_IF_NAME.io_diffCommits_info_207_pdest = RTL_PATH.io_diffCommits_info_207_pdest; \
        force U_IF_NAME.io_diffCommits_info_207_rfWen = RTL_PATH.io_diffCommits_info_207_rfWen; \
        force U_IF_NAME.io_diffCommits_info_207_fpWen = RTL_PATH.io_diffCommits_info_207_fpWen; \
        force U_IF_NAME.io_diffCommits_info_207_vecWen = RTL_PATH.io_diffCommits_info_207_vecWen; \
        force U_IF_NAME.io_diffCommits_info_207_v0Wen = RTL_PATH.io_diffCommits_info_207_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_207_vlWen = RTL_PATH.io_diffCommits_info_207_vlWen; \
        force U_IF_NAME.io_diffCommits_info_208_ldest = RTL_PATH.io_diffCommits_info_208_ldest; \
        force U_IF_NAME.io_diffCommits_info_208_pdest = RTL_PATH.io_diffCommits_info_208_pdest; \
        force U_IF_NAME.io_diffCommits_info_208_rfWen = RTL_PATH.io_diffCommits_info_208_rfWen; \
        force U_IF_NAME.io_diffCommits_info_208_fpWen = RTL_PATH.io_diffCommits_info_208_fpWen; \
        force U_IF_NAME.io_diffCommits_info_208_vecWen = RTL_PATH.io_diffCommits_info_208_vecWen; \
        force U_IF_NAME.io_diffCommits_info_208_v0Wen = RTL_PATH.io_diffCommits_info_208_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_208_vlWen = RTL_PATH.io_diffCommits_info_208_vlWen; \
        force U_IF_NAME.io_diffCommits_info_209_ldest = RTL_PATH.io_diffCommits_info_209_ldest; \
        force U_IF_NAME.io_diffCommits_info_209_pdest = RTL_PATH.io_diffCommits_info_209_pdest; \
        force U_IF_NAME.io_diffCommits_info_209_rfWen = RTL_PATH.io_diffCommits_info_209_rfWen; \
        force U_IF_NAME.io_diffCommits_info_209_fpWen = RTL_PATH.io_diffCommits_info_209_fpWen; \
        force U_IF_NAME.io_diffCommits_info_209_vecWen = RTL_PATH.io_diffCommits_info_209_vecWen; \
        force U_IF_NAME.io_diffCommits_info_209_v0Wen = RTL_PATH.io_diffCommits_info_209_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_209_vlWen = RTL_PATH.io_diffCommits_info_209_vlWen; \
        force U_IF_NAME.io_diffCommits_info_210_ldest = RTL_PATH.io_diffCommits_info_210_ldest; \
        force U_IF_NAME.io_diffCommits_info_210_pdest = RTL_PATH.io_diffCommits_info_210_pdest; \
        force U_IF_NAME.io_diffCommits_info_210_rfWen = RTL_PATH.io_diffCommits_info_210_rfWen; \
        force U_IF_NAME.io_diffCommits_info_210_fpWen = RTL_PATH.io_diffCommits_info_210_fpWen; \
        force U_IF_NAME.io_diffCommits_info_210_vecWen = RTL_PATH.io_diffCommits_info_210_vecWen; \
        force U_IF_NAME.io_diffCommits_info_210_v0Wen = RTL_PATH.io_diffCommits_info_210_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_210_vlWen = RTL_PATH.io_diffCommits_info_210_vlWen; \
        force U_IF_NAME.io_diffCommits_info_211_ldest = RTL_PATH.io_diffCommits_info_211_ldest; \
        force U_IF_NAME.io_diffCommits_info_211_pdest = RTL_PATH.io_diffCommits_info_211_pdest; \
        force U_IF_NAME.io_diffCommits_info_211_rfWen = RTL_PATH.io_diffCommits_info_211_rfWen; \
        force U_IF_NAME.io_diffCommits_info_211_fpWen = RTL_PATH.io_diffCommits_info_211_fpWen; \
        force U_IF_NAME.io_diffCommits_info_211_vecWen = RTL_PATH.io_diffCommits_info_211_vecWen; \
        force U_IF_NAME.io_diffCommits_info_211_v0Wen = RTL_PATH.io_diffCommits_info_211_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_211_vlWen = RTL_PATH.io_diffCommits_info_211_vlWen; \
        force U_IF_NAME.io_diffCommits_info_212_ldest = RTL_PATH.io_diffCommits_info_212_ldest; \
        force U_IF_NAME.io_diffCommits_info_212_pdest = RTL_PATH.io_diffCommits_info_212_pdest; \
        force U_IF_NAME.io_diffCommits_info_212_rfWen = RTL_PATH.io_diffCommits_info_212_rfWen; \
        force U_IF_NAME.io_diffCommits_info_212_fpWen = RTL_PATH.io_diffCommits_info_212_fpWen; \
        force U_IF_NAME.io_diffCommits_info_212_vecWen = RTL_PATH.io_diffCommits_info_212_vecWen; \
        force U_IF_NAME.io_diffCommits_info_212_v0Wen = RTL_PATH.io_diffCommits_info_212_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_212_vlWen = RTL_PATH.io_diffCommits_info_212_vlWen; \
        force U_IF_NAME.io_diffCommits_info_213_ldest = RTL_PATH.io_diffCommits_info_213_ldest; \
        force U_IF_NAME.io_diffCommits_info_213_pdest = RTL_PATH.io_diffCommits_info_213_pdest; \
        force U_IF_NAME.io_diffCommits_info_213_rfWen = RTL_PATH.io_diffCommits_info_213_rfWen; \
        force U_IF_NAME.io_diffCommits_info_213_fpWen = RTL_PATH.io_diffCommits_info_213_fpWen; \
        force U_IF_NAME.io_diffCommits_info_213_vecWen = RTL_PATH.io_diffCommits_info_213_vecWen; \
        force U_IF_NAME.io_diffCommits_info_213_v0Wen = RTL_PATH.io_diffCommits_info_213_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_213_vlWen = RTL_PATH.io_diffCommits_info_213_vlWen; \
        force U_IF_NAME.io_diffCommits_info_214_ldest = RTL_PATH.io_diffCommits_info_214_ldest; \
        force U_IF_NAME.io_diffCommits_info_214_pdest = RTL_PATH.io_diffCommits_info_214_pdest; \
        force U_IF_NAME.io_diffCommits_info_214_rfWen = RTL_PATH.io_diffCommits_info_214_rfWen; \
        force U_IF_NAME.io_diffCommits_info_214_fpWen = RTL_PATH.io_diffCommits_info_214_fpWen; \
        force U_IF_NAME.io_diffCommits_info_214_vecWen = RTL_PATH.io_diffCommits_info_214_vecWen; \
        force U_IF_NAME.io_diffCommits_info_214_v0Wen = RTL_PATH.io_diffCommits_info_214_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_214_vlWen = RTL_PATH.io_diffCommits_info_214_vlWen; \
        force U_IF_NAME.io_diffCommits_info_215_ldest = RTL_PATH.io_diffCommits_info_215_ldest; \
        force U_IF_NAME.io_diffCommits_info_215_pdest = RTL_PATH.io_diffCommits_info_215_pdest; \
        force U_IF_NAME.io_diffCommits_info_215_rfWen = RTL_PATH.io_diffCommits_info_215_rfWen; \
        force U_IF_NAME.io_diffCommits_info_215_fpWen = RTL_PATH.io_diffCommits_info_215_fpWen; \
        force U_IF_NAME.io_diffCommits_info_215_vecWen = RTL_PATH.io_diffCommits_info_215_vecWen; \
        force U_IF_NAME.io_diffCommits_info_215_v0Wen = RTL_PATH.io_diffCommits_info_215_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_215_vlWen = RTL_PATH.io_diffCommits_info_215_vlWen; \
        force U_IF_NAME.io_diffCommits_info_216_ldest = RTL_PATH.io_diffCommits_info_216_ldest; \
        force U_IF_NAME.io_diffCommits_info_216_pdest = RTL_PATH.io_diffCommits_info_216_pdest; \
        force U_IF_NAME.io_diffCommits_info_216_rfWen = RTL_PATH.io_diffCommits_info_216_rfWen; \
        force U_IF_NAME.io_diffCommits_info_216_fpWen = RTL_PATH.io_diffCommits_info_216_fpWen; \
        force U_IF_NAME.io_diffCommits_info_216_vecWen = RTL_PATH.io_diffCommits_info_216_vecWen; \
        force U_IF_NAME.io_diffCommits_info_216_v0Wen = RTL_PATH.io_diffCommits_info_216_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_216_vlWen = RTL_PATH.io_diffCommits_info_216_vlWen; \
        force U_IF_NAME.io_diffCommits_info_217_ldest = RTL_PATH.io_diffCommits_info_217_ldest; \
        force U_IF_NAME.io_diffCommits_info_217_pdest = RTL_PATH.io_diffCommits_info_217_pdest; \
        force U_IF_NAME.io_diffCommits_info_217_rfWen = RTL_PATH.io_diffCommits_info_217_rfWen; \
        force U_IF_NAME.io_diffCommits_info_217_fpWen = RTL_PATH.io_diffCommits_info_217_fpWen; \
        force U_IF_NAME.io_diffCommits_info_217_vecWen = RTL_PATH.io_diffCommits_info_217_vecWen; \
        force U_IF_NAME.io_diffCommits_info_217_v0Wen = RTL_PATH.io_diffCommits_info_217_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_217_vlWen = RTL_PATH.io_diffCommits_info_217_vlWen; \
        force U_IF_NAME.io_diffCommits_info_218_ldest = RTL_PATH.io_diffCommits_info_218_ldest; \
        force U_IF_NAME.io_diffCommits_info_218_pdest = RTL_PATH.io_diffCommits_info_218_pdest; \
        force U_IF_NAME.io_diffCommits_info_218_rfWen = RTL_PATH.io_diffCommits_info_218_rfWen; \
        force U_IF_NAME.io_diffCommits_info_218_fpWen = RTL_PATH.io_diffCommits_info_218_fpWen; \
        force U_IF_NAME.io_diffCommits_info_218_vecWen = RTL_PATH.io_diffCommits_info_218_vecWen; \
        force U_IF_NAME.io_diffCommits_info_218_v0Wen = RTL_PATH.io_diffCommits_info_218_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_218_vlWen = RTL_PATH.io_diffCommits_info_218_vlWen; \
        force U_IF_NAME.io_diffCommits_info_219_ldest = RTL_PATH.io_diffCommits_info_219_ldest; \
        force U_IF_NAME.io_diffCommits_info_219_pdest = RTL_PATH.io_diffCommits_info_219_pdest; \
        force U_IF_NAME.io_diffCommits_info_219_rfWen = RTL_PATH.io_diffCommits_info_219_rfWen; \
        force U_IF_NAME.io_diffCommits_info_219_fpWen = RTL_PATH.io_diffCommits_info_219_fpWen; \
        force U_IF_NAME.io_diffCommits_info_219_vecWen = RTL_PATH.io_diffCommits_info_219_vecWen; \
        force U_IF_NAME.io_diffCommits_info_219_v0Wen = RTL_PATH.io_diffCommits_info_219_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_219_vlWen = RTL_PATH.io_diffCommits_info_219_vlWen; \
        force U_IF_NAME.io_diffCommits_info_220_ldest = RTL_PATH.io_diffCommits_info_220_ldest; \
        force U_IF_NAME.io_diffCommits_info_220_pdest = RTL_PATH.io_diffCommits_info_220_pdest; \
        force U_IF_NAME.io_diffCommits_info_220_rfWen = RTL_PATH.io_diffCommits_info_220_rfWen; \
        force U_IF_NAME.io_diffCommits_info_220_fpWen = RTL_PATH.io_diffCommits_info_220_fpWen; \
        force U_IF_NAME.io_diffCommits_info_220_vecWen = RTL_PATH.io_diffCommits_info_220_vecWen; \
        force U_IF_NAME.io_diffCommits_info_220_v0Wen = RTL_PATH.io_diffCommits_info_220_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_220_vlWen = RTL_PATH.io_diffCommits_info_220_vlWen; \
        force U_IF_NAME.io_diffCommits_info_221_ldest = RTL_PATH.io_diffCommits_info_221_ldest; \
        force U_IF_NAME.io_diffCommits_info_221_pdest = RTL_PATH.io_diffCommits_info_221_pdest; \
        force U_IF_NAME.io_diffCommits_info_221_rfWen = RTL_PATH.io_diffCommits_info_221_rfWen; \
        force U_IF_NAME.io_diffCommits_info_221_fpWen = RTL_PATH.io_diffCommits_info_221_fpWen; \
        force U_IF_NAME.io_diffCommits_info_221_vecWen = RTL_PATH.io_diffCommits_info_221_vecWen; \
        force U_IF_NAME.io_diffCommits_info_221_v0Wen = RTL_PATH.io_diffCommits_info_221_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_221_vlWen = RTL_PATH.io_diffCommits_info_221_vlWen; \
        force U_IF_NAME.io_diffCommits_info_222_ldest = RTL_PATH.io_diffCommits_info_222_ldest; \
        force U_IF_NAME.io_diffCommits_info_222_pdest = RTL_PATH.io_diffCommits_info_222_pdest; \
        force U_IF_NAME.io_diffCommits_info_222_rfWen = RTL_PATH.io_diffCommits_info_222_rfWen; \
        force U_IF_NAME.io_diffCommits_info_222_fpWen = RTL_PATH.io_diffCommits_info_222_fpWen; \
        force U_IF_NAME.io_diffCommits_info_222_vecWen = RTL_PATH.io_diffCommits_info_222_vecWen; \
        force U_IF_NAME.io_diffCommits_info_222_v0Wen = RTL_PATH.io_diffCommits_info_222_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_222_vlWen = RTL_PATH.io_diffCommits_info_222_vlWen; \
        force U_IF_NAME.io_diffCommits_info_223_ldest = RTL_PATH.io_diffCommits_info_223_ldest; \
        force U_IF_NAME.io_diffCommits_info_223_pdest = RTL_PATH.io_diffCommits_info_223_pdest; \
        force U_IF_NAME.io_diffCommits_info_223_rfWen = RTL_PATH.io_diffCommits_info_223_rfWen; \
        force U_IF_NAME.io_diffCommits_info_223_fpWen = RTL_PATH.io_diffCommits_info_223_fpWen; \
        force U_IF_NAME.io_diffCommits_info_223_vecWen = RTL_PATH.io_diffCommits_info_223_vecWen; \
        force U_IF_NAME.io_diffCommits_info_223_v0Wen = RTL_PATH.io_diffCommits_info_223_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_223_vlWen = RTL_PATH.io_diffCommits_info_223_vlWen; \
        force U_IF_NAME.io_diffCommits_info_224_ldest = RTL_PATH.io_diffCommits_info_224_ldest; \
        force U_IF_NAME.io_diffCommits_info_224_pdest = RTL_PATH.io_diffCommits_info_224_pdest; \
        force U_IF_NAME.io_diffCommits_info_224_rfWen = RTL_PATH.io_diffCommits_info_224_rfWen; \
        force U_IF_NAME.io_diffCommits_info_224_fpWen = RTL_PATH.io_diffCommits_info_224_fpWen; \
        force U_IF_NAME.io_diffCommits_info_224_vecWen = RTL_PATH.io_diffCommits_info_224_vecWen; \
        force U_IF_NAME.io_diffCommits_info_224_v0Wen = RTL_PATH.io_diffCommits_info_224_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_224_vlWen = RTL_PATH.io_diffCommits_info_224_vlWen; \
        force U_IF_NAME.io_diffCommits_info_225_ldest = RTL_PATH.io_diffCommits_info_225_ldest; \
        force U_IF_NAME.io_diffCommits_info_225_pdest = RTL_PATH.io_diffCommits_info_225_pdest; \
        force U_IF_NAME.io_diffCommits_info_225_rfWen = RTL_PATH.io_diffCommits_info_225_rfWen; \
        force U_IF_NAME.io_diffCommits_info_225_fpWen = RTL_PATH.io_diffCommits_info_225_fpWen; \
        force U_IF_NAME.io_diffCommits_info_225_vecWen = RTL_PATH.io_diffCommits_info_225_vecWen; \
        force U_IF_NAME.io_diffCommits_info_225_v0Wen = RTL_PATH.io_diffCommits_info_225_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_225_vlWen = RTL_PATH.io_diffCommits_info_225_vlWen; \
        force U_IF_NAME.io_diffCommits_info_226_ldest = RTL_PATH.io_diffCommits_info_226_ldest; \
        force U_IF_NAME.io_diffCommits_info_226_pdest = RTL_PATH.io_diffCommits_info_226_pdest; \
        force U_IF_NAME.io_diffCommits_info_226_rfWen = RTL_PATH.io_diffCommits_info_226_rfWen; \
        force U_IF_NAME.io_diffCommits_info_226_fpWen = RTL_PATH.io_diffCommits_info_226_fpWen; \
        force U_IF_NAME.io_diffCommits_info_226_vecWen = RTL_PATH.io_diffCommits_info_226_vecWen; \
        force U_IF_NAME.io_diffCommits_info_226_v0Wen = RTL_PATH.io_diffCommits_info_226_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_226_vlWen = RTL_PATH.io_diffCommits_info_226_vlWen; \
        force U_IF_NAME.io_diffCommits_info_227_ldest = RTL_PATH.io_diffCommits_info_227_ldest; \
        force U_IF_NAME.io_diffCommits_info_227_pdest = RTL_PATH.io_diffCommits_info_227_pdest; \
        force U_IF_NAME.io_diffCommits_info_227_rfWen = RTL_PATH.io_diffCommits_info_227_rfWen; \
        force U_IF_NAME.io_diffCommits_info_227_fpWen = RTL_PATH.io_diffCommits_info_227_fpWen; \
        force U_IF_NAME.io_diffCommits_info_227_vecWen = RTL_PATH.io_diffCommits_info_227_vecWen; \
        force U_IF_NAME.io_diffCommits_info_227_v0Wen = RTL_PATH.io_diffCommits_info_227_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_227_vlWen = RTL_PATH.io_diffCommits_info_227_vlWen; \
        force U_IF_NAME.io_diffCommits_info_228_ldest = RTL_PATH.io_diffCommits_info_228_ldest; \
        force U_IF_NAME.io_diffCommits_info_228_pdest = RTL_PATH.io_diffCommits_info_228_pdest; \
        force U_IF_NAME.io_diffCommits_info_228_rfWen = RTL_PATH.io_diffCommits_info_228_rfWen; \
        force U_IF_NAME.io_diffCommits_info_228_fpWen = RTL_PATH.io_diffCommits_info_228_fpWen; \
        force U_IF_NAME.io_diffCommits_info_228_vecWen = RTL_PATH.io_diffCommits_info_228_vecWen; \
        force U_IF_NAME.io_diffCommits_info_228_v0Wen = RTL_PATH.io_diffCommits_info_228_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_228_vlWen = RTL_PATH.io_diffCommits_info_228_vlWen; \
        force U_IF_NAME.io_diffCommits_info_229_ldest = RTL_PATH.io_diffCommits_info_229_ldest; \
        force U_IF_NAME.io_diffCommits_info_229_pdest = RTL_PATH.io_diffCommits_info_229_pdest; \
        force U_IF_NAME.io_diffCommits_info_229_rfWen = RTL_PATH.io_diffCommits_info_229_rfWen; \
        force U_IF_NAME.io_diffCommits_info_229_fpWen = RTL_PATH.io_diffCommits_info_229_fpWen; \
        force U_IF_NAME.io_diffCommits_info_229_vecWen = RTL_PATH.io_diffCommits_info_229_vecWen; \
        force U_IF_NAME.io_diffCommits_info_229_v0Wen = RTL_PATH.io_diffCommits_info_229_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_229_vlWen = RTL_PATH.io_diffCommits_info_229_vlWen; \
        force U_IF_NAME.io_diffCommits_info_230_ldest = RTL_PATH.io_diffCommits_info_230_ldest; \
        force U_IF_NAME.io_diffCommits_info_230_pdest = RTL_PATH.io_diffCommits_info_230_pdest; \
        force U_IF_NAME.io_diffCommits_info_230_rfWen = RTL_PATH.io_diffCommits_info_230_rfWen; \
        force U_IF_NAME.io_diffCommits_info_230_fpWen = RTL_PATH.io_diffCommits_info_230_fpWen; \
        force U_IF_NAME.io_diffCommits_info_230_vecWen = RTL_PATH.io_diffCommits_info_230_vecWen; \
        force U_IF_NAME.io_diffCommits_info_230_v0Wen = RTL_PATH.io_diffCommits_info_230_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_230_vlWen = RTL_PATH.io_diffCommits_info_230_vlWen; \
        force U_IF_NAME.io_diffCommits_info_231_ldest = RTL_PATH.io_diffCommits_info_231_ldest; \
        force U_IF_NAME.io_diffCommits_info_231_pdest = RTL_PATH.io_diffCommits_info_231_pdest; \
        force U_IF_NAME.io_diffCommits_info_231_rfWen = RTL_PATH.io_diffCommits_info_231_rfWen; \
        force U_IF_NAME.io_diffCommits_info_231_fpWen = RTL_PATH.io_diffCommits_info_231_fpWen; \
        force U_IF_NAME.io_diffCommits_info_231_vecWen = RTL_PATH.io_diffCommits_info_231_vecWen; \
        force U_IF_NAME.io_diffCommits_info_231_v0Wen = RTL_PATH.io_diffCommits_info_231_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_231_vlWen = RTL_PATH.io_diffCommits_info_231_vlWen; \
        force U_IF_NAME.io_diffCommits_info_232_ldest = RTL_PATH.io_diffCommits_info_232_ldest; \
        force U_IF_NAME.io_diffCommits_info_232_pdest = RTL_PATH.io_diffCommits_info_232_pdest; \
        force U_IF_NAME.io_diffCommits_info_232_rfWen = RTL_PATH.io_diffCommits_info_232_rfWen; \
        force U_IF_NAME.io_diffCommits_info_232_fpWen = RTL_PATH.io_diffCommits_info_232_fpWen; \
        force U_IF_NAME.io_diffCommits_info_232_vecWen = RTL_PATH.io_diffCommits_info_232_vecWen; \
        force U_IF_NAME.io_diffCommits_info_232_v0Wen = RTL_PATH.io_diffCommits_info_232_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_232_vlWen = RTL_PATH.io_diffCommits_info_232_vlWen; \
        force U_IF_NAME.io_diffCommits_info_233_ldest = RTL_PATH.io_diffCommits_info_233_ldest; \
        force U_IF_NAME.io_diffCommits_info_233_pdest = RTL_PATH.io_diffCommits_info_233_pdest; \
        force U_IF_NAME.io_diffCommits_info_233_rfWen = RTL_PATH.io_diffCommits_info_233_rfWen; \
        force U_IF_NAME.io_diffCommits_info_233_fpWen = RTL_PATH.io_diffCommits_info_233_fpWen; \
        force U_IF_NAME.io_diffCommits_info_233_vecWen = RTL_PATH.io_diffCommits_info_233_vecWen; \
        force U_IF_NAME.io_diffCommits_info_233_v0Wen = RTL_PATH.io_diffCommits_info_233_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_233_vlWen = RTL_PATH.io_diffCommits_info_233_vlWen; \
        force U_IF_NAME.io_diffCommits_info_234_ldest = RTL_PATH.io_diffCommits_info_234_ldest; \
        force U_IF_NAME.io_diffCommits_info_234_pdest = RTL_PATH.io_diffCommits_info_234_pdest; \
        force U_IF_NAME.io_diffCommits_info_234_rfWen = RTL_PATH.io_diffCommits_info_234_rfWen; \
        force U_IF_NAME.io_diffCommits_info_234_fpWen = RTL_PATH.io_diffCommits_info_234_fpWen; \
        force U_IF_NAME.io_diffCommits_info_234_vecWen = RTL_PATH.io_diffCommits_info_234_vecWen; \
        force U_IF_NAME.io_diffCommits_info_234_v0Wen = RTL_PATH.io_diffCommits_info_234_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_234_vlWen = RTL_PATH.io_diffCommits_info_234_vlWen; \
        force U_IF_NAME.io_diffCommits_info_235_ldest = RTL_PATH.io_diffCommits_info_235_ldest; \
        force U_IF_NAME.io_diffCommits_info_235_pdest = RTL_PATH.io_diffCommits_info_235_pdest; \
        force U_IF_NAME.io_diffCommits_info_235_rfWen = RTL_PATH.io_diffCommits_info_235_rfWen; \
        force U_IF_NAME.io_diffCommits_info_235_fpWen = RTL_PATH.io_diffCommits_info_235_fpWen; \
        force U_IF_NAME.io_diffCommits_info_235_vecWen = RTL_PATH.io_diffCommits_info_235_vecWen; \
        force U_IF_NAME.io_diffCommits_info_235_v0Wen = RTL_PATH.io_diffCommits_info_235_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_235_vlWen = RTL_PATH.io_diffCommits_info_235_vlWen; \
        force U_IF_NAME.io_diffCommits_info_236_ldest = RTL_PATH.io_diffCommits_info_236_ldest; \
        force U_IF_NAME.io_diffCommits_info_236_pdest = RTL_PATH.io_diffCommits_info_236_pdest; \
        force U_IF_NAME.io_diffCommits_info_236_rfWen = RTL_PATH.io_diffCommits_info_236_rfWen; \
        force U_IF_NAME.io_diffCommits_info_236_fpWen = RTL_PATH.io_diffCommits_info_236_fpWen; \
        force U_IF_NAME.io_diffCommits_info_236_vecWen = RTL_PATH.io_diffCommits_info_236_vecWen; \
        force U_IF_NAME.io_diffCommits_info_236_v0Wen = RTL_PATH.io_diffCommits_info_236_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_236_vlWen = RTL_PATH.io_diffCommits_info_236_vlWen; \
        force U_IF_NAME.io_diffCommits_info_237_ldest = RTL_PATH.io_diffCommits_info_237_ldest; \
        force U_IF_NAME.io_diffCommits_info_237_pdest = RTL_PATH.io_diffCommits_info_237_pdest; \
        force U_IF_NAME.io_diffCommits_info_237_rfWen = RTL_PATH.io_diffCommits_info_237_rfWen; \
        force U_IF_NAME.io_diffCommits_info_237_fpWen = RTL_PATH.io_diffCommits_info_237_fpWen; \
        force U_IF_NAME.io_diffCommits_info_237_vecWen = RTL_PATH.io_diffCommits_info_237_vecWen; \
        force U_IF_NAME.io_diffCommits_info_237_v0Wen = RTL_PATH.io_diffCommits_info_237_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_237_vlWen = RTL_PATH.io_diffCommits_info_237_vlWen; \
        force U_IF_NAME.io_diffCommits_info_238_ldest = RTL_PATH.io_diffCommits_info_238_ldest; \
        force U_IF_NAME.io_diffCommits_info_238_pdest = RTL_PATH.io_diffCommits_info_238_pdest; \
        force U_IF_NAME.io_diffCommits_info_238_rfWen = RTL_PATH.io_diffCommits_info_238_rfWen; \
        force U_IF_NAME.io_diffCommits_info_238_fpWen = RTL_PATH.io_diffCommits_info_238_fpWen; \
        force U_IF_NAME.io_diffCommits_info_238_vecWen = RTL_PATH.io_diffCommits_info_238_vecWen; \
        force U_IF_NAME.io_diffCommits_info_238_v0Wen = RTL_PATH.io_diffCommits_info_238_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_238_vlWen = RTL_PATH.io_diffCommits_info_238_vlWen; \
        force U_IF_NAME.io_diffCommits_info_239_ldest = RTL_PATH.io_diffCommits_info_239_ldest; \
        force U_IF_NAME.io_diffCommits_info_239_pdest = RTL_PATH.io_diffCommits_info_239_pdest; \
        force U_IF_NAME.io_diffCommits_info_239_rfWen = RTL_PATH.io_diffCommits_info_239_rfWen; \
        force U_IF_NAME.io_diffCommits_info_239_fpWen = RTL_PATH.io_diffCommits_info_239_fpWen; \
        force U_IF_NAME.io_diffCommits_info_239_vecWen = RTL_PATH.io_diffCommits_info_239_vecWen; \
        force U_IF_NAME.io_diffCommits_info_239_v0Wen = RTL_PATH.io_diffCommits_info_239_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_239_vlWen = RTL_PATH.io_diffCommits_info_239_vlWen; \
        force U_IF_NAME.io_diffCommits_info_240_ldest = RTL_PATH.io_diffCommits_info_240_ldest; \
        force U_IF_NAME.io_diffCommits_info_240_pdest = RTL_PATH.io_diffCommits_info_240_pdest; \
        force U_IF_NAME.io_diffCommits_info_240_rfWen = RTL_PATH.io_diffCommits_info_240_rfWen; \
        force U_IF_NAME.io_diffCommits_info_240_fpWen = RTL_PATH.io_diffCommits_info_240_fpWen; \
        force U_IF_NAME.io_diffCommits_info_240_vecWen = RTL_PATH.io_diffCommits_info_240_vecWen; \
        force U_IF_NAME.io_diffCommits_info_240_v0Wen = RTL_PATH.io_diffCommits_info_240_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_240_vlWen = RTL_PATH.io_diffCommits_info_240_vlWen; \
        force U_IF_NAME.io_diffCommits_info_241_ldest = RTL_PATH.io_diffCommits_info_241_ldest; \
        force U_IF_NAME.io_diffCommits_info_241_pdest = RTL_PATH.io_diffCommits_info_241_pdest; \
        force U_IF_NAME.io_diffCommits_info_241_rfWen = RTL_PATH.io_diffCommits_info_241_rfWen; \
        force U_IF_NAME.io_diffCommits_info_241_fpWen = RTL_PATH.io_diffCommits_info_241_fpWen; \
        force U_IF_NAME.io_diffCommits_info_241_vecWen = RTL_PATH.io_diffCommits_info_241_vecWen; \
        force U_IF_NAME.io_diffCommits_info_241_v0Wen = RTL_PATH.io_diffCommits_info_241_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_241_vlWen = RTL_PATH.io_diffCommits_info_241_vlWen; \
        force U_IF_NAME.io_diffCommits_info_242_ldest = RTL_PATH.io_diffCommits_info_242_ldest; \
        force U_IF_NAME.io_diffCommits_info_242_pdest = RTL_PATH.io_diffCommits_info_242_pdest; \
        force U_IF_NAME.io_diffCommits_info_242_rfWen = RTL_PATH.io_diffCommits_info_242_rfWen; \
        force U_IF_NAME.io_diffCommits_info_242_fpWen = RTL_PATH.io_diffCommits_info_242_fpWen; \
        force U_IF_NAME.io_diffCommits_info_242_vecWen = RTL_PATH.io_diffCommits_info_242_vecWen; \
        force U_IF_NAME.io_diffCommits_info_242_v0Wen = RTL_PATH.io_diffCommits_info_242_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_242_vlWen = RTL_PATH.io_diffCommits_info_242_vlWen; \
        force U_IF_NAME.io_diffCommits_info_243_ldest = RTL_PATH.io_diffCommits_info_243_ldest; \
        force U_IF_NAME.io_diffCommits_info_243_pdest = RTL_PATH.io_diffCommits_info_243_pdest; \
        force U_IF_NAME.io_diffCommits_info_243_rfWen = RTL_PATH.io_diffCommits_info_243_rfWen; \
        force U_IF_NAME.io_diffCommits_info_243_fpWen = RTL_PATH.io_diffCommits_info_243_fpWen; \
        force U_IF_NAME.io_diffCommits_info_243_vecWen = RTL_PATH.io_diffCommits_info_243_vecWen; \
        force U_IF_NAME.io_diffCommits_info_243_v0Wen = RTL_PATH.io_diffCommits_info_243_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_243_vlWen = RTL_PATH.io_diffCommits_info_243_vlWen; \
        force U_IF_NAME.io_diffCommits_info_244_ldest = RTL_PATH.io_diffCommits_info_244_ldest; \
        force U_IF_NAME.io_diffCommits_info_244_pdest = RTL_PATH.io_diffCommits_info_244_pdest; \
        force U_IF_NAME.io_diffCommits_info_244_rfWen = RTL_PATH.io_diffCommits_info_244_rfWen; \
        force U_IF_NAME.io_diffCommits_info_244_fpWen = RTL_PATH.io_diffCommits_info_244_fpWen; \
        force U_IF_NAME.io_diffCommits_info_244_vecWen = RTL_PATH.io_diffCommits_info_244_vecWen; \
        force U_IF_NAME.io_diffCommits_info_244_v0Wen = RTL_PATH.io_diffCommits_info_244_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_244_vlWen = RTL_PATH.io_diffCommits_info_244_vlWen; \
        force U_IF_NAME.io_diffCommits_info_245_ldest = RTL_PATH.io_diffCommits_info_245_ldest; \
        force U_IF_NAME.io_diffCommits_info_245_pdest = RTL_PATH.io_diffCommits_info_245_pdest; \
        force U_IF_NAME.io_diffCommits_info_245_rfWen = RTL_PATH.io_diffCommits_info_245_rfWen; \
        force U_IF_NAME.io_diffCommits_info_245_fpWen = RTL_PATH.io_diffCommits_info_245_fpWen; \
        force U_IF_NAME.io_diffCommits_info_245_vecWen = RTL_PATH.io_diffCommits_info_245_vecWen; \
        force U_IF_NAME.io_diffCommits_info_245_v0Wen = RTL_PATH.io_diffCommits_info_245_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_245_vlWen = RTL_PATH.io_diffCommits_info_245_vlWen; \
        force U_IF_NAME.io_diffCommits_info_246_ldest = RTL_PATH.io_diffCommits_info_246_ldest; \
        force U_IF_NAME.io_diffCommits_info_246_pdest = RTL_PATH.io_diffCommits_info_246_pdest; \
        force U_IF_NAME.io_diffCommits_info_246_rfWen = RTL_PATH.io_diffCommits_info_246_rfWen; \
        force U_IF_NAME.io_diffCommits_info_246_fpWen = RTL_PATH.io_diffCommits_info_246_fpWen; \
        force U_IF_NAME.io_diffCommits_info_246_vecWen = RTL_PATH.io_diffCommits_info_246_vecWen; \
        force U_IF_NAME.io_diffCommits_info_246_v0Wen = RTL_PATH.io_diffCommits_info_246_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_246_vlWen = RTL_PATH.io_diffCommits_info_246_vlWen; \
        force U_IF_NAME.io_diffCommits_info_247_ldest = RTL_PATH.io_diffCommits_info_247_ldest; \
        force U_IF_NAME.io_diffCommits_info_247_pdest = RTL_PATH.io_diffCommits_info_247_pdest; \
        force U_IF_NAME.io_diffCommits_info_247_rfWen = RTL_PATH.io_diffCommits_info_247_rfWen; \
        force U_IF_NAME.io_diffCommits_info_247_fpWen = RTL_PATH.io_diffCommits_info_247_fpWen; \
        force U_IF_NAME.io_diffCommits_info_247_vecWen = RTL_PATH.io_diffCommits_info_247_vecWen; \
        force U_IF_NAME.io_diffCommits_info_247_v0Wen = RTL_PATH.io_diffCommits_info_247_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_247_vlWen = RTL_PATH.io_diffCommits_info_247_vlWen; \
        force U_IF_NAME.io_diffCommits_info_248_ldest = RTL_PATH.io_diffCommits_info_248_ldest; \
        force U_IF_NAME.io_diffCommits_info_248_pdest = RTL_PATH.io_diffCommits_info_248_pdest; \
        force U_IF_NAME.io_diffCommits_info_248_rfWen = RTL_PATH.io_diffCommits_info_248_rfWen; \
        force U_IF_NAME.io_diffCommits_info_248_fpWen = RTL_PATH.io_diffCommits_info_248_fpWen; \
        force U_IF_NAME.io_diffCommits_info_248_vecWen = RTL_PATH.io_diffCommits_info_248_vecWen; \
        force U_IF_NAME.io_diffCommits_info_248_v0Wen = RTL_PATH.io_diffCommits_info_248_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_248_vlWen = RTL_PATH.io_diffCommits_info_248_vlWen; \
        force U_IF_NAME.io_diffCommits_info_249_ldest = RTL_PATH.io_diffCommits_info_249_ldest; \
        force U_IF_NAME.io_diffCommits_info_249_pdest = RTL_PATH.io_diffCommits_info_249_pdest; \
        force U_IF_NAME.io_diffCommits_info_249_rfWen = RTL_PATH.io_diffCommits_info_249_rfWen; \
        force U_IF_NAME.io_diffCommits_info_249_fpWen = RTL_PATH.io_diffCommits_info_249_fpWen; \
        force U_IF_NAME.io_diffCommits_info_249_vecWen = RTL_PATH.io_diffCommits_info_249_vecWen; \
        force U_IF_NAME.io_diffCommits_info_249_v0Wen = RTL_PATH.io_diffCommits_info_249_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_249_vlWen = RTL_PATH.io_diffCommits_info_249_vlWen; \
        force U_IF_NAME.io_diffCommits_info_250_ldest = RTL_PATH.io_diffCommits_info_250_ldest; \
        force U_IF_NAME.io_diffCommits_info_250_pdest = RTL_PATH.io_diffCommits_info_250_pdest; \
        force U_IF_NAME.io_diffCommits_info_250_rfWen = RTL_PATH.io_diffCommits_info_250_rfWen; \
        force U_IF_NAME.io_diffCommits_info_250_fpWen = RTL_PATH.io_diffCommits_info_250_fpWen; \
        force U_IF_NAME.io_diffCommits_info_250_vecWen = RTL_PATH.io_diffCommits_info_250_vecWen; \
        force U_IF_NAME.io_diffCommits_info_250_v0Wen = RTL_PATH.io_diffCommits_info_250_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_250_vlWen = RTL_PATH.io_diffCommits_info_250_vlWen; \
        force U_IF_NAME.io_diffCommits_info_251_ldest = RTL_PATH.io_diffCommits_info_251_ldest; \
        force U_IF_NAME.io_diffCommits_info_251_pdest = RTL_PATH.io_diffCommits_info_251_pdest; \
        force U_IF_NAME.io_diffCommits_info_251_rfWen = RTL_PATH.io_diffCommits_info_251_rfWen; \
        force U_IF_NAME.io_diffCommits_info_251_fpWen = RTL_PATH.io_diffCommits_info_251_fpWen; \
        force U_IF_NAME.io_diffCommits_info_251_vecWen = RTL_PATH.io_diffCommits_info_251_vecWen; \
        force U_IF_NAME.io_diffCommits_info_251_v0Wen = RTL_PATH.io_diffCommits_info_251_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_251_vlWen = RTL_PATH.io_diffCommits_info_251_vlWen; \
        force U_IF_NAME.io_diffCommits_info_252_ldest = RTL_PATH.io_diffCommits_info_252_ldest; \
        force U_IF_NAME.io_diffCommits_info_252_pdest = RTL_PATH.io_diffCommits_info_252_pdest; \
        force U_IF_NAME.io_diffCommits_info_252_rfWen = RTL_PATH.io_diffCommits_info_252_rfWen; \
        force U_IF_NAME.io_diffCommits_info_252_fpWen = RTL_PATH.io_diffCommits_info_252_fpWen; \
        force U_IF_NAME.io_diffCommits_info_252_vecWen = RTL_PATH.io_diffCommits_info_252_vecWen; \
        force U_IF_NAME.io_diffCommits_info_252_v0Wen = RTL_PATH.io_diffCommits_info_252_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_252_vlWen = RTL_PATH.io_diffCommits_info_252_vlWen; \
        force U_IF_NAME.io_diffCommits_info_253_ldest = RTL_PATH.io_diffCommits_info_253_ldest; \
        force U_IF_NAME.io_diffCommits_info_253_pdest = RTL_PATH.io_diffCommits_info_253_pdest; \
        force U_IF_NAME.io_diffCommits_info_253_rfWen = RTL_PATH.io_diffCommits_info_253_rfWen; \
        force U_IF_NAME.io_diffCommits_info_253_fpWen = RTL_PATH.io_diffCommits_info_253_fpWen; \
        force U_IF_NAME.io_diffCommits_info_253_vecWen = RTL_PATH.io_diffCommits_info_253_vecWen; \
        force U_IF_NAME.io_diffCommits_info_253_v0Wen = RTL_PATH.io_diffCommits_info_253_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_253_vlWen = RTL_PATH.io_diffCommits_info_253_vlWen; \
        force U_IF_NAME.io_diffCommits_info_254_ldest = RTL_PATH.io_diffCommits_info_254_ldest; \
        force U_IF_NAME.io_diffCommits_info_254_pdest = RTL_PATH.io_diffCommits_info_254_pdest; \
        force U_IF_NAME.io_diffCommits_info_254_rfWen = RTL_PATH.io_diffCommits_info_254_rfWen; \
        force U_IF_NAME.io_diffCommits_info_254_fpWen = RTL_PATH.io_diffCommits_info_254_fpWen; \
        force U_IF_NAME.io_diffCommits_info_254_vecWen = RTL_PATH.io_diffCommits_info_254_vecWen; \
        force U_IF_NAME.io_diffCommits_info_254_v0Wen = RTL_PATH.io_diffCommits_info_254_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_254_vlWen = RTL_PATH.io_diffCommits_info_254_vlWen; \
        force U_IF_NAME.io_diffCommits_info_255_ldest = RTL_PATH.io_diffCommits_info_255_ldest; \
        force U_IF_NAME.io_diffCommits_info_255_pdest = RTL_PATH.io_diffCommits_info_255_pdest; \
        force U_IF_NAME.io_diffCommits_info_256_ldest = RTL_PATH.io_diffCommits_info_256_ldest; \
        force U_IF_NAME.io_diffCommits_info_256_pdest = RTL_PATH.io_diffCommits_info_256_pdest; \
        force U_IF_NAME.io_diffCommits_info_257_ldest = RTL_PATH.io_diffCommits_info_257_ldest; \
        force U_IF_NAME.io_diffCommits_info_257_pdest = RTL_PATH.io_diffCommits_info_257_pdest; \
        force U_IF_NAME.io_diffCommits_info_258_ldest = RTL_PATH.io_diffCommits_info_258_ldest; \
        force U_IF_NAME.io_diffCommits_info_258_pdest = RTL_PATH.io_diffCommits_info_258_pdest; \
        force U_IF_NAME.io_diffCommits_info_259_ldest = RTL_PATH.io_diffCommits_info_259_ldest; \
        force U_IF_NAME.io_diffCommits_info_259_pdest = RTL_PATH.io_diffCommits_info_259_pdest; \
        force U_IF_NAME.io_diffCommits_info_260_ldest = RTL_PATH.io_diffCommits_info_260_ldest; \
        force U_IF_NAME.io_diffCommits_info_260_pdest = RTL_PATH.io_diffCommits_info_260_pdest; \
        force U_IF_NAME.io_diffCommits_info_261_ldest = RTL_PATH.io_diffCommits_info_261_ldest; \
        force U_IF_NAME.io_diffCommits_info_261_pdest = RTL_PATH.io_diffCommits_info_261_pdest; \
        force U_IF_NAME.io_diffCommits_info_262_ldest = RTL_PATH.io_diffCommits_info_262_ldest; \
        force U_IF_NAME.io_diffCommits_info_262_pdest = RTL_PATH.io_diffCommits_info_262_pdest; \
        force U_IF_NAME.io_diffCommits_info_263_ldest = RTL_PATH.io_diffCommits_info_263_ldest; \
        force U_IF_NAME.io_diffCommits_info_263_pdest = RTL_PATH.io_diffCommits_info_263_pdest; \
        force U_IF_NAME.io_diffCommits_info_264_ldest = RTL_PATH.io_diffCommits_info_264_ldest; \
        force U_IF_NAME.io_diffCommits_info_264_pdest = RTL_PATH.io_diffCommits_info_264_pdest; \
        force U_IF_NAME.io_diffCommits_info_265_ldest = RTL_PATH.io_diffCommits_info_265_ldest; \
        force U_IF_NAME.io_diffCommits_info_265_pdest = RTL_PATH.io_diffCommits_info_265_pdest; \
        force U_IF_NAME.io_diffCommits_info_266_ldest = RTL_PATH.io_diffCommits_info_266_ldest; \
        force U_IF_NAME.io_diffCommits_info_266_pdest = RTL_PATH.io_diffCommits_info_266_pdest; \
        force U_IF_NAME.io_diffCommits_info_267_ldest = RTL_PATH.io_diffCommits_info_267_ldest; \
        force U_IF_NAME.io_diffCommits_info_267_pdest = RTL_PATH.io_diffCommits_info_267_pdest; \
        force U_IF_NAME.io_diffCommits_info_268_ldest = RTL_PATH.io_diffCommits_info_268_ldest; \
        force U_IF_NAME.io_diffCommits_info_268_pdest = RTL_PATH.io_diffCommits_info_268_pdest; \
        force U_IF_NAME.io_diffCommits_info_269_ldest = RTL_PATH.io_diffCommits_info_269_ldest; \
        force U_IF_NAME.io_diffCommits_info_269_pdest = RTL_PATH.io_diffCommits_info_269_pdest; \
        force U_IF_NAME.io_diffCommits_info_270_ldest = RTL_PATH.io_diffCommits_info_270_ldest; \
        force U_IF_NAME.io_diffCommits_info_270_pdest = RTL_PATH.io_diffCommits_info_270_pdest; \
        force U_IF_NAME.io_diffCommits_info_271_ldest = RTL_PATH.io_diffCommits_info_271_ldest; \
        force U_IF_NAME.io_diffCommits_info_271_pdest = RTL_PATH.io_diffCommits_info_271_pdest; \
        force U_IF_NAME.io_diffCommits_info_272_ldest = RTL_PATH.io_diffCommits_info_272_ldest; \
        force U_IF_NAME.io_diffCommits_info_272_pdest = RTL_PATH.io_diffCommits_info_272_pdest; \
        force U_IF_NAME.io_diffCommits_info_273_ldest = RTL_PATH.io_diffCommits_info_273_ldest; \
        force U_IF_NAME.io_diffCommits_info_273_pdest = RTL_PATH.io_diffCommits_info_273_pdest; \
        force U_IF_NAME.io_diffCommits_info_274_ldest = RTL_PATH.io_diffCommits_info_274_ldest; \
        force U_IF_NAME.io_diffCommits_info_274_pdest = RTL_PATH.io_diffCommits_info_274_pdest; \
        force U_IF_NAME.io_diffCommits_info_275_ldest = RTL_PATH.io_diffCommits_info_275_ldest; \
        force U_IF_NAME.io_diffCommits_info_275_pdest = RTL_PATH.io_diffCommits_info_275_pdest; \
        force U_IF_NAME.io_diffCommits_info_276_ldest = RTL_PATH.io_diffCommits_info_276_ldest; \
        force U_IF_NAME.io_diffCommits_info_276_pdest = RTL_PATH.io_diffCommits_info_276_pdest; \
        force U_IF_NAME.io_diffCommits_info_277_ldest = RTL_PATH.io_diffCommits_info_277_ldest; \
        force U_IF_NAME.io_diffCommits_info_277_pdest = RTL_PATH.io_diffCommits_info_277_pdest; \
        force U_IF_NAME.io_diffCommits_info_278_ldest = RTL_PATH.io_diffCommits_info_278_ldest; \
        force U_IF_NAME.io_diffCommits_info_278_pdest = RTL_PATH.io_diffCommits_info_278_pdest; \
        force U_IF_NAME.io_diffCommits_info_279_ldest = RTL_PATH.io_diffCommits_info_279_ldest; \
        force U_IF_NAME.io_diffCommits_info_279_pdest = RTL_PATH.io_diffCommits_info_279_pdest; \
        force U_IF_NAME.io_diffCommits_info_280_ldest = RTL_PATH.io_diffCommits_info_280_ldest; \
        force U_IF_NAME.io_diffCommits_info_280_pdest = RTL_PATH.io_diffCommits_info_280_pdest; \
        force U_IF_NAME.io_diffCommits_info_281_ldest = RTL_PATH.io_diffCommits_info_281_ldest; \
        force U_IF_NAME.io_diffCommits_info_281_pdest = RTL_PATH.io_diffCommits_info_281_pdest; \
        force U_IF_NAME.io_diffCommits_info_282_ldest = RTL_PATH.io_diffCommits_info_282_ldest; \
        force U_IF_NAME.io_diffCommits_info_282_pdest = RTL_PATH.io_diffCommits_info_282_pdest; \
        force U_IF_NAME.io_diffCommits_info_283_ldest = RTL_PATH.io_diffCommits_info_283_ldest; \
        force U_IF_NAME.io_diffCommits_info_283_pdest = RTL_PATH.io_diffCommits_info_283_pdest; \
        force U_IF_NAME.io_diffCommits_info_284_ldest = RTL_PATH.io_diffCommits_info_284_ldest; \
        force U_IF_NAME.io_diffCommits_info_284_pdest = RTL_PATH.io_diffCommits_info_284_pdest; \
        force U_IF_NAME.io_diffCommits_info_285_ldest = RTL_PATH.io_diffCommits_info_285_ldest; \
        force U_IF_NAME.io_diffCommits_info_285_pdest = RTL_PATH.io_diffCommits_info_285_pdest; \
        force U_IF_NAME.io_diffCommits_info_286_ldest = RTL_PATH.io_diffCommits_info_286_ldest; \
        force U_IF_NAME.io_diffCommits_info_286_pdest = RTL_PATH.io_diffCommits_info_286_pdest; \
        force U_IF_NAME.io_diffCommits_info_287_ldest = RTL_PATH.io_diffCommits_info_287_ldest; \
        force U_IF_NAME.io_diffCommits_info_287_pdest = RTL_PATH.io_diffCommits_info_287_pdest; \
        force U_IF_NAME.io_diffCommits_info_288_ldest = RTL_PATH.io_diffCommits_info_288_ldest; \
        force U_IF_NAME.io_diffCommits_info_288_pdest = RTL_PATH.io_diffCommits_info_288_pdest; \
        force U_IF_NAME.io_diffCommits_info_289_ldest = RTL_PATH.io_diffCommits_info_289_ldest; \
        force U_IF_NAME.io_diffCommits_info_289_pdest = RTL_PATH.io_diffCommits_info_289_pdest; \
        force U_IF_NAME.io_diffCommits_info_290_ldest = RTL_PATH.io_diffCommits_info_290_ldest; \
        force U_IF_NAME.io_diffCommits_info_290_pdest = RTL_PATH.io_diffCommits_info_290_pdest; \
        force U_IF_NAME.io_diffCommits_info_291_ldest = RTL_PATH.io_diffCommits_info_291_ldest; \
        force U_IF_NAME.io_diffCommits_info_291_pdest = RTL_PATH.io_diffCommits_info_291_pdest; \
        force U_IF_NAME.io_diffCommits_info_292_ldest = RTL_PATH.io_diffCommits_info_292_ldest; \
        force U_IF_NAME.io_diffCommits_info_292_pdest = RTL_PATH.io_diffCommits_info_292_pdest; \
        force U_IF_NAME.io_diffCommits_info_293_ldest = RTL_PATH.io_diffCommits_info_293_ldest; \
        force U_IF_NAME.io_diffCommits_info_293_pdest = RTL_PATH.io_diffCommits_info_293_pdest; \
        force U_IF_NAME.io_diffCommits_info_294_ldest = RTL_PATH.io_diffCommits_info_294_ldest; \
        force U_IF_NAME.io_diffCommits_info_294_pdest = RTL_PATH.io_diffCommits_info_294_pdest; \
        force U_IF_NAME.io_diffCommits_info_295_ldest = RTL_PATH.io_diffCommits_info_295_ldest; \
        force U_IF_NAME.io_diffCommits_info_295_pdest = RTL_PATH.io_diffCommits_info_295_pdest; \
        force U_IF_NAME.io_diffCommits_info_296_ldest = RTL_PATH.io_diffCommits_info_296_ldest; \
        force U_IF_NAME.io_diffCommits_info_296_pdest = RTL_PATH.io_diffCommits_info_296_pdest; \
        force U_IF_NAME.io_diffCommits_info_297_ldest = RTL_PATH.io_diffCommits_info_297_ldest; \
        force U_IF_NAME.io_diffCommits_info_297_pdest = RTL_PATH.io_diffCommits_info_297_pdest; \
        force U_IF_NAME.io_diffCommits_info_298_ldest = RTL_PATH.io_diffCommits_info_298_ldest; \
        force U_IF_NAME.io_diffCommits_info_298_pdest = RTL_PATH.io_diffCommits_info_298_pdest; \
        force U_IF_NAME.io_diffCommits_info_299_ldest = RTL_PATH.io_diffCommits_info_299_ldest; \
        force U_IF_NAME.io_diffCommits_info_299_pdest = RTL_PATH.io_diffCommits_info_299_pdest; \
        force U_IF_NAME.io_diffCommits_info_300_ldest = RTL_PATH.io_diffCommits_info_300_ldest; \
        force U_IF_NAME.io_diffCommits_info_300_pdest = RTL_PATH.io_diffCommits_info_300_pdest; \
        force U_IF_NAME.io_diffCommits_info_301_ldest = RTL_PATH.io_diffCommits_info_301_ldest; \
        force U_IF_NAME.io_diffCommits_info_301_pdest = RTL_PATH.io_diffCommits_info_301_pdest; \
        force U_IF_NAME.io_diffCommits_info_302_ldest = RTL_PATH.io_diffCommits_info_302_ldest; \
        force U_IF_NAME.io_diffCommits_info_302_pdest = RTL_PATH.io_diffCommits_info_302_pdest; \
        force U_IF_NAME.io_diffCommits_info_303_ldest = RTL_PATH.io_diffCommits_info_303_ldest; \
        force U_IF_NAME.io_diffCommits_info_303_pdest = RTL_PATH.io_diffCommits_info_303_pdest; \
        force U_IF_NAME.io_diffCommits_info_304_ldest = RTL_PATH.io_diffCommits_info_304_ldest; \
        force U_IF_NAME.io_diffCommits_info_304_pdest = RTL_PATH.io_diffCommits_info_304_pdest; \
        force U_IF_NAME.io_diffCommits_info_305_ldest = RTL_PATH.io_diffCommits_info_305_ldest; \
        force U_IF_NAME.io_diffCommits_info_305_pdest = RTL_PATH.io_diffCommits_info_305_pdest; \
        force U_IF_NAME.io_diffCommits_info_306_ldest = RTL_PATH.io_diffCommits_info_306_ldest; \
        force U_IF_NAME.io_diffCommits_info_306_pdest = RTL_PATH.io_diffCommits_info_306_pdest; \
        force U_IF_NAME.io_diffCommits_info_307_ldest = RTL_PATH.io_diffCommits_info_307_ldest; \
        force U_IF_NAME.io_diffCommits_info_307_pdest = RTL_PATH.io_diffCommits_info_307_pdest; \
        force U_IF_NAME.io_diffCommits_info_308_ldest = RTL_PATH.io_diffCommits_info_308_ldest; \
        force U_IF_NAME.io_diffCommits_info_308_pdest = RTL_PATH.io_diffCommits_info_308_pdest; \
        force U_IF_NAME.io_diffCommits_info_309_ldest = RTL_PATH.io_diffCommits_info_309_ldest; \
        force U_IF_NAME.io_diffCommits_info_309_pdest = RTL_PATH.io_diffCommits_info_309_pdest; \
        force U_IF_NAME.io_diffCommits_info_310_ldest = RTL_PATH.io_diffCommits_info_310_ldest; \
        force U_IF_NAME.io_diffCommits_info_310_pdest = RTL_PATH.io_diffCommits_info_310_pdest; \
        force U_IF_NAME.io_diffCommits_info_311_ldest = RTL_PATH.io_diffCommits_info_311_ldest; \
        force U_IF_NAME.io_diffCommits_info_311_pdest = RTL_PATH.io_diffCommits_info_311_pdest; \
        force U_IF_NAME.io_diffCommits_info_312_ldest = RTL_PATH.io_diffCommits_info_312_ldest; \
        force U_IF_NAME.io_diffCommits_info_312_pdest = RTL_PATH.io_diffCommits_info_312_pdest; \
        force U_IF_NAME.io_diffCommits_info_313_ldest = RTL_PATH.io_diffCommits_info_313_ldest; \
        force U_IF_NAME.io_diffCommits_info_313_pdest = RTL_PATH.io_diffCommits_info_313_pdest; \
        force U_IF_NAME.io_diffCommits_info_314_ldest = RTL_PATH.io_diffCommits_info_314_ldest; \
        force U_IF_NAME.io_diffCommits_info_314_pdest = RTL_PATH.io_diffCommits_info_314_pdest; \
        force U_IF_NAME.io_diffCommits_info_315_ldest = RTL_PATH.io_diffCommits_info_315_ldest; \
        force U_IF_NAME.io_diffCommits_info_315_pdest = RTL_PATH.io_diffCommits_info_315_pdest; \
        force U_IF_NAME.io_diffCommits_info_316_ldest = RTL_PATH.io_diffCommits_info_316_ldest; \
        force U_IF_NAME.io_diffCommits_info_316_pdest = RTL_PATH.io_diffCommits_info_316_pdest; \
        force U_IF_NAME.io_diffCommits_info_317_ldest = RTL_PATH.io_diffCommits_info_317_ldest; \
        force U_IF_NAME.io_diffCommits_info_317_pdest = RTL_PATH.io_diffCommits_info_317_pdest; \
        force U_IF_NAME.io_diffCommits_info_318_ldest = RTL_PATH.io_diffCommits_info_318_ldest; \
        force U_IF_NAME.io_diffCommits_info_318_pdest = RTL_PATH.io_diffCommits_info_318_pdest; \
        force U_IF_NAME.io_diffCommits_info_319_ldest = RTL_PATH.io_diffCommits_info_319_ldest; \
        force U_IF_NAME.io_diffCommits_info_319_pdest = RTL_PATH.io_diffCommits_info_319_pdest; \
        force U_IF_NAME.io_diffCommits_info_320_ldest = RTL_PATH.io_diffCommits_info_320_ldest; \
        force U_IF_NAME.io_diffCommits_info_320_pdest = RTL_PATH.io_diffCommits_info_320_pdest; \
        force U_IF_NAME.io_diffCommits_info_321_ldest = RTL_PATH.io_diffCommits_info_321_ldest; \
        force U_IF_NAME.io_diffCommits_info_321_pdest = RTL_PATH.io_diffCommits_info_321_pdest; \
        force U_IF_NAME.io_diffCommits_info_322_ldest = RTL_PATH.io_diffCommits_info_322_ldest; \
        force U_IF_NAME.io_diffCommits_info_322_pdest = RTL_PATH.io_diffCommits_info_322_pdest; \
        force U_IF_NAME.io_diffCommits_info_323_ldest = RTL_PATH.io_diffCommits_info_323_ldest; \
        force U_IF_NAME.io_diffCommits_info_323_pdest = RTL_PATH.io_diffCommits_info_323_pdest; \
        force U_IF_NAME.io_diffCommits_info_324_ldest = RTL_PATH.io_diffCommits_info_324_ldest; \
        force U_IF_NAME.io_diffCommits_info_324_pdest = RTL_PATH.io_diffCommits_info_324_pdest; \
        force U_IF_NAME.io_diffCommits_info_325_ldest = RTL_PATH.io_diffCommits_info_325_ldest; \
        force U_IF_NAME.io_diffCommits_info_325_pdest = RTL_PATH.io_diffCommits_info_325_pdest; \
        force U_IF_NAME.io_diffCommits_info_326_ldest = RTL_PATH.io_diffCommits_info_326_ldest; \
        force U_IF_NAME.io_diffCommits_info_326_pdest = RTL_PATH.io_diffCommits_info_326_pdest; \
        force U_IF_NAME.io_diffCommits_info_327_ldest = RTL_PATH.io_diffCommits_info_327_ldest; \
        force U_IF_NAME.io_diffCommits_info_327_pdest = RTL_PATH.io_diffCommits_info_327_pdest; \
        force U_IF_NAME.io_diffCommits_info_328_ldest = RTL_PATH.io_diffCommits_info_328_ldest; \
        force U_IF_NAME.io_diffCommits_info_328_pdest = RTL_PATH.io_diffCommits_info_328_pdest; \
        force U_IF_NAME.io_diffCommits_info_329_ldest = RTL_PATH.io_diffCommits_info_329_ldest; \
        force U_IF_NAME.io_diffCommits_info_329_pdest = RTL_PATH.io_diffCommits_info_329_pdest; \
        force U_IF_NAME.io_diffCommits_info_330_ldest = RTL_PATH.io_diffCommits_info_330_ldest; \
        force U_IF_NAME.io_diffCommits_info_330_pdest = RTL_PATH.io_diffCommits_info_330_pdest; \
        force U_IF_NAME.io_diffCommits_info_331_ldest = RTL_PATH.io_diffCommits_info_331_ldest; \
        force U_IF_NAME.io_diffCommits_info_331_pdest = RTL_PATH.io_diffCommits_info_331_pdest; \
        force U_IF_NAME.io_diffCommits_info_332_ldest = RTL_PATH.io_diffCommits_info_332_ldest; \
        force U_IF_NAME.io_diffCommits_info_332_pdest = RTL_PATH.io_diffCommits_info_332_pdest; \
        force U_IF_NAME.io_diffCommits_info_333_ldest = RTL_PATH.io_diffCommits_info_333_ldest; \
        force U_IF_NAME.io_diffCommits_info_333_pdest = RTL_PATH.io_diffCommits_info_333_pdest; \
        force U_IF_NAME.io_diffCommits_info_334_ldest = RTL_PATH.io_diffCommits_info_334_ldest; \
        force U_IF_NAME.io_diffCommits_info_334_pdest = RTL_PATH.io_diffCommits_info_334_pdest; \
        force U_IF_NAME.io_diffCommits_info_335_ldest = RTL_PATH.io_diffCommits_info_335_ldest; \
        force U_IF_NAME.io_diffCommits_info_335_pdest = RTL_PATH.io_diffCommits_info_335_pdest; \
        force U_IF_NAME.io_diffCommits_info_336_ldest = RTL_PATH.io_diffCommits_info_336_ldest; \
        force U_IF_NAME.io_diffCommits_info_336_pdest = RTL_PATH.io_diffCommits_info_336_pdest; \
        force U_IF_NAME.io_diffCommits_info_337_ldest = RTL_PATH.io_diffCommits_info_337_ldest; \
        force U_IF_NAME.io_diffCommits_info_337_pdest = RTL_PATH.io_diffCommits_info_337_pdest; \
        force U_IF_NAME.io_diffCommits_info_338_ldest = RTL_PATH.io_diffCommits_info_338_ldest; \
        force U_IF_NAME.io_diffCommits_info_338_pdest = RTL_PATH.io_diffCommits_info_338_pdest; \
        force U_IF_NAME.io_diffCommits_info_339_ldest = RTL_PATH.io_diffCommits_info_339_ldest; \
        force U_IF_NAME.io_diffCommits_info_339_pdest = RTL_PATH.io_diffCommits_info_339_pdest; \
        force U_IF_NAME.io_diffCommits_info_340_ldest = RTL_PATH.io_diffCommits_info_340_ldest; \
        force U_IF_NAME.io_diffCommits_info_340_pdest = RTL_PATH.io_diffCommits_info_340_pdest; \
        force U_IF_NAME.io_diffCommits_info_341_ldest = RTL_PATH.io_diffCommits_info_341_ldest; \
        force U_IF_NAME.io_diffCommits_info_341_pdest = RTL_PATH.io_diffCommits_info_341_pdest; \
        force U_IF_NAME.io_diffCommits_info_342_ldest = RTL_PATH.io_diffCommits_info_342_ldest; \
        force U_IF_NAME.io_diffCommits_info_342_pdest = RTL_PATH.io_diffCommits_info_342_pdest; \
        force U_IF_NAME.io_diffCommits_info_343_ldest = RTL_PATH.io_diffCommits_info_343_ldest; \
        force U_IF_NAME.io_diffCommits_info_343_pdest = RTL_PATH.io_diffCommits_info_343_pdest; \
        force U_IF_NAME.io_diffCommits_info_344_ldest = RTL_PATH.io_diffCommits_info_344_ldest; \
        force U_IF_NAME.io_diffCommits_info_344_pdest = RTL_PATH.io_diffCommits_info_344_pdest; \
        force U_IF_NAME.io_diffCommits_info_345_ldest = RTL_PATH.io_diffCommits_info_345_ldest; \
        force U_IF_NAME.io_diffCommits_info_345_pdest = RTL_PATH.io_diffCommits_info_345_pdest; \
        force U_IF_NAME.io_diffCommits_info_346_ldest = RTL_PATH.io_diffCommits_info_346_ldest; \
        force U_IF_NAME.io_diffCommits_info_346_pdest = RTL_PATH.io_diffCommits_info_346_pdest; \
        force U_IF_NAME.io_diffCommits_info_347_ldest = RTL_PATH.io_diffCommits_info_347_ldest; \
        force U_IF_NAME.io_diffCommits_info_347_pdest = RTL_PATH.io_diffCommits_info_347_pdest; \
        force U_IF_NAME.io_diffCommits_info_348_ldest = RTL_PATH.io_diffCommits_info_348_ldest; \
        force U_IF_NAME.io_diffCommits_info_348_pdest = RTL_PATH.io_diffCommits_info_348_pdest; \
        force U_IF_NAME.io_diffCommits_info_349_ldest = RTL_PATH.io_diffCommits_info_349_ldest; \
        force U_IF_NAME.io_diffCommits_info_349_pdest = RTL_PATH.io_diffCommits_info_349_pdest; \
        force U_IF_NAME.io_diffCommits_info_350_ldest = RTL_PATH.io_diffCommits_info_350_ldest; \
        force U_IF_NAME.io_diffCommits_info_350_pdest = RTL_PATH.io_diffCommits_info_350_pdest; \
        force U_IF_NAME.io_diffCommits_info_351_ldest = RTL_PATH.io_diffCommits_info_351_ldest; \
        force U_IF_NAME.io_diffCommits_info_351_pdest = RTL_PATH.io_diffCommits_info_351_pdest; \
        force U_IF_NAME.io_diffCommits_info_352_ldest = RTL_PATH.io_diffCommits_info_352_ldest; \
        force U_IF_NAME.io_diffCommits_info_352_pdest = RTL_PATH.io_diffCommits_info_352_pdest; \
        force U_IF_NAME.io_diffCommits_info_353_ldest = RTL_PATH.io_diffCommits_info_353_ldest; \
        force U_IF_NAME.io_diffCommits_info_353_pdest = RTL_PATH.io_diffCommits_info_353_pdest; \
        force U_IF_NAME.io_diffCommits_info_354_ldest = RTL_PATH.io_diffCommits_info_354_ldest; \
        force U_IF_NAME.io_diffCommits_info_354_pdest = RTL_PATH.io_diffCommits_info_354_pdest; \
        force U_IF_NAME.io_diffCommits_info_355_ldest = RTL_PATH.io_diffCommits_info_355_ldest; \
        force U_IF_NAME.io_diffCommits_info_355_pdest = RTL_PATH.io_diffCommits_info_355_pdest; \
        force U_IF_NAME.io_diffCommits_info_356_ldest = RTL_PATH.io_diffCommits_info_356_ldest; \
        force U_IF_NAME.io_diffCommits_info_356_pdest = RTL_PATH.io_diffCommits_info_356_pdest; \
        force U_IF_NAME.io_diffCommits_info_357_ldest = RTL_PATH.io_diffCommits_info_357_ldest; \
        force U_IF_NAME.io_diffCommits_info_357_pdest = RTL_PATH.io_diffCommits_info_357_pdest; \
        force U_IF_NAME.io_diffCommits_info_358_ldest = RTL_PATH.io_diffCommits_info_358_ldest; \
        force U_IF_NAME.io_diffCommits_info_358_pdest = RTL_PATH.io_diffCommits_info_358_pdest; \
        force U_IF_NAME.io_diffCommits_info_359_ldest = RTL_PATH.io_diffCommits_info_359_ldest; \
        force U_IF_NAME.io_diffCommits_info_359_pdest = RTL_PATH.io_diffCommits_info_359_pdest; \
        force U_IF_NAME.io_diffCommits_info_360_ldest = RTL_PATH.io_diffCommits_info_360_ldest; \
        force U_IF_NAME.io_diffCommits_info_360_pdest = RTL_PATH.io_diffCommits_info_360_pdest; \
        force U_IF_NAME.io_diffCommits_info_361_ldest = RTL_PATH.io_diffCommits_info_361_ldest; \
        force U_IF_NAME.io_diffCommits_info_361_pdest = RTL_PATH.io_diffCommits_info_361_pdest; \
        force U_IF_NAME.io_diffCommits_info_362_ldest = RTL_PATH.io_diffCommits_info_362_ldest; \
        force U_IF_NAME.io_diffCommits_info_362_pdest = RTL_PATH.io_diffCommits_info_362_pdest; \
        force U_IF_NAME.io_diffCommits_info_363_ldest = RTL_PATH.io_diffCommits_info_363_ldest; \
        force U_IF_NAME.io_diffCommits_info_363_pdest = RTL_PATH.io_diffCommits_info_363_pdest; \
        force U_IF_NAME.io_diffCommits_info_364_ldest = RTL_PATH.io_diffCommits_info_364_ldest; \
        force U_IF_NAME.io_diffCommits_info_364_pdest = RTL_PATH.io_diffCommits_info_364_pdest; \
        force U_IF_NAME.io_diffCommits_info_365_ldest = RTL_PATH.io_diffCommits_info_365_ldest; \
        force U_IF_NAME.io_diffCommits_info_365_pdest = RTL_PATH.io_diffCommits_info_365_pdest; \
        force U_IF_NAME.io_diffCommits_info_366_ldest = RTL_PATH.io_diffCommits_info_366_ldest; \
        force U_IF_NAME.io_diffCommits_info_366_pdest = RTL_PATH.io_diffCommits_info_366_pdest; \
        force U_IF_NAME.io_diffCommits_info_367_ldest = RTL_PATH.io_diffCommits_info_367_ldest; \
        force U_IF_NAME.io_diffCommits_info_367_pdest = RTL_PATH.io_diffCommits_info_367_pdest; \
        force U_IF_NAME.io_diffCommits_info_368_ldest = RTL_PATH.io_diffCommits_info_368_ldest; \
        force U_IF_NAME.io_diffCommits_info_368_pdest = RTL_PATH.io_diffCommits_info_368_pdest; \
        force U_IF_NAME.io_diffCommits_info_369_ldest = RTL_PATH.io_diffCommits_info_369_ldest; \
        force U_IF_NAME.io_diffCommits_info_369_pdest = RTL_PATH.io_diffCommits_info_369_pdest; \
        force U_IF_NAME.io_diffCommits_info_370_ldest = RTL_PATH.io_diffCommits_info_370_ldest; \
        force U_IF_NAME.io_diffCommits_info_370_pdest = RTL_PATH.io_diffCommits_info_370_pdest; \
        force U_IF_NAME.io_diffCommits_info_371_ldest = RTL_PATH.io_diffCommits_info_371_ldest; \
        force U_IF_NAME.io_diffCommits_info_371_pdest = RTL_PATH.io_diffCommits_info_371_pdest; \
        force U_IF_NAME.io_diffCommits_info_372_ldest = RTL_PATH.io_diffCommits_info_372_ldest; \
        force U_IF_NAME.io_diffCommits_info_372_pdest = RTL_PATH.io_diffCommits_info_372_pdest; \
        force U_IF_NAME.io_diffCommits_info_373_ldest = RTL_PATH.io_diffCommits_info_373_ldest; \
        force U_IF_NAME.io_diffCommits_info_373_pdest = RTL_PATH.io_diffCommits_info_373_pdest; \
        force U_IF_NAME.io_diffCommits_info_374_ldest = RTL_PATH.io_diffCommits_info_374_ldest; \
        force U_IF_NAME.io_diffCommits_info_374_pdest = RTL_PATH.io_diffCommits_info_374_pdest; \
        force U_IF_NAME.io_diffCommits_info_375_ldest = RTL_PATH.io_diffCommits_info_375_ldest; \
        force U_IF_NAME.io_diffCommits_info_375_pdest = RTL_PATH.io_diffCommits_info_375_pdest; \
        force U_IF_NAME.io_diffCommits_info_376_ldest = RTL_PATH.io_diffCommits_info_376_ldest; \
        force U_IF_NAME.io_diffCommits_info_376_pdest = RTL_PATH.io_diffCommits_info_376_pdest; \
        force U_IF_NAME.io_diffCommits_info_377_ldest = RTL_PATH.io_diffCommits_info_377_ldest; \
        force U_IF_NAME.io_diffCommits_info_377_pdest = RTL_PATH.io_diffCommits_info_377_pdest; \
        force U_IF_NAME.io_diffCommits_info_378_ldest = RTL_PATH.io_diffCommits_info_378_ldest; \
        force U_IF_NAME.io_diffCommits_info_378_pdest = RTL_PATH.io_diffCommits_info_378_pdest; \
        force U_IF_NAME.io_diffCommits_info_379_ldest = RTL_PATH.io_diffCommits_info_379_ldest; \
        force U_IF_NAME.io_diffCommits_info_379_pdest = RTL_PATH.io_diffCommits_info_379_pdest; \
        force U_IF_NAME.io_diffCommits_info_380_ldest = RTL_PATH.io_diffCommits_info_380_ldest; \
        force U_IF_NAME.io_diffCommits_info_380_pdest = RTL_PATH.io_diffCommits_info_380_pdest; \
        force U_IF_NAME.io_diffCommits_info_381_ldest = RTL_PATH.io_diffCommits_info_381_ldest; \
        force U_IF_NAME.io_diffCommits_info_381_pdest = RTL_PATH.io_diffCommits_info_381_pdest; \
        force U_IF_NAME.io_diffCommits_info_382_ldest = RTL_PATH.io_diffCommits_info_382_ldest; \
        force U_IF_NAME.io_diffCommits_info_382_pdest = RTL_PATH.io_diffCommits_info_382_pdest; \
        force U_IF_NAME.io_diffCommits_info_383_ldest = RTL_PATH.io_diffCommits_info_383_ldest; \
        force U_IF_NAME.io_diffCommits_info_383_pdest = RTL_PATH.io_diffCommits_info_383_pdest; \
        force U_IF_NAME.io_diffCommits_info_384_ldest = RTL_PATH.io_diffCommits_info_384_ldest; \
        force U_IF_NAME.io_diffCommits_info_384_pdest = RTL_PATH.io_diffCommits_info_384_pdest; \
        force U_IF_NAME.io_diffCommits_info_385_ldest = RTL_PATH.io_diffCommits_info_385_ldest; \
        force U_IF_NAME.io_diffCommits_info_385_pdest = RTL_PATH.io_diffCommits_info_385_pdest; \
        force U_IF_NAME.io_diffCommits_info_386_ldest = RTL_PATH.io_diffCommits_info_386_ldest; \
        force U_IF_NAME.io_diffCommits_info_386_pdest = RTL_PATH.io_diffCommits_info_386_pdest; \
        force U_IF_NAME.io_diffCommits_info_387_ldest = RTL_PATH.io_diffCommits_info_387_ldest; \
        force U_IF_NAME.io_diffCommits_info_387_pdest = RTL_PATH.io_diffCommits_info_387_pdest; \
        force U_IF_NAME.io_diffCommits_info_388_ldest = RTL_PATH.io_diffCommits_info_388_ldest; \
        force U_IF_NAME.io_diffCommits_info_388_pdest = RTL_PATH.io_diffCommits_info_388_pdest; \
        force U_IF_NAME.io_diffCommits_info_389_ldest = RTL_PATH.io_diffCommits_info_389_ldest; \
        force U_IF_NAME.io_diffCommits_info_389_pdest = RTL_PATH.io_diffCommits_info_389_pdest; \
        force U_IF_NAME.io_lsq_scommit = RTL_PATH.io_lsq_scommit; \
        force U_IF_NAME.io_lsq_pendingMMIOld = RTL_PATH.io_lsq_pendingMMIOld; \
        force U_IF_NAME.io_lsq_pendingst = RTL_PATH.io_lsq_pendingst; \
        force U_IF_NAME.io_lsq_pendingPtr_flag = RTL_PATH.io_lsq_pendingPtr_flag; \
        force U_IF_NAME.io_lsq_pendingPtr_value = RTL_PATH.io_lsq_pendingPtr_value; \
        force U_IF_NAME.io_robDeqPtr_flag = RTL_PATH.io_robDeqPtr_flag; \
        force U_IF_NAME.io_robDeqPtr_value = RTL_PATH.io_robDeqPtr_value; \
        force U_IF_NAME.io_csr_fflags_valid = RTL_PATH.io_csr_fflags_valid; \
        force U_IF_NAME.io_csr_fflags_bits = RTL_PATH.io_csr_fflags_bits; \
        force U_IF_NAME.io_csr_vxsat_valid = RTL_PATH.io_csr_vxsat_valid; \
        force U_IF_NAME.io_csr_vxsat_bits = RTL_PATH.io_csr_vxsat_bits; \
        force U_IF_NAME.io_csr_vstart_valid = RTL_PATH.io_csr_vstart_valid; \
        force U_IF_NAME.io_csr_vstart_bits = RTL_PATH.io_csr_vstart_bits; \
        force U_IF_NAME.io_csr_dirty_fs = RTL_PATH.io_csr_dirty_fs; \
        force U_IF_NAME.io_csr_dirty_vs = RTL_PATH.io_csr_dirty_vs; \
        force U_IF_NAME.io_csr_perfinfo_retiredInstr = RTL_PATH.io_csr_perfinfo_retiredInstr; \
        force U_IF_NAME.io_cpu_halt = RTL_PATH.io_cpu_halt; \
        force U_IF_NAME.io_wfi_wfiReq = RTL_PATH.io_wfi_wfiReq; \
        force U_IF_NAME.io_toDecode_isResumeVType = RTL_PATH.io_toDecode_isResumeVType; \
        force U_IF_NAME.io_toDecode_walkToArchVType = RTL_PATH.io_toDecode_walkToArchVType; \
        force U_IF_NAME.io_toDecode_walkVType_valid = RTL_PATH.io_toDecode_walkVType_valid; \
        force U_IF_NAME.io_toDecode_walkVType_bits_illegal = RTL_PATH.io_toDecode_walkVType_bits_illegal; \
        force U_IF_NAME.io_toDecode_walkVType_bits_vma = RTL_PATH.io_toDecode_walkVType_bits_vma; \
        force U_IF_NAME.io_toDecode_walkVType_bits_vta = RTL_PATH.io_toDecode_walkVType_bits_vta; \
        force U_IF_NAME.io_toDecode_walkVType_bits_vsew = RTL_PATH.io_toDecode_walkVType_bits_vsew; \
        force U_IF_NAME.io_toDecode_walkVType_bits_vlmul = RTL_PATH.io_toDecode_walkVType_bits_vlmul; \
        force U_IF_NAME.io_toDecode_commitVType_vtype_valid = RTL_PATH.io_toDecode_commitVType_vtype_valid; \
        force U_IF_NAME.io_toDecode_commitVType_vtype_bits_illegal = RTL_PATH.io_toDecode_commitVType_vtype_bits_illegal; \
        force U_IF_NAME.io_toDecode_commitVType_vtype_bits_vma = RTL_PATH.io_toDecode_commitVType_vtype_bits_vma; \
        force U_IF_NAME.io_toDecode_commitVType_vtype_bits_vta = RTL_PATH.io_toDecode_commitVType_vtype_bits_vta; \
        force U_IF_NAME.io_toDecode_commitVType_vtype_bits_vsew = RTL_PATH.io_toDecode_commitVType_vtype_bits_vsew; \
        force U_IF_NAME.io_toDecode_commitVType_vtype_bits_vlmul = RTL_PATH.io_toDecode_commitVType_vtype_bits_vlmul; \
        force U_IF_NAME.io_toDecode_commitVType_hasVsetvl = RTL_PATH.io_toDecode_commitVType_hasVsetvl; \
        force U_IF_NAME.io_readGPAMemAddr_valid = RTL_PATH.io_readGPAMemAddr_valid; \
        force U_IF_NAME.io_readGPAMemAddr_bits_ftqPtr_value = RTL_PATH.io_readGPAMemAddr_bits_ftqPtr_value; \
        force U_IF_NAME.io_readGPAMemAddr_bits_ftqOffset = RTL_PATH.io_readGPAMemAddr_bits_ftqOffset; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_0_valid = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_0_valid; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_0_bits_lreg = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_0_bits_lreg; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_0_bits_preg = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_0_bits_preg; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_1_valid = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_1_valid; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_1_bits_lreg = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_1_bits_lreg; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_1_bits_preg = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_1_bits_preg; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_2_valid = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_2_valid; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_2_bits_lreg = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_2_bits_lreg; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_2_bits_preg = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_2_bits_preg; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_3_valid = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_3_valid; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_3_bits_lreg = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_3_bits_lreg; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_3_bits_preg = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_3_bits_preg; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_4_valid = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_4_valid; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_4_bits_lreg = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_4_bits_lreg; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_4_bits_preg = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_4_bits_preg; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_5_valid = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_5_valid; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_5_bits_lreg = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_5_bits_lreg; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_5_bits_preg = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_5_bits_preg; \
        force U_IF_NAME.io_toVecExcpMod_excpInfo_valid = RTL_PATH.io_toVecExcpMod_excpInfo_valid; \
        force U_IF_NAME.io_toVecExcpMod_excpInfo_bits_vstart = RTL_PATH.io_toVecExcpMod_excpInfo_bits_vstart; \
        force U_IF_NAME.io_toVecExcpMod_excpInfo_bits_vsew = RTL_PATH.io_toVecExcpMod_excpInfo_bits_vsew; \
        force U_IF_NAME.io_toVecExcpMod_excpInfo_bits_veew = RTL_PATH.io_toVecExcpMod_excpInfo_bits_veew; \
        force U_IF_NAME.io_toVecExcpMod_excpInfo_bits_vlmul = RTL_PATH.io_toVecExcpMod_excpInfo_bits_vlmul; \
        force U_IF_NAME.io_toVecExcpMod_excpInfo_bits_nf = RTL_PATH.io_toVecExcpMod_excpInfo_bits_nf; \
        force U_IF_NAME.io_toVecExcpMod_excpInfo_bits_isStride = RTL_PATH.io_toVecExcpMod_excpInfo_bits_isStride; \
        force U_IF_NAME.io_toVecExcpMod_excpInfo_bits_isIndexed = RTL_PATH.io_toVecExcpMod_excpInfo_bits_isIndexed; \
        force U_IF_NAME.io_toVecExcpMod_excpInfo_bits_isWhole = RTL_PATH.io_toVecExcpMod_excpInfo_bits_isWhole; \
        force U_IF_NAME.io_toVecExcpMod_excpInfo_bits_isVlm = RTL_PATH.io_toVecExcpMod_excpInfo_bits_isVlm; \
        force U_IF_NAME.io_storeDebugInfo_1_pc = RTL_PATH.io_storeDebugInfo_1_pc; \
        force U_IF_NAME.io_perf_0_value = RTL_PATH.io_perf_0_value; \
        force U_IF_NAME.io_perf_1_value = RTL_PATH.io_perf_1_value; \
        force U_IF_NAME.io_perf_2_value = RTL_PATH.io_perf_2_value; \
        force U_IF_NAME.io_perf_3_value = RTL_PATH.io_perf_3_value; \
        force U_IF_NAME.io_perf_4_value = RTL_PATH.io_perf_4_value; \
        force U_IF_NAME.io_perf_5_value = RTL_PATH.io_perf_5_value; \
        force U_IF_NAME.io_perf_6_value = RTL_PATH.io_perf_6_value; \
        force U_IF_NAME.io_perf_7_value = RTL_PATH.io_perf_7_value; \
        force U_IF_NAME.io_perf_8_value = RTL_PATH.io_perf_8_value; \
        force U_IF_NAME.io_perf_9_value = RTL_PATH.io_perf_9_value; \
        force U_IF_NAME.io_perf_10_value = RTL_PATH.io_perf_10_value; \
        force U_IF_NAME.io_perf_11_value = RTL_PATH.io_perf_11_value; \
        force U_IF_NAME.io_perf_12_value = RTL_PATH.io_perf_12_value; \
        force U_IF_NAME.io_perf_13_value = RTL_PATH.io_perf_13_value; \
        force U_IF_NAME.io_perf_14_value = RTL_PATH.io_perf_14_value; \
        force U_IF_NAME.io_perf_15_value = RTL_PATH.io_perf_15_value; \
        force U_IF_NAME.io_perf_16_value = RTL_PATH.io_perf_16_value; \
        force U_IF_NAME.io_perf_17_value = RTL_PATH.io_perf_17_value; \
        force U_IF_NAME.io_error_0 = RTL_PATH.io_error_0; \
    end \
    `else \
    initial begin \
        force U_IF_NAME.io_enq_canAccept = RTL_PATH.io_enq_canAccept; \
        force U_IF_NAME.io_enq_canAcceptForDispatch = RTL_PATH.io_enq_canAcceptForDispatch; \
        force U_IF_NAME.io_enq_isEmpty = RTL_PATH.io_enq_isEmpty; \
        force U_IF_NAME.io_flushOut_valid = RTL_PATH.io_flushOut_valid; \
        force U_IF_NAME.io_flushOut_bits_isRVC = RTL_PATH.io_flushOut_bits_isRVC; \
        force U_IF_NAME.io_flushOut_bits_robIdx_flag = RTL_PATH.io_flushOut_bits_robIdx_flag; \
        force U_IF_NAME.io_flushOut_bits_robIdx_value = RTL_PATH.io_flushOut_bits_robIdx_value; \
        force U_IF_NAME.io_flushOut_bits_ftqIdx_flag = RTL_PATH.io_flushOut_bits_ftqIdx_flag; \
        force U_IF_NAME.io_flushOut_bits_ftqIdx_value = RTL_PATH.io_flushOut_bits_ftqIdx_value; \
        force U_IF_NAME.io_flushOut_bits_ftqOffset = RTL_PATH.io_flushOut_bits_ftqOffset; \
        force U_IF_NAME.io_flushOut_bits_level = RTL_PATH.io_flushOut_bits_level; \
        force U_IF_NAME.io_exception_valid = RTL_PATH.io_exception_valid; \
        force U_IF_NAME.io_exception_bits_instr = RTL_PATH.io_exception_bits_instr; \
        force U_IF_NAME.io_exception_bits_commitType = RTL_PATH.io_exception_bits_commitType; \
        force U_IF_NAME.io_exception_bits_exceptionVec_0 = RTL_PATH.io_exception_bits_exceptionVec_0; \
        force U_IF_NAME.io_exception_bits_exceptionVec_1 = RTL_PATH.io_exception_bits_exceptionVec_1; \
        force U_IF_NAME.io_exception_bits_exceptionVec_2 = RTL_PATH.io_exception_bits_exceptionVec_2; \
        force U_IF_NAME.io_exception_bits_exceptionVec_3 = RTL_PATH.io_exception_bits_exceptionVec_3; \
        force U_IF_NAME.io_exception_bits_exceptionVec_4 = RTL_PATH.io_exception_bits_exceptionVec_4; \
        force U_IF_NAME.io_exception_bits_exceptionVec_5 = RTL_PATH.io_exception_bits_exceptionVec_5; \
        force U_IF_NAME.io_exception_bits_exceptionVec_6 = RTL_PATH.io_exception_bits_exceptionVec_6; \
        force U_IF_NAME.io_exception_bits_exceptionVec_7 = RTL_PATH.io_exception_bits_exceptionVec_7; \
        force U_IF_NAME.io_exception_bits_exceptionVec_8 = RTL_PATH.io_exception_bits_exceptionVec_8; \
        force U_IF_NAME.io_exception_bits_exceptionVec_9 = RTL_PATH.io_exception_bits_exceptionVec_9; \
        force U_IF_NAME.io_exception_bits_exceptionVec_10 = RTL_PATH.io_exception_bits_exceptionVec_10; \
        force U_IF_NAME.io_exception_bits_exceptionVec_11 = RTL_PATH.io_exception_bits_exceptionVec_11; \
        force U_IF_NAME.io_exception_bits_exceptionVec_12 = RTL_PATH.io_exception_bits_exceptionVec_12; \
        force U_IF_NAME.io_exception_bits_exceptionVec_13 = RTL_PATH.io_exception_bits_exceptionVec_13; \
        force U_IF_NAME.io_exception_bits_exceptionVec_14 = RTL_PATH.io_exception_bits_exceptionVec_14; \
        force U_IF_NAME.io_exception_bits_exceptionVec_15 = RTL_PATH.io_exception_bits_exceptionVec_15; \
        force U_IF_NAME.io_exception_bits_exceptionVec_16 = RTL_PATH.io_exception_bits_exceptionVec_16; \
        force U_IF_NAME.io_exception_bits_exceptionVec_17 = RTL_PATH.io_exception_bits_exceptionVec_17; \
        force U_IF_NAME.io_exception_bits_exceptionVec_18 = RTL_PATH.io_exception_bits_exceptionVec_18; \
        force U_IF_NAME.io_exception_bits_exceptionVec_19 = RTL_PATH.io_exception_bits_exceptionVec_19; \
        force U_IF_NAME.io_exception_bits_exceptionVec_20 = RTL_PATH.io_exception_bits_exceptionVec_20; \
        force U_IF_NAME.io_exception_bits_exceptionVec_21 = RTL_PATH.io_exception_bits_exceptionVec_21; \
        force U_IF_NAME.io_exception_bits_exceptionVec_22 = RTL_PATH.io_exception_bits_exceptionVec_22; \
        force U_IF_NAME.io_exception_bits_exceptionVec_23 = RTL_PATH.io_exception_bits_exceptionVec_23; \
        force U_IF_NAME.io_exception_bits_isPcBkpt = RTL_PATH.io_exception_bits_isPcBkpt; \
        force U_IF_NAME.io_exception_bits_isFetchMalAddr = RTL_PATH.io_exception_bits_isFetchMalAddr; \
        force U_IF_NAME.io_exception_bits_gpaddr = RTL_PATH.io_exception_bits_gpaddr; \
        force U_IF_NAME.io_exception_bits_singleStep = RTL_PATH.io_exception_bits_singleStep; \
        force U_IF_NAME.io_exception_bits_crossPageIPFFix = RTL_PATH.io_exception_bits_crossPageIPFFix; \
        force U_IF_NAME.io_exception_bits_isInterrupt = RTL_PATH.io_exception_bits_isInterrupt; \
        force U_IF_NAME.io_exception_bits_isHls = RTL_PATH.io_exception_bits_isHls; \
        force U_IF_NAME.io_exception_bits_trigger = RTL_PATH.io_exception_bits_trigger; \
        force U_IF_NAME.io_exception_bits_isForVSnonLeafPTE = RTL_PATH.io_exception_bits_isForVSnonLeafPTE; \
        force U_IF_NAME.io_commits_isCommit = RTL_PATH.io_commits_isCommit; \
        force U_IF_NAME.io_commits_commitValid_0 = RTL_PATH.io_commits_commitValid_0; \
        force U_IF_NAME.io_commits_commitValid_1 = RTL_PATH.io_commits_commitValid_1; \
        force U_IF_NAME.io_commits_commitValid_2 = RTL_PATH.io_commits_commitValid_2; \
        force U_IF_NAME.io_commits_commitValid_3 = RTL_PATH.io_commits_commitValid_3; \
        force U_IF_NAME.io_commits_commitValid_4 = RTL_PATH.io_commits_commitValid_4; \
        force U_IF_NAME.io_commits_commitValid_5 = RTL_PATH.io_commits_commitValid_5; \
        force U_IF_NAME.io_commits_commitValid_6 = RTL_PATH.io_commits_commitValid_6; \
        force U_IF_NAME.io_commits_commitValid_7 = RTL_PATH.io_commits_commitValid_7; \
        force U_IF_NAME.io_commits_isWalk = RTL_PATH.io_commits_isWalk; \
        force U_IF_NAME.io_commits_walkValid_0 = RTL_PATH.io_commits_walkValid_0; \
        force U_IF_NAME.io_commits_walkValid_1 = RTL_PATH.io_commits_walkValid_1; \
        force U_IF_NAME.io_commits_walkValid_2 = RTL_PATH.io_commits_walkValid_2; \
        force U_IF_NAME.io_commits_walkValid_3 = RTL_PATH.io_commits_walkValid_3; \
        force U_IF_NAME.io_commits_walkValid_4 = RTL_PATH.io_commits_walkValid_4; \
        force U_IF_NAME.io_commits_walkValid_5 = RTL_PATH.io_commits_walkValid_5; \
        force U_IF_NAME.io_commits_walkValid_6 = RTL_PATH.io_commits_walkValid_6; \
        force U_IF_NAME.io_commits_walkValid_7 = RTL_PATH.io_commits_walkValid_7; \
        force U_IF_NAME.io_commits_info_0_walk_v = RTL_PATH.io_commits_info_0_walk_v; \
        force U_IF_NAME.io_commits_info_0_commit_v = RTL_PATH.io_commits_info_0_commit_v; \
        force U_IF_NAME.io_commits_info_0_commit_w = RTL_PATH.io_commits_info_0_commit_w; \
        force U_IF_NAME.io_commits_info_0_realDestSize = RTL_PATH.io_commits_info_0_realDestSize; \
        force U_IF_NAME.io_commits_info_0_interrupt_safe = RTL_PATH.io_commits_info_0_interrupt_safe; \
        force U_IF_NAME.io_commits_info_0_wflags = RTL_PATH.io_commits_info_0_wflags; \
        force U_IF_NAME.io_commits_info_0_fflags = RTL_PATH.io_commits_info_0_fflags; \
        force U_IF_NAME.io_commits_info_0_vxsat = RTL_PATH.io_commits_info_0_vxsat; \
        force U_IF_NAME.io_commits_info_0_isRVC = RTL_PATH.io_commits_info_0_isRVC; \
        force U_IF_NAME.io_commits_info_0_isVset = RTL_PATH.io_commits_info_0_isVset; \
        force U_IF_NAME.io_commits_info_0_isHls = RTL_PATH.io_commits_info_0_isHls; \
        force U_IF_NAME.io_commits_info_0_isVls = RTL_PATH.io_commits_info_0_isVls; \
        force U_IF_NAME.io_commits_info_0_vls = RTL_PATH.io_commits_info_0_vls; \
        force U_IF_NAME.io_commits_info_0_mmio = RTL_PATH.io_commits_info_0_mmio; \
        force U_IF_NAME.io_commits_info_0_commitType = RTL_PATH.io_commits_info_0_commitType; \
        force U_IF_NAME.io_commits_info_0_ftqIdx_flag = RTL_PATH.io_commits_info_0_ftqIdx_flag; \
        force U_IF_NAME.io_commits_info_0_ftqIdx_value = RTL_PATH.io_commits_info_0_ftqIdx_value; \
        force U_IF_NAME.io_commits_info_0_ftqOffset = RTL_PATH.io_commits_info_0_ftqOffset; \
        force U_IF_NAME.io_commits_info_0_instrSize = RTL_PATH.io_commits_info_0_instrSize; \
        force U_IF_NAME.io_commits_info_0_fpWen = RTL_PATH.io_commits_info_0_fpWen; \
        force U_IF_NAME.io_commits_info_0_rfWen = RTL_PATH.io_commits_info_0_rfWen; \
        force U_IF_NAME.io_commits_info_0_needFlush = RTL_PATH.io_commits_info_0_needFlush; \
        force U_IF_NAME.io_commits_info_0_traceBlockInPipe_itype = RTL_PATH.io_commits_info_0_traceBlockInPipe_itype; \
        force U_IF_NAME.io_commits_info_0_traceBlockInPipe_iretire = RTL_PATH.io_commits_info_0_traceBlockInPipe_iretire; \
        force U_IF_NAME.io_commits_info_0_traceBlockInPipe_ilastsize = RTL_PATH.io_commits_info_0_traceBlockInPipe_ilastsize; \
        force U_IF_NAME.io_commits_info_0_debug_pc = RTL_PATH.io_commits_info_0_debug_pc; \
        force U_IF_NAME.io_commits_info_0_debug_instr = RTL_PATH.io_commits_info_0_debug_instr; \
        force U_IF_NAME.io_commits_info_0_debug_ldest = RTL_PATH.io_commits_info_0_debug_ldest; \
        force U_IF_NAME.io_commits_info_0_debug_pdest = RTL_PATH.io_commits_info_0_debug_pdest; \
        force U_IF_NAME.io_commits_info_0_debug_otherPdest_0 = RTL_PATH.io_commits_info_0_debug_otherPdest_0; \
        force U_IF_NAME.io_commits_info_0_debug_otherPdest_1 = RTL_PATH.io_commits_info_0_debug_otherPdest_1; \
        force U_IF_NAME.io_commits_info_0_debug_otherPdest_2 = RTL_PATH.io_commits_info_0_debug_otherPdest_2; \
        force U_IF_NAME.io_commits_info_0_debug_otherPdest_3 = RTL_PATH.io_commits_info_0_debug_otherPdest_3; \
        force U_IF_NAME.io_commits_info_0_debug_otherPdest_4 = RTL_PATH.io_commits_info_0_debug_otherPdest_4; \
        force U_IF_NAME.io_commits_info_0_debug_otherPdest_5 = RTL_PATH.io_commits_info_0_debug_otherPdest_5; \
        force U_IF_NAME.io_commits_info_0_debug_otherPdest_6 = RTL_PATH.io_commits_info_0_debug_otherPdest_6; \
        force U_IF_NAME.io_commits_info_0_debug_fuType = RTL_PATH.io_commits_info_0_debug_fuType; \
        force U_IF_NAME.io_commits_info_0_dirtyFs = RTL_PATH.io_commits_info_0_dirtyFs; \
        force U_IF_NAME.io_commits_info_0_dirtyVs = RTL_PATH.io_commits_info_0_dirtyVs; \
        force U_IF_NAME.io_commits_info_1_walk_v = RTL_PATH.io_commits_info_1_walk_v; \
        force U_IF_NAME.io_commits_info_1_commit_v = RTL_PATH.io_commits_info_1_commit_v; \
        force U_IF_NAME.io_commits_info_1_commit_w = RTL_PATH.io_commits_info_1_commit_w; \
        force U_IF_NAME.io_commits_info_1_realDestSize = RTL_PATH.io_commits_info_1_realDestSize; \
        force U_IF_NAME.io_commits_info_1_interrupt_safe = RTL_PATH.io_commits_info_1_interrupt_safe; \
        force U_IF_NAME.io_commits_info_1_wflags = RTL_PATH.io_commits_info_1_wflags; \
        force U_IF_NAME.io_commits_info_1_fflags = RTL_PATH.io_commits_info_1_fflags; \
        force U_IF_NAME.io_commits_info_1_vxsat = RTL_PATH.io_commits_info_1_vxsat; \
        force U_IF_NAME.io_commits_info_1_isRVC = RTL_PATH.io_commits_info_1_isRVC; \
        force U_IF_NAME.io_commits_info_1_isVset = RTL_PATH.io_commits_info_1_isVset; \
        force U_IF_NAME.io_commits_info_1_isHls = RTL_PATH.io_commits_info_1_isHls; \
        force U_IF_NAME.io_commits_info_1_isVls = RTL_PATH.io_commits_info_1_isVls; \
        force U_IF_NAME.io_commits_info_1_vls = RTL_PATH.io_commits_info_1_vls; \
        force U_IF_NAME.io_commits_info_1_mmio = RTL_PATH.io_commits_info_1_mmio; \
        force U_IF_NAME.io_commits_info_1_commitType = RTL_PATH.io_commits_info_1_commitType; \
        force U_IF_NAME.io_commits_info_1_ftqIdx_flag = RTL_PATH.io_commits_info_1_ftqIdx_flag; \
        force U_IF_NAME.io_commits_info_1_ftqIdx_value = RTL_PATH.io_commits_info_1_ftqIdx_value; \
        force U_IF_NAME.io_commits_info_1_ftqOffset = RTL_PATH.io_commits_info_1_ftqOffset; \
        force U_IF_NAME.io_commits_info_1_instrSize = RTL_PATH.io_commits_info_1_instrSize; \
        force U_IF_NAME.io_commits_info_1_fpWen = RTL_PATH.io_commits_info_1_fpWen; \
        force U_IF_NAME.io_commits_info_1_rfWen = RTL_PATH.io_commits_info_1_rfWen; \
        force U_IF_NAME.io_commits_info_1_needFlush = RTL_PATH.io_commits_info_1_needFlush; \
        force U_IF_NAME.io_commits_info_1_traceBlockInPipe_itype = RTL_PATH.io_commits_info_1_traceBlockInPipe_itype; \
        force U_IF_NAME.io_commits_info_1_traceBlockInPipe_iretire = RTL_PATH.io_commits_info_1_traceBlockInPipe_iretire; \
        force U_IF_NAME.io_commits_info_1_traceBlockInPipe_ilastsize = RTL_PATH.io_commits_info_1_traceBlockInPipe_ilastsize; \
        force U_IF_NAME.io_commits_info_1_debug_pc = RTL_PATH.io_commits_info_1_debug_pc; \
        force U_IF_NAME.io_commits_info_1_debug_instr = RTL_PATH.io_commits_info_1_debug_instr; \
        force U_IF_NAME.io_commits_info_1_debug_ldest = RTL_PATH.io_commits_info_1_debug_ldest; \
        force U_IF_NAME.io_commits_info_1_debug_pdest = RTL_PATH.io_commits_info_1_debug_pdest; \
        force U_IF_NAME.io_commits_info_1_debug_otherPdest_0 = RTL_PATH.io_commits_info_1_debug_otherPdest_0; \
        force U_IF_NAME.io_commits_info_1_debug_otherPdest_1 = RTL_PATH.io_commits_info_1_debug_otherPdest_1; \
        force U_IF_NAME.io_commits_info_1_debug_otherPdest_2 = RTL_PATH.io_commits_info_1_debug_otherPdest_2; \
        force U_IF_NAME.io_commits_info_1_debug_otherPdest_3 = RTL_PATH.io_commits_info_1_debug_otherPdest_3; \
        force U_IF_NAME.io_commits_info_1_debug_otherPdest_4 = RTL_PATH.io_commits_info_1_debug_otherPdest_4; \
        force U_IF_NAME.io_commits_info_1_debug_otherPdest_5 = RTL_PATH.io_commits_info_1_debug_otherPdest_5; \
        force U_IF_NAME.io_commits_info_1_debug_otherPdest_6 = RTL_PATH.io_commits_info_1_debug_otherPdest_6; \
        force U_IF_NAME.io_commits_info_1_debug_fuType = RTL_PATH.io_commits_info_1_debug_fuType; \
        force U_IF_NAME.io_commits_info_1_dirtyFs = RTL_PATH.io_commits_info_1_dirtyFs; \
        force U_IF_NAME.io_commits_info_1_dirtyVs = RTL_PATH.io_commits_info_1_dirtyVs; \
        force U_IF_NAME.io_commits_info_2_walk_v = RTL_PATH.io_commits_info_2_walk_v; \
        force U_IF_NAME.io_commits_info_2_commit_v = RTL_PATH.io_commits_info_2_commit_v; \
        force U_IF_NAME.io_commits_info_2_commit_w = RTL_PATH.io_commits_info_2_commit_w; \
        force U_IF_NAME.io_commits_info_2_realDestSize = RTL_PATH.io_commits_info_2_realDestSize; \
        force U_IF_NAME.io_commits_info_2_interrupt_safe = RTL_PATH.io_commits_info_2_interrupt_safe; \
        force U_IF_NAME.io_commits_info_2_wflags = RTL_PATH.io_commits_info_2_wflags; \
        force U_IF_NAME.io_commits_info_2_fflags = RTL_PATH.io_commits_info_2_fflags; \
        force U_IF_NAME.io_commits_info_2_vxsat = RTL_PATH.io_commits_info_2_vxsat; \
        force U_IF_NAME.io_commits_info_2_isRVC = RTL_PATH.io_commits_info_2_isRVC; \
        force U_IF_NAME.io_commits_info_2_isVset = RTL_PATH.io_commits_info_2_isVset; \
        force U_IF_NAME.io_commits_info_2_isHls = RTL_PATH.io_commits_info_2_isHls; \
        force U_IF_NAME.io_commits_info_2_isVls = RTL_PATH.io_commits_info_2_isVls; \
        force U_IF_NAME.io_commits_info_2_vls = RTL_PATH.io_commits_info_2_vls; \
        force U_IF_NAME.io_commits_info_2_mmio = RTL_PATH.io_commits_info_2_mmio; \
        force U_IF_NAME.io_commits_info_2_commitType = RTL_PATH.io_commits_info_2_commitType; \
        force U_IF_NAME.io_commits_info_2_ftqIdx_flag = RTL_PATH.io_commits_info_2_ftqIdx_flag; \
        force U_IF_NAME.io_commits_info_2_ftqIdx_value = RTL_PATH.io_commits_info_2_ftqIdx_value; \
        force U_IF_NAME.io_commits_info_2_ftqOffset = RTL_PATH.io_commits_info_2_ftqOffset; \
        force U_IF_NAME.io_commits_info_2_instrSize = RTL_PATH.io_commits_info_2_instrSize; \
        force U_IF_NAME.io_commits_info_2_fpWen = RTL_PATH.io_commits_info_2_fpWen; \
        force U_IF_NAME.io_commits_info_2_rfWen = RTL_PATH.io_commits_info_2_rfWen; \
        force U_IF_NAME.io_commits_info_2_needFlush = RTL_PATH.io_commits_info_2_needFlush; \
        force U_IF_NAME.io_commits_info_2_traceBlockInPipe_itype = RTL_PATH.io_commits_info_2_traceBlockInPipe_itype; \
        force U_IF_NAME.io_commits_info_2_traceBlockInPipe_iretire = RTL_PATH.io_commits_info_2_traceBlockInPipe_iretire; \
        force U_IF_NAME.io_commits_info_2_traceBlockInPipe_ilastsize = RTL_PATH.io_commits_info_2_traceBlockInPipe_ilastsize; \
        force U_IF_NAME.io_commits_info_2_debug_pc = RTL_PATH.io_commits_info_2_debug_pc; \
        force U_IF_NAME.io_commits_info_2_debug_instr = RTL_PATH.io_commits_info_2_debug_instr; \
        force U_IF_NAME.io_commits_info_2_debug_ldest = RTL_PATH.io_commits_info_2_debug_ldest; \
        force U_IF_NAME.io_commits_info_2_debug_pdest = RTL_PATH.io_commits_info_2_debug_pdest; \
        force U_IF_NAME.io_commits_info_2_debug_otherPdest_0 = RTL_PATH.io_commits_info_2_debug_otherPdest_0; \
        force U_IF_NAME.io_commits_info_2_debug_otherPdest_1 = RTL_PATH.io_commits_info_2_debug_otherPdest_1; \
        force U_IF_NAME.io_commits_info_2_debug_otherPdest_2 = RTL_PATH.io_commits_info_2_debug_otherPdest_2; \
        force U_IF_NAME.io_commits_info_2_debug_otherPdest_3 = RTL_PATH.io_commits_info_2_debug_otherPdest_3; \
        force U_IF_NAME.io_commits_info_2_debug_otherPdest_4 = RTL_PATH.io_commits_info_2_debug_otherPdest_4; \
        force U_IF_NAME.io_commits_info_2_debug_otherPdest_5 = RTL_PATH.io_commits_info_2_debug_otherPdest_5; \
        force U_IF_NAME.io_commits_info_2_debug_otherPdest_6 = RTL_PATH.io_commits_info_2_debug_otherPdest_6; \
        force U_IF_NAME.io_commits_info_2_debug_fuType = RTL_PATH.io_commits_info_2_debug_fuType; \
        force U_IF_NAME.io_commits_info_2_dirtyFs = RTL_PATH.io_commits_info_2_dirtyFs; \
        force U_IF_NAME.io_commits_info_2_dirtyVs = RTL_PATH.io_commits_info_2_dirtyVs; \
        force U_IF_NAME.io_commits_info_3_walk_v = RTL_PATH.io_commits_info_3_walk_v; \
        force U_IF_NAME.io_commits_info_3_commit_v = RTL_PATH.io_commits_info_3_commit_v; \
        force U_IF_NAME.io_commits_info_3_commit_w = RTL_PATH.io_commits_info_3_commit_w; \
        force U_IF_NAME.io_commits_info_3_realDestSize = RTL_PATH.io_commits_info_3_realDestSize; \
        force U_IF_NAME.io_commits_info_3_interrupt_safe = RTL_PATH.io_commits_info_3_interrupt_safe; \
        force U_IF_NAME.io_commits_info_3_wflags = RTL_PATH.io_commits_info_3_wflags; \
        force U_IF_NAME.io_commits_info_3_fflags = RTL_PATH.io_commits_info_3_fflags; \
        force U_IF_NAME.io_commits_info_3_vxsat = RTL_PATH.io_commits_info_3_vxsat; \
        force U_IF_NAME.io_commits_info_3_isRVC = RTL_PATH.io_commits_info_3_isRVC; \
        force U_IF_NAME.io_commits_info_3_isVset = RTL_PATH.io_commits_info_3_isVset; \
        force U_IF_NAME.io_commits_info_3_isHls = RTL_PATH.io_commits_info_3_isHls; \
        force U_IF_NAME.io_commits_info_3_isVls = RTL_PATH.io_commits_info_3_isVls; \
        force U_IF_NAME.io_commits_info_3_vls = RTL_PATH.io_commits_info_3_vls; \
        force U_IF_NAME.io_commits_info_3_mmio = RTL_PATH.io_commits_info_3_mmio; \
        force U_IF_NAME.io_commits_info_3_commitType = RTL_PATH.io_commits_info_3_commitType; \
        force U_IF_NAME.io_commits_info_3_ftqIdx_flag = RTL_PATH.io_commits_info_3_ftqIdx_flag; \
        force U_IF_NAME.io_commits_info_3_ftqIdx_value = RTL_PATH.io_commits_info_3_ftqIdx_value; \
        force U_IF_NAME.io_commits_info_3_ftqOffset = RTL_PATH.io_commits_info_3_ftqOffset; \
        force U_IF_NAME.io_commits_info_3_instrSize = RTL_PATH.io_commits_info_3_instrSize; \
        force U_IF_NAME.io_commits_info_3_fpWen = RTL_PATH.io_commits_info_3_fpWen; \
        force U_IF_NAME.io_commits_info_3_rfWen = RTL_PATH.io_commits_info_3_rfWen; \
        force U_IF_NAME.io_commits_info_3_needFlush = RTL_PATH.io_commits_info_3_needFlush; \
        force U_IF_NAME.io_commits_info_3_traceBlockInPipe_itype = RTL_PATH.io_commits_info_3_traceBlockInPipe_itype; \
        force U_IF_NAME.io_commits_info_3_traceBlockInPipe_iretire = RTL_PATH.io_commits_info_3_traceBlockInPipe_iretire; \
        force U_IF_NAME.io_commits_info_3_traceBlockInPipe_ilastsize = RTL_PATH.io_commits_info_3_traceBlockInPipe_ilastsize; \
        force U_IF_NAME.io_commits_info_3_debug_pc = RTL_PATH.io_commits_info_3_debug_pc; \
        force U_IF_NAME.io_commits_info_3_debug_instr = RTL_PATH.io_commits_info_3_debug_instr; \
        force U_IF_NAME.io_commits_info_3_debug_ldest = RTL_PATH.io_commits_info_3_debug_ldest; \
        force U_IF_NAME.io_commits_info_3_debug_pdest = RTL_PATH.io_commits_info_3_debug_pdest; \
        force U_IF_NAME.io_commits_info_3_debug_otherPdest_0 = RTL_PATH.io_commits_info_3_debug_otherPdest_0; \
        force U_IF_NAME.io_commits_info_3_debug_otherPdest_1 = RTL_PATH.io_commits_info_3_debug_otherPdest_1; \
        force U_IF_NAME.io_commits_info_3_debug_otherPdest_2 = RTL_PATH.io_commits_info_3_debug_otherPdest_2; \
        force U_IF_NAME.io_commits_info_3_debug_otherPdest_3 = RTL_PATH.io_commits_info_3_debug_otherPdest_3; \
        force U_IF_NAME.io_commits_info_3_debug_otherPdest_4 = RTL_PATH.io_commits_info_3_debug_otherPdest_4; \
        force U_IF_NAME.io_commits_info_3_debug_otherPdest_5 = RTL_PATH.io_commits_info_3_debug_otherPdest_5; \
        force U_IF_NAME.io_commits_info_3_debug_otherPdest_6 = RTL_PATH.io_commits_info_3_debug_otherPdest_6; \
        force U_IF_NAME.io_commits_info_3_debug_fuType = RTL_PATH.io_commits_info_3_debug_fuType; \
        force U_IF_NAME.io_commits_info_3_dirtyFs = RTL_PATH.io_commits_info_3_dirtyFs; \
        force U_IF_NAME.io_commits_info_3_dirtyVs = RTL_PATH.io_commits_info_3_dirtyVs; \
        force U_IF_NAME.io_commits_info_4_walk_v = RTL_PATH.io_commits_info_4_walk_v; \
        force U_IF_NAME.io_commits_info_4_commit_v = RTL_PATH.io_commits_info_4_commit_v; \
        force U_IF_NAME.io_commits_info_4_commit_w = RTL_PATH.io_commits_info_4_commit_w; \
        force U_IF_NAME.io_commits_info_4_realDestSize = RTL_PATH.io_commits_info_4_realDestSize; \
        force U_IF_NAME.io_commits_info_4_interrupt_safe = RTL_PATH.io_commits_info_4_interrupt_safe; \
        force U_IF_NAME.io_commits_info_4_wflags = RTL_PATH.io_commits_info_4_wflags; \
        force U_IF_NAME.io_commits_info_4_fflags = RTL_PATH.io_commits_info_4_fflags; \
        force U_IF_NAME.io_commits_info_4_vxsat = RTL_PATH.io_commits_info_4_vxsat; \
        force U_IF_NAME.io_commits_info_4_isRVC = RTL_PATH.io_commits_info_4_isRVC; \
        force U_IF_NAME.io_commits_info_4_isVset = RTL_PATH.io_commits_info_4_isVset; \
        force U_IF_NAME.io_commits_info_4_isHls = RTL_PATH.io_commits_info_4_isHls; \
        force U_IF_NAME.io_commits_info_4_isVls = RTL_PATH.io_commits_info_4_isVls; \
        force U_IF_NAME.io_commits_info_4_vls = RTL_PATH.io_commits_info_4_vls; \
        force U_IF_NAME.io_commits_info_4_mmio = RTL_PATH.io_commits_info_4_mmio; \
        force U_IF_NAME.io_commits_info_4_commitType = RTL_PATH.io_commits_info_4_commitType; \
        force U_IF_NAME.io_commits_info_4_ftqIdx_flag = RTL_PATH.io_commits_info_4_ftqIdx_flag; \
        force U_IF_NAME.io_commits_info_4_ftqIdx_value = RTL_PATH.io_commits_info_4_ftqIdx_value; \
        force U_IF_NAME.io_commits_info_4_ftqOffset = RTL_PATH.io_commits_info_4_ftqOffset; \
        force U_IF_NAME.io_commits_info_4_instrSize = RTL_PATH.io_commits_info_4_instrSize; \
        force U_IF_NAME.io_commits_info_4_fpWen = RTL_PATH.io_commits_info_4_fpWen; \
        force U_IF_NAME.io_commits_info_4_rfWen = RTL_PATH.io_commits_info_4_rfWen; \
        force U_IF_NAME.io_commits_info_4_needFlush = RTL_PATH.io_commits_info_4_needFlush; \
        force U_IF_NAME.io_commits_info_4_traceBlockInPipe_itype = RTL_PATH.io_commits_info_4_traceBlockInPipe_itype; \
        force U_IF_NAME.io_commits_info_4_traceBlockInPipe_iretire = RTL_PATH.io_commits_info_4_traceBlockInPipe_iretire; \
        force U_IF_NAME.io_commits_info_4_traceBlockInPipe_ilastsize = RTL_PATH.io_commits_info_4_traceBlockInPipe_ilastsize; \
        force U_IF_NAME.io_commits_info_4_debug_pc = RTL_PATH.io_commits_info_4_debug_pc; \
        force U_IF_NAME.io_commits_info_4_debug_instr = RTL_PATH.io_commits_info_4_debug_instr; \
        force U_IF_NAME.io_commits_info_4_debug_ldest = RTL_PATH.io_commits_info_4_debug_ldest; \
        force U_IF_NAME.io_commits_info_4_debug_pdest = RTL_PATH.io_commits_info_4_debug_pdest; \
        force U_IF_NAME.io_commits_info_4_debug_otherPdest_0 = RTL_PATH.io_commits_info_4_debug_otherPdest_0; \
        force U_IF_NAME.io_commits_info_4_debug_otherPdest_1 = RTL_PATH.io_commits_info_4_debug_otherPdest_1; \
        force U_IF_NAME.io_commits_info_4_debug_otherPdest_2 = RTL_PATH.io_commits_info_4_debug_otherPdest_2; \
        force U_IF_NAME.io_commits_info_4_debug_otherPdest_3 = RTL_PATH.io_commits_info_4_debug_otherPdest_3; \
        force U_IF_NAME.io_commits_info_4_debug_otherPdest_4 = RTL_PATH.io_commits_info_4_debug_otherPdest_4; \
        force U_IF_NAME.io_commits_info_4_debug_otherPdest_5 = RTL_PATH.io_commits_info_4_debug_otherPdest_5; \
        force U_IF_NAME.io_commits_info_4_debug_otherPdest_6 = RTL_PATH.io_commits_info_4_debug_otherPdest_6; \
        force U_IF_NAME.io_commits_info_4_debug_fuType = RTL_PATH.io_commits_info_4_debug_fuType; \
        force U_IF_NAME.io_commits_info_4_dirtyFs = RTL_PATH.io_commits_info_4_dirtyFs; \
        force U_IF_NAME.io_commits_info_4_dirtyVs = RTL_PATH.io_commits_info_4_dirtyVs; \
        force U_IF_NAME.io_commits_info_5_walk_v = RTL_PATH.io_commits_info_5_walk_v; \
        force U_IF_NAME.io_commits_info_5_commit_v = RTL_PATH.io_commits_info_5_commit_v; \
        force U_IF_NAME.io_commits_info_5_commit_w = RTL_PATH.io_commits_info_5_commit_w; \
        force U_IF_NAME.io_commits_info_5_realDestSize = RTL_PATH.io_commits_info_5_realDestSize; \
        force U_IF_NAME.io_commits_info_5_interrupt_safe = RTL_PATH.io_commits_info_5_interrupt_safe; \
        force U_IF_NAME.io_commits_info_5_wflags = RTL_PATH.io_commits_info_5_wflags; \
        force U_IF_NAME.io_commits_info_5_fflags = RTL_PATH.io_commits_info_5_fflags; \
        force U_IF_NAME.io_commits_info_5_vxsat = RTL_PATH.io_commits_info_5_vxsat; \
        force U_IF_NAME.io_commits_info_5_isRVC = RTL_PATH.io_commits_info_5_isRVC; \
        force U_IF_NAME.io_commits_info_5_isVset = RTL_PATH.io_commits_info_5_isVset; \
        force U_IF_NAME.io_commits_info_5_isHls = RTL_PATH.io_commits_info_5_isHls; \
        force U_IF_NAME.io_commits_info_5_isVls = RTL_PATH.io_commits_info_5_isVls; \
        force U_IF_NAME.io_commits_info_5_vls = RTL_PATH.io_commits_info_5_vls; \
        force U_IF_NAME.io_commits_info_5_mmio = RTL_PATH.io_commits_info_5_mmio; \
        force U_IF_NAME.io_commits_info_5_commitType = RTL_PATH.io_commits_info_5_commitType; \
        force U_IF_NAME.io_commits_info_5_ftqIdx_flag = RTL_PATH.io_commits_info_5_ftqIdx_flag; \
        force U_IF_NAME.io_commits_info_5_ftqIdx_value = RTL_PATH.io_commits_info_5_ftqIdx_value; \
        force U_IF_NAME.io_commits_info_5_ftqOffset = RTL_PATH.io_commits_info_5_ftqOffset; \
        force U_IF_NAME.io_commits_info_5_instrSize = RTL_PATH.io_commits_info_5_instrSize; \
        force U_IF_NAME.io_commits_info_5_fpWen = RTL_PATH.io_commits_info_5_fpWen; \
        force U_IF_NAME.io_commits_info_5_rfWen = RTL_PATH.io_commits_info_5_rfWen; \
        force U_IF_NAME.io_commits_info_5_needFlush = RTL_PATH.io_commits_info_5_needFlush; \
        force U_IF_NAME.io_commits_info_5_traceBlockInPipe_itype = RTL_PATH.io_commits_info_5_traceBlockInPipe_itype; \
        force U_IF_NAME.io_commits_info_5_traceBlockInPipe_iretire = RTL_PATH.io_commits_info_5_traceBlockInPipe_iretire; \
        force U_IF_NAME.io_commits_info_5_traceBlockInPipe_ilastsize = RTL_PATH.io_commits_info_5_traceBlockInPipe_ilastsize; \
        force U_IF_NAME.io_commits_info_5_debug_pc = RTL_PATH.io_commits_info_5_debug_pc; \
        force U_IF_NAME.io_commits_info_5_debug_instr = RTL_PATH.io_commits_info_5_debug_instr; \
        force U_IF_NAME.io_commits_info_5_debug_ldest = RTL_PATH.io_commits_info_5_debug_ldest; \
        force U_IF_NAME.io_commits_info_5_debug_pdest = RTL_PATH.io_commits_info_5_debug_pdest; \
        force U_IF_NAME.io_commits_info_5_debug_otherPdest_0 = RTL_PATH.io_commits_info_5_debug_otherPdest_0; \
        force U_IF_NAME.io_commits_info_5_debug_otherPdest_1 = RTL_PATH.io_commits_info_5_debug_otherPdest_1; \
        force U_IF_NAME.io_commits_info_5_debug_otherPdest_2 = RTL_PATH.io_commits_info_5_debug_otherPdest_2; \
        force U_IF_NAME.io_commits_info_5_debug_otherPdest_3 = RTL_PATH.io_commits_info_5_debug_otherPdest_3; \
        force U_IF_NAME.io_commits_info_5_debug_otherPdest_4 = RTL_PATH.io_commits_info_5_debug_otherPdest_4; \
        force U_IF_NAME.io_commits_info_5_debug_otherPdest_5 = RTL_PATH.io_commits_info_5_debug_otherPdest_5; \
        force U_IF_NAME.io_commits_info_5_debug_otherPdest_6 = RTL_PATH.io_commits_info_5_debug_otherPdest_6; \
        force U_IF_NAME.io_commits_info_5_debug_fuType = RTL_PATH.io_commits_info_5_debug_fuType; \
        force U_IF_NAME.io_commits_info_5_dirtyFs = RTL_PATH.io_commits_info_5_dirtyFs; \
        force U_IF_NAME.io_commits_info_5_dirtyVs = RTL_PATH.io_commits_info_5_dirtyVs; \
        force U_IF_NAME.io_commits_info_6_walk_v = RTL_PATH.io_commits_info_6_walk_v; \
        force U_IF_NAME.io_commits_info_6_commit_v = RTL_PATH.io_commits_info_6_commit_v; \
        force U_IF_NAME.io_commits_info_6_commit_w = RTL_PATH.io_commits_info_6_commit_w; \
        force U_IF_NAME.io_commits_info_6_realDestSize = RTL_PATH.io_commits_info_6_realDestSize; \
        force U_IF_NAME.io_commits_info_6_interrupt_safe = RTL_PATH.io_commits_info_6_interrupt_safe; \
        force U_IF_NAME.io_commits_info_6_wflags = RTL_PATH.io_commits_info_6_wflags; \
        force U_IF_NAME.io_commits_info_6_fflags = RTL_PATH.io_commits_info_6_fflags; \
        force U_IF_NAME.io_commits_info_6_vxsat = RTL_PATH.io_commits_info_6_vxsat; \
        force U_IF_NAME.io_commits_info_6_isRVC = RTL_PATH.io_commits_info_6_isRVC; \
        force U_IF_NAME.io_commits_info_6_isVset = RTL_PATH.io_commits_info_6_isVset; \
        force U_IF_NAME.io_commits_info_6_isHls = RTL_PATH.io_commits_info_6_isHls; \
        force U_IF_NAME.io_commits_info_6_isVls = RTL_PATH.io_commits_info_6_isVls; \
        force U_IF_NAME.io_commits_info_6_vls = RTL_PATH.io_commits_info_6_vls; \
        force U_IF_NAME.io_commits_info_6_mmio = RTL_PATH.io_commits_info_6_mmio; \
        force U_IF_NAME.io_commits_info_6_commitType = RTL_PATH.io_commits_info_6_commitType; \
        force U_IF_NAME.io_commits_info_6_ftqIdx_flag = RTL_PATH.io_commits_info_6_ftqIdx_flag; \
        force U_IF_NAME.io_commits_info_6_ftqIdx_value = RTL_PATH.io_commits_info_6_ftqIdx_value; \
        force U_IF_NAME.io_commits_info_6_ftqOffset = RTL_PATH.io_commits_info_6_ftqOffset; \
        force U_IF_NAME.io_commits_info_6_instrSize = RTL_PATH.io_commits_info_6_instrSize; \
        force U_IF_NAME.io_commits_info_6_fpWen = RTL_PATH.io_commits_info_6_fpWen; \
        force U_IF_NAME.io_commits_info_6_rfWen = RTL_PATH.io_commits_info_6_rfWen; \
        force U_IF_NAME.io_commits_info_6_needFlush = RTL_PATH.io_commits_info_6_needFlush; \
        force U_IF_NAME.io_commits_info_6_traceBlockInPipe_itype = RTL_PATH.io_commits_info_6_traceBlockInPipe_itype; \
        force U_IF_NAME.io_commits_info_6_traceBlockInPipe_iretire = RTL_PATH.io_commits_info_6_traceBlockInPipe_iretire; \
        force U_IF_NAME.io_commits_info_6_traceBlockInPipe_ilastsize = RTL_PATH.io_commits_info_6_traceBlockInPipe_ilastsize; \
        force U_IF_NAME.io_commits_info_6_debug_pc = RTL_PATH.io_commits_info_6_debug_pc; \
        force U_IF_NAME.io_commits_info_6_debug_instr = RTL_PATH.io_commits_info_6_debug_instr; \
        force U_IF_NAME.io_commits_info_6_debug_ldest = RTL_PATH.io_commits_info_6_debug_ldest; \
        force U_IF_NAME.io_commits_info_6_debug_pdest = RTL_PATH.io_commits_info_6_debug_pdest; \
        force U_IF_NAME.io_commits_info_6_debug_otherPdest_0 = RTL_PATH.io_commits_info_6_debug_otherPdest_0; \
        force U_IF_NAME.io_commits_info_6_debug_otherPdest_1 = RTL_PATH.io_commits_info_6_debug_otherPdest_1; \
        force U_IF_NAME.io_commits_info_6_debug_otherPdest_2 = RTL_PATH.io_commits_info_6_debug_otherPdest_2; \
        force U_IF_NAME.io_commits_info_6_debug_otherPdest_3 = RTL_PATH.io_commits_info_6_debug_otherPdest_3; \
        force U_IF_NAME.io_commits_info_6_debug_otherPdest_4 = RTL_PATH.io_commits_info_6_debug_otherPdest_4; \
        force U_IF_NAME.io_commits_info_6_debug_otherPdest_5 = RTL_PATH.io_commits_info_6_debug_otherPdest_5; \
        force U_IF_NAME.io_commits_info_6_debug_otherPdest_6 = RTL_PATH.io_commits_info_6_debug_otherPdest_6; \
        force U_IF_NAME.io_commits_info_6_debug_fuType = RTL_PATH.io_commits_info_6_debug_fuType; \
        force U_IF_NAME.io_commits_info_6_dirtyFs = RTL_PATH.io_commits_info_6_dirtyFs; \
        force U_IF_NAME.io_commits_info_6_dirtyVs = RTL_PATH.io_commits_info_6_dirtyVs; \
        force U_IF_NAME.io_commits_info_7_walk_v = RTL_PATH.io_commits_info_7_walk_v; \
        force U_IF_NAME.io_commits_info_7_commit_v = RTL_PATH.io_commits_info_7_commit_v; \
        force U_IF_NAME.io_commits_info_7_commit_w = RTL_PATH.io_commits_info_7_commit_w; \
        force U_IF_NAME.io_commits_info_7_realDestSize = RTL_PATH.io_commits_info_7_realDestSize; \
        force U_IF_NAME.io_commits_info_7_interrupt_safe = RTL_PATH.io_commits_info_7_interrupt_safe; \
        force U_IF_NAME.io_commits_info_7_wflags = RTL_PATH.io_commits_info_7_wflags; \
        force U_IF_NAME.io_commits_info_7_fflags = RTL_PATH.io_commits_info_7_fflags; \
        force U_IF_NAME.io_commits_info_7_vxsat = RTL_PATH.io_commits_info_7_vxsat; \
        force U_IF_NAME.io_commits_info_7_isRVC = RTL_PATH.io_commits_info_7_isRVC; \
        force U_IF_NAME.io_commits_info_7_isVset = RTL_PATH.io_commits_info_7_isVset; \
        force U_IF_NAME.io_commits_info_7_isHls = RTL_PATH.io_commits_info_7_isHls; \
        force U_IF_NAME.io_commits_info_7_isVls = RTL_PATH.io_commits_info_7_isVls; \
        force U_IF_NAME.io_commits_info_7_vls = RTL_PATH.io_commits_info_7_vls; \
        force U_IF_NAME.io_commits_info_7_mmio = RTL_PATH.io_commits_info_7_mmio; \
        force U_IF_NAME.io_commits_info_7_commitType = RTL_PATH.io_commits_info_7_commitType; \
        force U_IF_NAME.io_commits_info_7_ftqIdx_flag = RTL_PATH.io_commits_info_7_ftqIdx_flag; \
        force U_IF_NAME.io_commits_info_7_ftqIdx_value = RTL_PATH.io_commits_info_7_ftqIdx_value; \
        force U_IF_NAME.io_commits_info_7_ftqOffset = RTL_PATH.io_commits_info_7_ftqOffset; \
        force U_IF_NAME.io_commits_info_7_instrSize = RTL_PATH.io_commits_info_7_instrSize; \
        force U_IF_NAME.io_commits_info_7_fpWen = RTL_PATH.io_commits_info_7_fpWen; \
        force U_IF_NAME.io_commits_info_7_rfWen = RTL_PATH.io_commits_info_7_rfWen; \
        force U_IF_NAME.io_commits_info_7_needFlush = RTL_PATH.io_commits_info_7_needFlush; \
        force U_IF_NAME.io_commits_info_7_traceBlockInPipe_itype = RTL_PATH.io_commits_info_7_traceBlockInPipe_itype; \
        force U_IF_NAME.io_commits_info_7_traceBlockInPipe_iretire = RTL_PATH.io_commits_info_7_traceBlockInPipe_iretire; \
        force U_IF_NAME.io_commits_info_7_traceBlockInPipe_ilastsize = RTL_PATH.io_commits_info_7_traceBlockInPipe_ilastsize; \
        force U_IF_NAME.io_commits_info_7_debug_pc = RTL_PATH.io_commits_info_7_debug_pc; \
        force U_IF_NAME.io_commits_info_7_debug_instr = RTL_PATH.io_commits_info_7_debug_instr; \
        force U_IF_NAME.io_commits_info_7_debug_ldest = RTL_PATH.io_commits_info_7_debug_ldest; \
        force U_IF_NAME.io_commits_info_7_debug_pdest = RTL_PATH.io_commits_info_7_debug_pdest; \
        force U_IF_NAME.io_commits_info_7_debug_otherPdest_0 = RTL_PATH.io_commits_info_7_debug_otherPdest_0; \
        force U_IF_NAME.io_commits_info_7_debug_otherPdest_1 = RTL_PATH.io_commits_info_7_debug_otherPdest_1; \
        force U_IF_NAME.io_commits_info_7_debug_otherPdest_2 = RTL_PATH.io_commits_info_7_debug_otherPdest_2; \
        force U_IF_NAME.io_commits_info_7_debug_otherPdest_3 = RTL_PATH.io_commits_info_7_debug_otherPdest_3; \
        force U_IF_NAME.io_commits_info_7_debug_otherPdest_4 = RTL_PATH.io_commits_info_7_debug_otherPdest_4; \
        force U_IF_NAME.io_commits_info_7_debug_otherPdest_5 = RTL_PATH.io_commits_info_7_debug_otherPdest_5; \
        force U_IF_NAME.io_commits_info_7_debug_otherPdest_6 = RTL_PATH.io_commits_info_7_debug_otherPdest_6; \
        force U_IF_NAME.io_commits_info_7_debug_fuType = RTL_PATH.io_commits_info_7_debug_fuType; \
        force U_IF_NAME.io_commits_info_7_dirtyFs = RTL_PATH.io_commits_info_7_dirtyFs; \
        force U_IF_NAME.io_commits_info_7_dirtyVs = RTL_PATH.io_commits_info_7_dirtyVs; \
        force U_IF_NAME.io_commits_robIdx_0_flag = RTL_PATH.io_commits_robIdx_0_flag; \
        force U_IF_NAME.io_commits_robIdx_0_value = RTL_PATH.io_commits_robIdx_0_value; \
        force U_IF_NAME.io_commits_robIdx_1_flag = RTL_PATH.io_commits_robIdx_1_flag; \
        force U_IF_NAME.io_commits_robIdx_1_value = RTL_PATH.io_commits_robIdx_1_value; \
        force U_IF_NAME.io_commits_robIdx_2_flag = RTL_PATH.io_commits_robIdx_2_flag; \
        force U_IF_NAME.io_commits_robIdx_2_value = RTL_PATH.io_commits_robIdx_2_value; \
        force U_IF_NAME.io_commits_robIdx_3_flag = RTL_PATH.io_commits_robIdx_3_flag; \
        force U_IF_NAME.io_commits_robIdx_3_value = RTL_PATH.io_commits_robIdx_3_value; \
        force U_IF_NAME.io_commits_robIdx_4_flag = RTL_PATH.io_commits_robIdx_4_flag; \
        force U_IF_NAME.io_commits_robIdx_4_value = RTL_PATH.io_commits_robIdx_4_value; \
        force U_IF_NAME.io_commits_robIdx_5_flag = RTL_PATH.io_commits_robIdx_5_flag; \
        force U_IF_NAME.io_commits_robIdx_5_value = RTL_PATH.io_commits_robIdx_5_value; \
        force U_IF_NAME.io_commits_robIdx_6_flag = RTL_PATH.io_commits_robIdx_6_flag; \
        force U_IF_NAME.io_commits_robIdx_6_value = RTL_PATH.io_commits_robIdx_6_value; \
        force U_IF_NAME.io_commits_robIdx_7_flag = RTL_PATH.io_commits_robIdx_7_flag; \
        force U_IF_NAME.io_commits_robIdx_7_value = RTL_PATH.io_commits_robIdx_7_value; \
        force U_IF_NAME.io_trace_blockCommit = RTL_PATH.io_trace_blockCommit; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_0_valid = RTL_PATH.io_trace_traceCommitInfo_blocks_0_valid; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value = RTL_PATH.io_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_0_bits_ftqOffset = RTL_PATH.io_trace_traceCommitInfo_blocks_0_bits_ftqOffset; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype = RTL_PATH.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire = RTL_PATH.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize = RTL_PATH.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_1_valid = RTL_PATH.io_trace_traceCommitInfo_blocks_1_valid; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value = RTL_PATH.io_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_1_bits_ftqOffset = RTL_PATH.io_trace_traceCommitInfo_blocks_1_bits_ftqOffset; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype = RTL_PATH.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire = RTL_PATH.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize = RTL_PATH.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_2_valid = RTL_PATH.io_trace_traceCommitInfo_blocks_2_valid; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value = RTL_PATH.io_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_2_bits_ftqOffset = RTL_PATH.io_trace_traceCommitInfo_blocks_2_bits_ftqOffset; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype = RTL_PATH.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire = RTL_PATH.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize = RTL_PATH.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_3_valid = RTL_PATH.io_trace_traceCommitInfo_blocks_3_valid; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value = RTL_PATH.io_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_3_bits_ftqOffset = RTL_PATH.io_trace_traceCommitInfo_blocks_3_bits_ftqOffset; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype = RTL_PATH.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire = RTL_PATH.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize = RTL_PATH.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_4_valid = RTL_PATH.io_trace_traceCommitInfo_blocks_4_valid; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value = RTL_PATH.io_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_4_bits_ftqOffset = RTL_PATH.io_trace_traceCommitInfo_blocks_4_bits_ftqOffset; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype = RTL_PATH.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire = RTL_PATH.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize = RTL_PATH.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_5_valid = RTL_PATH.io_trace_traceCommitInfo_blocks_5_valid; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value = RTL_PATH.io_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_5_bits_ftqOffset = RTL_PATH.io_trace_traceCommitInfo_blocks_5_bits_ftqOffset; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype = RTL_PATH.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire = RTL_PATH.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize = RTL_PATH.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_6_valid = RTL_PATH.io_trace_traceCommitInfo_blocks_6_valid; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value = RTL_PATH.io_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_6_bits_ftqOffset = RTL_PATH.io_trace_traceCommitInfo_blocks_6_bits_ftqOffset; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype = RTL_PATH.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire = RTL_PATH.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize = RTL_PATH.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_7_valid = RTL_PATH.io_trace_traceCommitInfo_blocks_7_valid; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value = RTL_PATH.io_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_7_bits_ftqOffset = RTL_PATH.io_trace_traceCommitInfo_blocks_7_bits_ftqOffset; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype = RTL_PATH.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire = RTL_PATH.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire; \
        force U_IF_NAME.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize = RTL_PATH.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize; \
        force U_IF_NAME.io_rabCommits_isCommit = RTL_PATH.io_rabCommits_isCommit; \
        force U_IF_NAME.io_rabCommits_commitValid_0 = RTL_PATH.io_rabCommits_commitValid_0; \
        force U_IF_NAME.io_rabCommits_commitValid_1 = RTL_PATH.io_rabCommits_commitValid_1; \
        force U_IF_NAME.io_rabCommits_commitValid_2 = RTL_PATH.io_rabCommits_commitValid_2; \
        force U_IF_NAME.io_rabCommits_commitValid_3 = RTL_PATH.io_rabCommits_commitValid_3; \
        force U_IF_NAME.io_rabCommits_commitValid_4 = RTL_PATH.io_rabCommits_commitValid_4; \
        force U_IF_NAME.io_rabCommits_commitValid_5 = RTL_PATH.io_rabCommits_commitValid_5; \
        force U_IF_NAME.io_rabCommits_isWalk = RTL_PATH.io_rabCommits_isWalk; \
        force U_IF_NAME.io_rabCommits_walkValid_0 = RTL_PATH.io_rabCommits_walkValid_0; \
        force U_IF_NAME.io_rabCommits_walkValid_1 = RTL_PATH.io_rabCommits_walkValid_1; \
        force U_IF_NAME.io_rabCommits_walkValid_2 = RTL_PATH.io_rabCommits_walkValid_2; \
        force U_IF_NAME.io_rabCommits_walkValid_3 = RTL_PATH.io_rabCommits_walkValid_3; \
        force U_IF_NAME.io_rabCommits_walkValid_4 = RTL_PATH.io_rabCommits_walkValid_4; \
        force U_IF_NAME.io_rabCommits_walkValid_5 = RTL_PATH.io_rabCommits_walkValid_5; \
        force U_IF_NAME.io_rabCommits_info_0_ldest = RTL_PATH.io_rabCommits_info_0_ldest; \
        force U_IF_NAME.io_rabCommits_info_0_pdest = RTL_PATH.io_rabCommits_info_0_pdest; \
        force U_IF_NAME.io_rabCommits_info_0_rfWen = RTL_PATH.io_rabCommits_info_0_rfWen; \
        force U_IF_NAME.io_rabCommits_info_0_fpWen = RTL_PATH.io_rabCommits_info_0_fpWen; \
        force U_IF_NAME.io_rabCommits_info_0_vecWen = RTL_PATH.io_rabCommits_info_0_vecWen; \
        force U_IF_NAME.io_rabCommits_info_0_v0Wen = RTL_PATH.io_rabCommits_info_0_v0Wen; \
        force U_IF_NAME.io_rabCommits_info_0_vlWen = RTL_PATH.io_rabCommits_info_0_vlWen; \
        force U_IF_NAME.io_rabCommits_info_0_isMove = RTL_PATH.io_rabCommits_info_0_isMove; \
        force U_IF_NAME.io_rabCommits_info_1_ldest = RTL_PATH.io_rabCommits_info_1_ldest; \
        force U_IF_NAME.io_rabCommits_info_1_pdest = RTL_PATH.io_rabCommits_info_1_pdest; \
        force U_IF_NAME.io_rabCommits_info_1_rfWen = RTL_PATH.io_rabCommits_info_1_rfWen; \
        force U_IF_NAME.io_rabCommits_info_1_fpWen = RTL_PATH.io_rabCommits_info_1_fpWen; \
        force U_IF_NAME.io_rabCommits_info_1_vecWen = RTL_PATH.io_rabCommits_info_1_vecWen; \
        force U_IF_NAME.io_rabCommits_info_1_v0Wen = RTL_PATH.io_rabCommits_info_1_v0Wen; \
        force U_IF_NAME.io_rabCommits_info_1_vlWen = RTL_PATH.io_rabCommits_info_1_vlWen; \
        force U_IF_NAME.io_rabCommits_info_1_isMove = RTL_PATH.io_rabCommits_info_1_isMove; \
        force U_IF_NAME.io_rabCommits_info_2_ldest = RTL_PATH.io_rabCommits_info_2_ldest; \
        force U_IF_NAME.io_rabCommits_info_2_pdest = RTL_PATH.io_rabCommits_info_2_pdest; \
        force U_IF_NAME.io_rabCommits_info_2_rfWen = RTL_PATH.io_rabCommits_info_2_rfWen; \
        force U_IF_NAME.io_rabCommits_info_2_fpWen = RTL_PATH.io_rabCommits_info_2_fpWen; \
        force U_IF_NAME.io_rabCommits_info_2_vecWen = RTL_PATH.io_rabCommits_info_2_vecWen; \
        force U_IF_NAME.io_rabCommits_info_2_v0Wen = RTL_PATH.io_rabCommits_info_2_v0Wen; \
        force U_IF_NAME.io_rabCommits_info_2_vlWen = RTL_PATH.io_rabCommits_info_2_vlWen; \
        force U_IF_NAME.io_rabCommits_info_2_isMove = RTL_PATH.io_rabCommits_info_2_isMove; \
        force U_IF_NAME.io_rabCommits_info_3_ldest = RTL_PATH.io_rabCommits_info_3_ldest; \
        force U_IF_NAME.io_rabCommits_info_3_pdest = RTL_PATH.io_rabCommits_info_3_pdest; \
        force U_IF_NAME.io_rabCommits_info_3_rfWen = RTL_PATH.io_rabCommits_info_3_rfWen; \
        force U_IF_NAME.io_rabCommits_info_3_fpWen = RTL_PATH.io_rabCommits_info_3_fpWen; \
        force U_IF_NAME.io_rabCommits_info_3_vecWen = RTL_PATH.io_rabCommits_info_3_vecWen; \
        force U_IF_NAME.io_rabCommits_info_3_v0Wen = RTL_PATH.io_rabCommits_info_3_v0Wen; \
        force U_IF_NAME.io_rabCommits_info_3_vlWen = RTL_PATH.io_rabCommits_info_3_vlWen; \
        force U_IF_NAME.io_rabCommits_info_3_isMove = RTL_PATH.io_rabCommits_info_3_isMove; \
        force U_IF_NAME.io_rabCommits_info_4_ldest = RTL_PATH.io_rabCommits_info_4_ldest; \
        force U_IF_NAME.io_rabCommits_info_4_pdest = RTL_PATH.io_rabCommits_info_4_pdest; \
        force U_IF_NAME.io_rabCommits_info_4_rfWen = RTL_PATH.io_rabCommits_info_4_rfWen; \
        force U_IF_NAME.io_rabCommits_info_4_fpWen = RTL_PATH.io_rabCommits_info_4_fpWen; \
        force U_IF_NAME.io_rabCommits_info_4_vecWen = RTL_PATH.io_rabCommits_info_4_vecWen; \
        force U_IF_NAME.io_rabCommits_info_4_v0Wen = RTL_PATH.io_rabCommits_info_4_v0Wen; \
        force U_IF_NAME.io_rabCommits_info_4_vlWen = RTL_PATH.io_rabCommits_info_4_vlWen; \
        force U_IF_NAME.io_rabCommits_info_4_isMove = RTL_PATH.io_rabCommits_info_4_isMove; \
        force U_IF_NAME.io_rabCommits_info_5_ldest = RTL_PATH.io_rabCommits_info_5_ldest; \
        force U_IF_NAME.io_rabCommits_info_5_pdest = RTL_PATH.io_rabCommits_info_5_pdest; \
        force U_IF_NAME.io_rabCommits_info_5_rfWen = RTL_PATH.io_rabCommits_info_5_rfWen; \
        force U_IF_NAME.io_rabCommits_info_5_fpWen = RTL_PATH.io_rabCommits_info_5_fpWen; \
        force U_IF_NAME.io_rabCommits_info_5_vecWen = RTL_PATH.io_rabCommits_info_5_vecWen; \
        force U_IF_NAME.io_rabCommits_info_5_v0Wen = RTL_PATH.io_rabCommits_info_5_v0Wen; \
        force U_IF_NAME.io_rabCommits_info_5_vlWen = RTL_PATH.io_rabCommits_info_5_vlWen; \
        force U_IF_NAME.io_rabCommits_info_5_isMove = RTL_PATH.io_rabCommits_info_5_isMove; \
        force U_IF_NAME.io_diffCommits_commitValid_0 = RTL_PATH.io_diffCommits_commitValid_0; \
        force U_IF_NAME.io_diffCommits_commitValid_1 = RTL_PATH.io_diffCommits_commitValid_1; \
        force U_IF_NAME.io_diffCommits_commitValid_2 = RTL_PATH.io_diffCommits_commitValid_2; \
        force U_IF_NAME.io_diffCommits_commitValid_3 = RTL_PATH.io_diffCommits_commitValid_3; \
        force U_IF_NAME.io_diffCommits_commitValid_4 = RTL_PATH.io_diffCommits_commitValid_4; \
        force U_IF_NAME.io_diffCommits_commitValid_5 = RTL_PATH.io_diffCommits_commitValid_5; \
        force U_IF_NAME.io_diffCommits_commitValid_6 = RTL_PATH.io_diffCommits_commitValid_6; \
        force U_IF_NAME.io_diffCommits_commitValid_7 = RTL_PATH.io_diffCommits_commitValid_7; \
        force U_IF_NAME.io_diffCommits_commitValid_8 = RTL_PATH.io_diffCommits_commitValid_8; \
        force U_IF_NAME.io_diffCommits_commitValid_9 = RTL_PATH.io_diffCommits_commitValid_9; \
        force U_IF_NAME.io_diffCommits_commitValid_10 = RTL_PATH.io_diffCommits_commitValid_10; \
        force U_IF_NAME.io_diffCommits_commitValid_11 = RTL_PATH.io_diffCommits_commitValid_11; \
        force U_IF_NAME.io_diffCommits_commitValid_12 = RTL_PATH.io_diffCommits_commitValid_12; \
        force U_IF_NAME.io_diffCommits_commitValid_13 = RTL_PATH.io_diffCommits_commitValid_13; \
        force U_IF_NAME.io_diffCommits_commitValid_14 = RTL_PATH.io_diffCommits_commitValid_14; \
        force U_IF_NAME.io_diffCommits_commitValid_15 = RTL_PATH.io_diffCommits_commitValid_15; \
        force U_IF_NAME.io_diffCommits_commitValid_16 = RTL_PATH.io_diffCommits_commitValid_16; \
        force U_IF_NAME.io_diffCommits_commitValid_17 = RTL_PATH.io_diffCommits_commitValid_17; \
        force U_IF_NAME.io_diffCommits_commitValid_18 = RTL_PATH.io_diffCommits_commitValid_18; \
        force U_IF_NAME.io_diffCommits_commitValid_19 = RTL_PATH.io_diffCommits_commitValid_19; \
        force U_IF_NAME.io_diffCommits_commitValid_20 = RTL_PATH.io_diffCommits_commitValid_20; \
        force U_IF_NAME.io_diffCommits_commitValid_21 = RTL_PATH.io_diffCommits_commitValid_21; \
        force U_IF_NAME.io_diffCommits_commitValid_22 = RTL_PATH.io_diffCommits_commitValid_22; \
        force U_IF_NAME.io_diffCommits_commitValid_23 = RTL_PATH.io_diffCommits_commitValid_23; \
        force U_IF_NAME.io_diffCommits_commitValid_24 = RTL_PATH.io_diffCommits_commitValid_24; \
        force U_IF_NAME.io_diffCommits_commitValid_25 = RTL_PATH.io_diffCommits_commitValid_25; \
        force U_IF_NAME.io_diffCommits_commitValid_26 = RTL_PATH.io_diffCommits_commitValid_26; \
        force U_IF_NAME.io_diffCommits_commitValid_27 = RTL_PATH.io_diffCommits_commitValid_27; \
        force U_IF_NAME.io_diffCommits_commitValid_28 = RTL_PATH.io_diffCommits_commitValid_28; \
        force U_IF_NAME.io_diffCommits_commitValid_29 = RTL_PATH.io_diffCommits_commitValid_29; \
        force U_IF_NAME.io_diffCommits_commitValid_30 = RTL_PATH.io_diffCommits_commitValid_30; \
        force U_IF_NAME.io_diffCommits_commitValid_31 = RTL_PATH.io_diffCommits_commitValid_31; \
        force U_IF_NAME.io_diffCommits_commitValid_32 = RTL_PATH.io_diffCommits_commitValid_32; \
        force U_IF_NAME.io_diffCommits_commitValid_33 = RTL_PATH.io_diffCommits_commitValid_33; \
        force U_IF_NAME.io_diffCommits_commitValid_34 = RTL_PATH.io_diffCommits_commitValid_34; \
        force U_IF_NAME.io_diffCommits_commitValid_35 = RTL_PATH.io_diffCommits_commitValid_35; \
        force U_IF_NAME.io_diffCommits_commitValid_36 = RTL_PATH.io_diffCommits_commitValid_36; \
        force U_IF_NAME.io_diffCommits_commitValid_37 = RTL_PATH.io_diffCommits_commitValid_37; \
        force U_IF_NAME.io_diffCommits_commitValid_38 = RTL_PATH.io_diffCommits_commitValid_38; \
        force U_IF_NAME.io_diffCommits_commitValid_39 = RTL_PATH.io_diffCommits_commitValid_39; \
        force U_IF_NAME.io_diffCommits_commitValid_40 = RTL_PATH.io_diffCommits_commitValid_40; \
        force U_IF_NAME.io_diffCommits_commitValid_41 = RTL_PATH.io_diffCommits_commitValid_41; \
        force U_IF_NAME.io_diffCommits_commitValid_42 = RTL_PATH.io_diffCommits_commitValid_42; \
        force U_IF_NAME.io_diffCommits_commitValid_43 = RTL_PATH.io_diffCommits_commitValid_43; \
        force U_IF_NAME.io_diffCommits_commitValid_44 = RTL_PATH.io_diffCommits_commitValid_44; \
        force U_IF_NAME.io_diffCommits_commitValid_45 = RTL_PATH.io_diffCommits_commitValid_45; \
        force U_IF_NAME.io_diffCommits_commitValid_46 = RTL_PATH.io_diffCommits_commitValid_46; \
        force U_IF_NAME.io_diffCommits_commitValid_47 = RTL_PATH.io_diffCommits_commitValid_47; \
        force U_IF_NAME.io_diffCommits_commitValid_48 = RTL_PATH.io_diffCommits_commitValid_48; \
        force U_IF_NAME.io_diffCommits_commitValid_49 = RTL_PATH.io_diffCommits_commitValid_49; \
        force U_IF_NAME.io_diffCommits_commitValid_50 = RTL_PATH.io_diffCommits_commitValid_50; \
        force U_IF_NAME.io_diffCommits_commitValid_51 = RTL_PATH.io_diffCommits_commitValid_51; \
        force U_IF_NAME.io_diffCommits_commitValid_52 = RTL_PATH.io_diffCommits_commitValid_52; \
        force U_IF_NAME.io_diffCommits_commitValid_53 = RTL_PATH.io_diffCommits_commitValid_53; \
        force U_IF_NAME.io_diffCommits_commitValid_54 = RTL_PATH.io_diffCommits_commitValid_54; \
        force U_IF_NAME.io_diffCommits_commitValid_55 = RTL_PATH.io_diffCommits_commitValid_55; \
        force U_IF_NAME.io_diffCommits_commitValid_56 = RTL_PATH.io_diffCommits_commitValid_56; \
        force U_IF_NAME.io_diffCommits_commitValid_57 = RTL_PATH.io_diffCommits_commitValid_57; \
        force U_IF_NAME.io_diffCommits_commitValid_58 = RTL_PATH.io_diffCommits_commitValid_58; \
        force U_IF_NAME.io_diffCommits_commitValid_59 = RTL_PATH.io_diffCommits_commitValid_59; \
        force U_IF_NAME.io_diffCommits_commitValid_60 = RTL_PATH.io_diffCommits_commitValid_60; \
        force U_IF_NAME.io_diffCommits_commitValid_61 = RTL_PATH.io_diffCommits_commitValid_61; \
        force U_IF_NAME.io_diffCommits_commitValid_62 = RTL_PATH.io_diffCommits_commitValid_62; \
        force U_IF_NAME.io_diffCommits_commitValid_63 = RTL_PATH.io_diffCommits_commitValid_63; \
        force U_IF_NAME.io_diffCommits_commitValid_64 = RTL_PATH.io_diffCommits_commitValid_64; \
        force U_IF_NAME.io_diffCommits_commitValid_65 = RTL_PATH.io_diffCommits_commitValid_65; \
        force U_IF_NAME.io_diffCommits_commitValid_66 = RTL_PATH.io_diffCommits_commitValid_66; \
        force U_IF_NAME.io_diffCommits_commitValid_67 = RTL_PATH.io_diffCommits_commitValid_67; \
        force U_IF_NAME.io_diffCommits_commitValid_68 = RTL_PATH.io_diffCommits_commitValid_68; \
        force U_IF_NAME.io_diffCommits_commitValid_69 = RTL_PATH.io_diffCommits_commitValid_69; \
        force U_IF_NAME.io_diffCommits_commitValid_70 = RTL_PATH.io_diffCommits_commitValid_70; \
        force U_IF_NAME.io_diffCommits_commitValid_71 = RTL_PATH.io_diffCommits_commitValid_71; \
        force U_IF_NAME.io_diffCommits_commitValid_72 = RTL_PATH.io_diffCommits_commitValid_72; \
        force U_IF_NAME.io_diffCommits_commitValid_73 = RTL_PATH.io_diffCommits_commitValid_73; \
        force U_IF_NAME.io_diffCommits_commitValid_74 = RTL_PATH.io_diffCommits_commitValid_74; \
        force U_IF_NAME.io_diffCommits_commitValid_75 = RTL_PATH.io_diffCommits_commitValid_75; \
        force U_IF_NAME.io_diffCommits_commitValid_76 = RTL_PATH.io_diffCommits_commitValid_76; \
        force U_IF_NAME.io_diffCommits_commitValid_77 = RTL_PATH.io_diffCommits_commitValid_77; \
        force U_IF_NAME.io_diffCommits_commitValid_78 = RTL_PATH.io_diffCommits_commitValid_78; \
        force U_IF_NAME.io_diffCommits_commitValid_79 = RTL_PATH.io_diffCommits_commitValid_79; \
        force U_IF_NAME.io_diffCommits_commitValid_80 = RTL_PATH.io_diffCommits_commitValid_80; \
        force U_IF_NAME.io_diffCommits_commitValid_81 = RTL_PATH.io_diffCommits_commitValid_81; \
        force U_IF_NAME.io_diffCommits_commitValid_82 = RTL_PATH.io_diffCommits_commitValid_82; \
        force U_IF_NAME.io_diffCommits_commitValid_83 = RTL_PATH.io_diffCommits_commitValid_83; \
        force U_IF_NAME.io_diffCommits_commitValid_84 = RTL_PATH.io_diffCommits_commitValid_84; \
        force U_IF_NAME.io_diffCommits_commitValid_85 = RTL_PATH.io_diffCommits_commitValid_85; \
        force U_IF_NAME.io_diffCommits_commitValid_86 = RTL_PATH.io_diffCommits_commitValid_86; \
        force U_IF_NAME.io_diffCommits_commitValid_87 = RTL_PATH.io_diffCommits_commitValid_87; \
        force U_IF_NAME.io_diffCommits_commitValid_88 = RTL_PATH.io_diffCommits_commitValid_88; \
        force U_IF_NAME.io_diffCommits_commitValid_89 = RTL_PATH.io_diffCommits_commitValid_89; \
        force U_IF_NAME.io_diffCommits_commitValid_90 = RTL_PATH.io_diffCommits_commitValid_90; \
        force U_IF_NAME.io_diffCommits_commitValid_91 = RTL_PATH.io_diffCommits_commitValid_91; \
        force U_IF_NAME.io_diffCommits_commitValid_92 = RTL_PATH.io_diffCommits_commitValid_92; \
        force U_IF_NAME.io_diffCommits_commitValid_93 = RTL_PATH.io_diffCommits_commitValid_93; \
        force U_IF_NAME.io_diffCommits_commitValid_94 = RTL_PATH.io_diffCommits_commitValid_94; \
        force U_IF_NAME.io_diffCommits_commitValid_95 = RTL_PATH.io_diffCommits_commitValid_95; \
        force U_IF_NAME.io_diffCommits_commitValid_96 = RTL_PATH.io_diffCommits_commitValid_96; \
        force U_IF_NAME.io_diffCommits_commitValid_97 = RTL_PATH.io_diffCommits_commitValid_97; \
        force U_IF_NAME.io_diffCommits_commitValid_98 = RTL_PATH.io_diffCommits_commitValid_98; \
        force U_IF_NAME.io_diffCommits_commitValid_99 = RTL_PATH.io_diffCommits_commitValid_99; \
        force U_IF_NAME.io_diffCommits_commitValid_100 = RTL_PATH.io_diffCommits_commitValid_100; \
        force U_IF_NAME.io_diffCommits_commitValid_101 = RTL_PATH.io_diffCommits_commitValid_101; \
        force U_IF_NAME.io_diffCommits_commitValid_102 = RTL_PATH.io_diffCommits_commitValid_102; \
        force U_IF_NAME.io_diffCommits_commitValid_103 = RTL_PATH.io_diffCommits_commitValid_103; \
        force U_IF_NAME.io_diffCommits_commitValid_104 = RTL_PATH.io_diffCommits_commitValid_104; \
        force U_IF_NAME.io_diffCommits_commitValid_105 = RTL_PATH.io_diffCommits_commitValid_105; \
        force U_IF_NAME.io_diffCommits_commitValid_106 = RTL_PATH.io_diffCommits_commitValid_106; \
        force U_IF_NAME.io_diffCommits_commitValid_107 = RTL_PATH.io_diffCommits_commitValid_107; \
        force U_IF_NAME.io_diffCommits_commitValid_108 = RTL_PATH.io_diffCommits_commitValid_108; \
        force U_IF_NAME.io_diffCommits_commitValid_109 = RTL_PATH.io_diffCommits_commitValid_109; \
        force U_IF_NAME.io_diffCommits_commitValid_110 = RTL_PATH.io_diffCommits_commitValid_110; \
        force U_IF_NAME.io_diffCommits_commitValid_111 = RTL_PATH.io_diffCommits_commitValid_111; \
        force U_IF_NAME.io_diffCommits_commitValid_112 = RTL_PATH.io_diffCommits_commitValid_112; \
        force U_IF_NAME.io_diffCommits_commitValid_113 = RTL_PATH.io_diffCommits_commitValid_113; \
        force U_IF_NAME.io_diffCommits_commitValid_114 = RTL_PATH.io_diffCommits_commitValid_114; \
        force U_IF_NAME.io_diffCommits_commitValid_115 = RTL_PATH.io_diffCommits_commitValid_115; \
        force U_IF_NAME.io_diffCommits_commitValid_116 = RTL_PATH.io_diffCommits_commitValid_116; \
        force U_IF_NAME.io_diffCommits_commitValid_117 = RTL_PATH.io_diffCommits_commitValid_117; \
        force U_IF_NAME.io_diffCommits_commitValid_118 = RTL_PATH.io_diffCommits_commitValid_118; \
        force U_IF_NAME.io_diffCommits_commitValid_119 = RTL_PATH.io_diffCommits_commitValid_119; \
        force U_IF_NAME.io_diffCommits_commitValid_120 = RTL_PATH.io_diffCommits_commitValid_120; \
        force U_IF_NAME.io_diffCommits_commitValid_121 = RTL_PATH.io_diffCommits_commitValid_121; \
        force U_IF_NAME.io_diffCommits_commitValid_122 = RTL_PATH.io_diffCommits_commitValid_122; \
        force U_IF_NAME.io_diffCommits_commitValid_123 = RTL_PATH.io_diffCommits_commitValid_123; \
        force U_IF_NAME.io_diffCommits_commitValid_124 = RTL_PATH.io_diffCommits_commitValid_124; \
        force U_IF_NAME.io_diffCommits_commitValid_125 = RTL_PATH.io_diffCommits_commitValid_125; \
        force U_IF_NAME.io_diffCommits_commitValid_126 = RTL_PATH.io_diffCommits_commitValid_126; \
        force U_IF_NAME.io_diffCommits_commitValid_127 = RTL_PATH.io_diffCommits_commitValid_127; \
        force U_IF_NAME.io_diffCommits_commitValid_128 = RTL_PATH.io_diffCommits_commitValid_128; \
        force U_IF_NAME.io_diffCommits_commitValid_129 = RTL_PATH.io_diffCommits_commitValid_129; \
        force U_IF_NAME.io_diffCommits_commitValid_130 = RTL_PATH.io_diffCommits_commitValid_130; \
        force U_IF_NAME.io_diffCommits_commitValid_131 = RTL_PATH.io_diffCommits_commitValid_131; \
        force U_IF_NAME.io_diffCommits_commitValid_132 = RTL_PATH.io_diffCommits_commitValid_132; \
        force U_IF_NAME.io_diffCommits_commitValid_133 = RTL_PATH.io_diffCommits_commitValid_133; \
        force U_IF_NAME.io_diffCommits_commitValid_134 = RTL_PATH.io_diffCommits_commitValid_134; \
        force U_IF_NAME.io_diffCommits_commitValid_135 = RTL_PATH.io_diffCommits_commitValid_135; \
        force U_IF_NAME.io_diffCommits_commitValid_136 = RTL_PATH.io_diffCommits_commitValid_136; \
        force U_IF_NAME.io_diffCommits_commitValid_137 = RTL_PATH.io_diffCommits_commitValid_137; \
        force U_IF_NAME.io_diffCommits_commitValid_138 = RTL_PATH.io_diffCommits_commitValid_138; \
        force U_IF_NAME.io_diffCommits_commitValid_139 = RTL_PATH.io_diffCommits_commitValid_139; \
        force U_IF_NAME.io_diffCommits_commitValid_140 = RTL_PATH.io_diffCommits_commitValid_140; \
        force U_IF_NAME.io_diffCommits_commitValid_141 = RTL_PATH.io_diffCommits_commitValid_141; \
        force U_IF_NAME.io_diffCommits_commitValid_142 = RTL_PATH.io_diffCommits_commitValid_142; \
        force U_IF_NAME.io_diffCommits_commitValid_143 = RTL_PATH.io_diffCommits_commitValid_143; \
        force U_IF_NAME.io_diffCommits_commitValid_144 = RTL_PATH.io_diffCommits_commitValid_144; \
        force U_IF_NAME.io_diffCommits_commitValid_145 = RTL_PATH.io_diffCommits_commitValid_145; \
        force U_IF_NAME.io_diffCommits_commitValid_146 = RTL_PATH.io_diffCommits_commitValid_146; \
        force U_IF_NAME.io_diffCommits_commitValid_147 = RTL_PATH.io_diffCommits_commitValid_147; \
        force U_IF_NAME.io_diffCommits_commitValid_148 = RTL_PATH.io_diffCommits_commitValid_148; \
        force U_IF_NAME.io_diffCommits_commitValid_149 = RTL_PATH.io_diffCommits_commitValid_149; \
        force U_IF_NAME.io_diffCommits_commitValid_150 = RTL_PATH.io_diffCommits_commitValid_150; \
        force U_IF_NAME.io_diffCommits_commitValid_151 = RTL_PATH.io_diffCommits_commitValid_151; \
        force U_IF_NAME.io_diffCommits_commitValid_152 = RTL_PATH.io_diffCommits_commitValid_152; \
        force U_IF_NAME.io_diffCommits_commitValid_153 = RTL_PATH.io_diffCommits_commitValid_153; \
        force U_IF_NAME.io_diffCommits_commitValid_154 = RTL_PATH.io_diffCommits_commitValid_154; \
        force U_IF_NAME.io_diffCommits_commitValid_155 = RTL_PATH.io_diffCommits_commitValid_155; \
        force U_IF_NAME.io_diffCommits_commitValid_156 = RTL_PATH.io_diffCommits_commitValid_156; \
        force U_IF_NAME.io_diffCommits_commitValid_157 = RTL_PATH.io_diffCommits_commitValid_157; \
        force U_IF_NAME.io_diffCommits_commitValid_158 = RTL_PATH.io_diffCommits_commitValid_158; \
        force U_IF_NAME.io_diffCommits_commitValid_159 = RTL_PATH.io_diffCommits_commitValid_159; \
        force U_IF_NAME.io_diffCommits_commitValid_160 = RTL_PATH.io_diffCommits_commitValid_160; \
        force U_IF_NAME.io_diffCommits_commitValid_161 = RTL_PATH.io_diffCommits_commitValid_161; \
        force U_IF_NAME.io_diffCommits_commitValid_162 = RTL_PATH.io_diffCommits_commitValid_162; \
        force U_IF_NAME.io_diffCommits_commitValid_163 = RTL_PATH.io_diffCommits_commitValid_163; \
        force U_IF_NAME.io_diffCommits_commitValid_164 = RTL_PATH.io_diffCommits_commitValid_164; \
        force U_IF_NAME.io_diffCommits_commitValid_165 = RTL_PATH.io_diffCommits_commitValid_165; \
        force U_IF_NAME.io_diffCommits_commitValid_166 = RTL_PATH.io_diffCommits_commitValid_166; \
        force U_IF_NAME.io_diffCommits_commitValid_167 = RTL_PATH.io_diffCommits_commitValid_167; \
        force U_IF_NAME.io_diffCommits_commitValid_168 = RTL_PATH.io_diffCommits_commitValid_168; \
        force U_IF_NAME.io_diffCommits_commitValid_169 = RTL_PATH.io_diffCommits_commitValid_169; \
        force U_IF_NAME.io_diffCommits_commitValid_170 = RTL_PATH.io_diffCommits_commitValid_170; \
        force U_IF_NAME.io_diffCommits_commitValid_171 = RTL_PATH.io_diffCommits_commitValid_171; \
        force U_IF_NAME.io_diffCommits_commitValid_172 = RTL_PATH.io_diffCommits_commitValid_172; \
        force U_IF_NAME.io_diffCommits_commitValid_173 = RTL_PATH.io_diffCommits_commitValid_173; \
        force U_IF_NAME.io_diffCommits_commitValid_174 = RTL_PATH.io_diffCommits_commitValid_174; \
        force U_IF_NAME.io_diffCommits_commitValid_175 = RTL_PATH.io_diffCommits_commitValid_175; \
        force U_IF_NAME.io_diffCommits_commitValid_176 = RTL_PATH.io_diffCommits_commitValid_176; \
        force U_IF_NAME.io_diffCommits_commitValid_177 = RTL_PATH.io_diffCommits_commitValid_177; \
        force U_IF_NAME.io_diffCommits_commitValid_178 = RTL_PATH.io_diffCommits_commitValid_178; \
        force U_IF_NAME.io_diffCommits_commitValid_179 = RTL_PATH.io_diffCommits_commitValid_179; \
        force U_IF_NAME.io_diffCommits_commitValid_180 = RTL_PATH.io_diffCommits_commitValid_180; \
        force U_IF_NAME.io_diffCommits_commitValid_181 = RTL_PATH.io_diffCommits_commitValid_181; \
        force U_IF_NAME.io_diffCommits_commitValid_182 = RTL_PATH.io_diffCommits_commitValid_182; \
        force U_IF_NAME.io_diffCommits_commitValid_183 = RTL_PATH.io_diffCommits_commitValid_183; \
        force U_IF_NAME.io_diffCommits_commitValid_184 = RTL_PATH.io_diffCommits_commitValid_184; \
        force U_IF_NAME.io_diffCommits_commitValid_185 = RTL_PATH.io_diffCommits_commitValid_185; \
        force U_IF_NAME.io_diffCommits_commitValid_186 = RTL_PATH.io_diffCommits_commitValid_186; \
        force U_IF_NAME.io_diffCommits_commitValid_187 = RTL_PATH.io_diffCommits_commitValid_187; \
        force U_IF_NAME.io_diffCommits_commitValid_188 = RTL_PATH.io_diffCommits_commitValid_188; \
        force U_IF_NAME.io_diffCommits_commitValid_189 = RTL_PATH.io_diffCommits_commitValid_189; \
        force U_IF_NAME.io_diffCommits_commitValid_190 = RTL_PATH.io_diffCommits_commitValid_190; \
        force U_IF_NAME.io_diffCommits_commitValid_191 = RTL_PATH.io_diffCommits_commitValid_191; \
        force U_IF_NAME.io_diffCommits_commitValid_192 = RTL_PATH.io_diffCommits_commitValid_192; \
        force U_IF_NAME.io_diffCommits_commitValid_193 = RTL_PATH.io_diffCommits_commitValid_193; \
        force U_IF_NAME.io_diffCommits_commitValid_194 = RTL_PATH.io_diffCommits_commitValid_194; \
        force U_IF_NAME.io_diffCommits_commitValid_195 = RTL_PATH.io_diffCommits_commitValid_195; \
        force U_IF_NAME.io_diffCommits_commitValid_196 = RTL_PATH.io_diffCommits_commitValid_196; \
        force U_IF_NAME.io_diffCommits_commitValid_197 = RTL_PATH.io_diffCommits_commitValid_197; \
        force U_IF_NAME.io_diffCommits_commitValid_198 = RTL_PATH.io_diffCommits_commitValid_198; \
        force U_IF_NAME.io_diffCommits_commitValid_199 = RTL_PATH.io_diffCommits_commitValid_199; \
        force U_IF_NAME.io_diffCommits_commitValid_200 = RTL_PATH.io_diffCommits_commitValid_200; \
        force U_IF_NAME.io_diffCommits_commitValid_201 = RTL_PATH.io_diffCommits_commitValid_201; \
        force U_IF_NAME.io_diffCommits_commitValid_202 = RTL_PATH.io_diffCommits_commitValid_202; \
        force U_IF_NAME.io_diffCommits_commitValid_203 = RTL_PATH.io_diffCommits_commitValid_203; \
        force U_IF_NAME.io_diffCommits_commitValid_204 = RTL_PATH.io_diffCommits_commitValid_204; \
        force U_IF_NAME.io_diffCommits_commitValid_205 = RTL_PATH.io_diffCommits_commitValid_205; \
        force U_IF_NAME.io_diffCommits_commitValid_206 = RTL_PATH.io_diffCommits_commitValid_206; \
        force U_IF_NAME.io_diffCommits_commitValid_207 = RTL_PATH.io_diffCommits_commitValid_207; \
        force U_IF_NAME.io_diffCommits_commitValid_208 = RTL_PATH.io_diffCommits_commitValid_208; \
        force U_IF_NAME.io_diffCommits_commitValid_209 = RTL_PATH.io_diffCommits_commitValid_209; \
        force U_IF_NAME.io_diffCommits_commitValid_210 = RTL_PATH.io_diffCommits_commitValid_210; \
        force U_IF_NAME.io_diffCommits_commitValid_211 = RTL_PATH.io_diffCommits_commitValid_211; \
        force U_IF_NAME.io_diffCommits_commitValid_212 = RTL_PATH.io_diffCommits_commitValid_212; \
        force U_IF_NAME.io_diffCommits_commitValid_213 = RTL_PATH.io_diffCommits_commitValid_213; \
        force U_IF_NAME.io_diffCommits_commitValid_214 = RTL_PATH.io_diffCommits_commitValid_214; \
        force U_IF_NAME.io_diffCommits_commitValid_215 = RTL_PATH.io_diffCommits_commitValid_215; \
        force U_IF_NAME.io_diffCommits_commitValid_216 = RTL_PATH.io_diffCommits_commitValid_216; \
        force U_IF_NAME.io_diffCommits_commitValid_217 = RTL_PATH.io_diffCommits_commitValid_217; \
        force U_IF_NAME.io_diffCommits_commitValid_218 = RTL_PATH.io_diffCommits_commitValid_218; \
        force U_IF_NAME.io_diffCommits_commitValid_219 = RTL_PATH.io_diffCommits_commitValid_219; \
        force U_IF_NAME.io_diffCommits_commitValid_220 = RTL_PATH.io_diffCommits_commitValid_220; \
        force U_IF_NAME.io_diffCommits_commitValid_221 = RTL_PATH.io_diffCommits_commitValid_221; \
        force U_IF_NAME.io_diffCommits_commitValid_222 = RTL_PATH.io_diffCommits_commitValid_222; \
        force U_IF_NAME.io_diffCommits_commitValid_223 = RTL_PATH.io_diffCommits_commitValid_223; \
        force U_IF_NAME.io_diffCommits_commitValid_224 = RTL_PATH.io_diffCommits_commitValid_224; \
        force U_IF_NAME.io_diffCommits_commitValid_225 = RTL_PATH.io_diffCommits_commitValid_225; \
        force U_IF_NAME.io_diffCommits_commitValid_226 = RTL_PATH.io_diffCommits_commitValid_226; \
        force U_IF_NAME.io_diffCommits_commitValid_227 = RTL_PATH.io_diffCommits_commitValid_227; \
        force U_IF_NAME.io_diffCommits_commitValid_228 = RTL_PATH.io_diffCommits_commitValid_228; \
        force U_IF_NAME.io_diffCommits_commitValid_229 = RTL_PATH.io_diffCommits_commitValid_229; \
        force U_IF_NAME.io_diffCommits_commitValid_230 = RTL_PATH.io_diffCommits_commitValid_230; \
        force U_IF_NAME.io_diffCommits_commitValid_231 = RTL_PATH.io_diffCommits_commitValid_231; \
        force U_IF_NAME.io_diffCommits_commitValid_232 = RTL_PATH.io_diffCommits_commitValid_232; \
        force U_IF_NAME.io_diffCommits_commitValid_233 = RTL_PATH.io_diffCommits_commitValid_233; \
        force U_IF_NAME.io_diffCommits_commitValid_234 = RTL_PATH.io_diffCommits_commitValid_234; \
        force U_IF_NAME.io_diffCommits_commitValid_235 = RTL_PATH.io_diffCommits_commitValid_235; \
        force U_IF_NAME.io_diffCommits_commitValid_236 = RTL_PATH.io_diffCommits_commitValid_236; \
        force U_IF_NAME.io_diffCommits_commitValid_237 = RTL_PATH.io_diffCommits_commitValid_237; \
        force U_IF_NAME.io_diffCommits_commitValid_238 = RTL_PATH.io_diffCommits_commitValid_238; \
        force U_IF_NAME.io_diffCommits_commitValid_239 = RTL_PATH.io_diffCommits_commitValid_239; \
        force U_IF_NAME.io_diffCommits_commitValid_240 = RTL_PATH.io_diffCommits_commitValid_240; \
        force U_IF_NAME.io_diffCommits_commitValid_241 = RTL_PATH.io_diffCommits_commitValid_241; \
        force U_IF_NAME.io_diffCommits_commitValid_242 = RTL_PATH.io_diffCommits_commitValid_242; \
        force U_IF_NAME.io_diffCommits_commitValid_243 = RTL_PATH.io_diffCommits_commitValid_243; \
        force U_IF_NAME.io_diffCommits_commitValid_244 = RTL_PATH.io_diffCommits_commitValid_244; \
        force U_IF_NAME.io_diffCommits_commitValid_245 = RTL_PATH.io_diffCommits_commitValid_245; \
        force U_IF_NAME.io_diffCommits_commitValid_246 = RTL_PATH.io_diffCommits_commitValid_246; \
        force U_IF_NAME.io_diffCommits_commitValid_247 = RTL_PATH.io_diffCommits_commitValid_247; \
        force U_IF_NAME.io_diffCommits_commitValid_248 = RTL_PATH.io_diffCommits_commitValid_248; \
        force U_IF_NAME.io_diffCommits_commitValid_249 = RTL_PATH.io_diffCommits_commitValid_249; \
        force U_IF_NAME.io_diffCommits_commitValid_250 = RTL_PATH.io_diffCommits_commitValid_250; \
        force U_IF_NAME.io_diffCommits_commitValid_251 = RTL_PATH.io_diffCommits_commitValid_251; \
        force U_IF_NAME.io_diffCommits_commitValid_252 = RTL_PATH.io_diffCommits_commitValid_252; \
        force U_IF_NAME.io_diffCommits_commitValid_253 = RTL_PATH.io_diffCommits_commitValid_253; \
        force U_IF_NAME.io_diffCommits_commitValid_254 = RTL_PATH.io_diffCommits_commitValid_254; \
        force U_IF_NAME.io_diffCommits_info_0_ldest = RTL_PATH.io_diffCommits_info_0_ldest; \
        force U_IF_NAME.io_diffCommits_info_0_pdest = RTL_PATH.io_diffCommits_info_0_pdest; \
        force U_IF_NAME.io_diffCommits_info_0_rfWen = RTL_PATH.io_diffCommits_info_0_rfWen; \
        force U_IF_NAME.io_diffCommits_info_0_fpWen = RTL_PATH.io_diffCommits_info_0_fpWen; \
        force U_IF_NAME.io_diffCommits_info_0_vecWen = RTL_PATH.io_diffCommits_info_0_vecWen; \
        force U_IF_NAME.io_diffCommits_info_0_v0Wen = RTL_PATH.io_diffCommits_info_0_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_0_vlWen = RTL_PATH.io_diffCommits_info_0_vlWen; \
        force U_IF_NAME.io_diffCommits_info_1_ldest = RTL_PATH.io_diffCommits_info_1_ldest; \
        force U_IF_NAME.io_diffCommits_info_1_pdest = RTL_PATH.io_diffCommits_info_1_pdest; \
        force U_IF_NAME.io_diffCommits_info_1_rfWen = RTL_PATH.io_diffCommits_info_1_rfWen; \
        force U_IF_NAME.io_diffCommits_info_1_fpWen = RTL_PATH.io_diffCommits_info_1_fpWen; \
        force U_IF_NAME.io_diffCommits_info_1_vecWen = RTL_PATH.io_diffCommits_info_1_vecWen; \
        force U_IF_NAME.io_diffCommits_info_1_v0Wen = RTL_PATH.io_diffCommits_info_1_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_1_vlWen = RTL_PATH.io_diffCommits_info_1_vlWen; \
        force U_IF_NAME.io_diffCommits_info_2_ldest = RTL_PATH.io_diffCommits_info_2_ldest; \
        force U_IF_NAME.io_diffCommits_info_2_pdest = RTL_PATH.io_diffCommits_info_2_pdest; \
        force U_IF_NAME.io_diffCommits_info_2_rfWen = RTL_PATH.io_diffCommits_info_2_rfWen; \
        force U_IF_NAME.io_diffCommits_info_2_fpWen = RTL_PATH.io_diffCommits_info_2_fpWen; \
        force U_IF_NAME.io_diffCommits_info_2_vecWen = RTL_PATH.io_diffCommits_info_2_vecWen; \
        force U_IF_NAME.io_diffCommits_info_2_v0Wen = RTL_PATH.io_diffCommits_info_2_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_2_vlWen = RTL_PATH.io_diffCommits_info_2_vlWen; \
        force U_IF_NAME.io_diffCommits_info_3_ldest = RTL_PATH.io_diffCommits_info_3_ldest; \
        force U_IF_NAME.io_diffCommits_info_3_pdest = RTL_PATH.io_diffCommits_info_3_pdest; \
        force U_IF_NAME.io_diffCommits_info_3_rfWen = RTL_PATH.io_diffCommits_info_3_rfWen; \
        force U_IF_NAME.io_diffCommits_info_3_fpWen = RTL_PATH.io_diffCommits_info_3_fpWen; \
        force U_IF_NAME.io_diffCommits_info_3_vecWen = RTL_PATH.io_diffCommits_info_3_vecWen; \
        force U_IF_NAME.io_diffCommits_info_3_v0Wen = RTL_PATH.io_diffCommits_info_3_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_3_vlWen = RTL_PATH.io_diffCommits_info_3_vlWen; \
        force U_IF_NAME.io_diffCommits_info_4_ldest = RTL_PATH.io_diffCommits_info_4_ldest; \
        force U_IF_NAME.io_diffCommits_info_4_pdest = RTL_PATH.io_diffCommits_info_4_pdest; \
        force U_IF_NAME.io_diffCommits_info_4_rfWen = RTL_PATH.io_diffCommits_info_4_rfWen; \
        force U_IF_NAME.io_diffCommits_info_4_fpWen = RTL_PATH.io_diffCommits_info_4_fpWen; \
        force U_IF_NAME.io_diffCommits_info_4_vecWen = RTL_PATH.io_diffCommits_info_4_vecWen; \
        force U_IF_NAME.io_diffCommits_info_4_v0Wen = RTL_PATH.io_diffCommits_info_4_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_4_vlWen = RTL_PATH.io_diffCommits_info_4_vlWen; \
        force U_IF_NAME.io_diffCommits_info_5_ldest = RTL_PATH.io_diffCommits_info_5_ldest; \
        force U_IF_NAME.io_diffCommits_info_5_pdest = RTL_PATH.io_diffCommits_info_5_pdest; \
        force U_IF_NAME.io_diffCommits_info_5_rfWen = RTL_PATH.io_diffCommits_info_5_rfWen; \
        force U_IF_NAME.io_diffCommits_info_5_fpWen = RTL_PATH.io_diffCommits_info_5_fpWen; \
        force U_IF_NAME.io_diffCommits_info_5_vecWen = RTL_PATH.io_diffCommits_info_5_vecWen; \
        force U_IF_NAME.io_diffCommits_info_5_v0Wen = RTL_PATH.io_diffCommits_info_5_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_5_vlWen = RTL_PATH.io_diffCommits_info_5_vlWen; \
        force U_IF_NAME.io_diffCommits_info_6_ldest = RTL_PATH.io_diffCommits_info_6_ldest; \
        force U_IF_NAME.io_diffCommits_info_6_pdest = RTL_PATH.io_diffCommits_info_6_pdest; \
        force U_IF_NAME.io_diffCommits_info_6_rfWen = RTL_PATH.io_diffCommits_info_6_rfWen; \
        force U_IF_NAME.io_diffCommits_info_6_fpWen = RTL_PATH.io_diffCommits_info_6_fpWen; \
        force U_IF_NAME.io_diffCommits_info_6_vecWen = RTL_PATH.io_diffCommits_info_6_vecWen; \
        force U_IF_NAME.io_diffCommits_info_6_v0Wen = RTL_PATH.io_diffCommits_info_6_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_6_vlWen = RTL_PATH.io_diffCommits_info_6_vlWen; \
        force U_IF_NAME.io_diffCommits_info_7_ldest = RTL_PATH.io_diffCommits_info_7_ldest; \
        force U_IF_NAME.io_diffCommits_info_7_pdest = RTL_PATH.io_diffCommits_info_7_pdest; \
        force U_IF_NAME.io_diffCommits_info_7_rfWen = RTL_PATH.io_diffCommits_info_7_rfWen; \
        force U_IF_NAME.io_diffCommits_info_7_fpWen = RTL_PATH.io_diffCommits_info_7_fpWen; \
        force U_IF_NAME.io_diffCommits_info_7_vecWen = RTL_PATH.io_diffCommits_info_7_vecWen; \
        force U_IF_NAME.io_diffCommits_info_7_v0Wen = RTL_PATH.io_diffCommits_info_7_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_7_vlWen = RTL_PATH.io_diffCommits_info_7_vlWen; \
        force U_IF_NAME.io_diffCommits_info_8_ldest = RTL_PATH.io_diffCommits_info_8_ldest; \
        force U_IF_NAME.io_diffCommits_info_8_pdest = RTL_PATH.io_diffCommits_info_8_pdest; \
        force U_IF_NAME.io_diffCommits_info_8_rfWen = RTL_PATH.io_diffCommits_info_8_rfWen; \
        force U_IF_NAME.io_diffCommits_info_8_fpWen = RTL_PATH.io_diffCommits_info_8_fpWen; \
        force U_IF_NAME.io_diffCommits_info_8_vecWen = RTL_PATH.io_diffCommits_info_8_vecWen; \
        force U_IF_NAME.io_diffCommits_info_8_v0Wen = RTL_PATH.io_diffCommits_info_8_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_8_vlWen = RTL_PATH.io_diffCommits_info_8_vlWen; \
        force U_IF_NAME.io_diffCommits_info_9_ldest = RTL_PATH.io_diffCommits_info_9_ldest; \
        force U_IF_NAME.io_diffCommits_info_9_pdest = RTL_PATH.io_diffCommits_info_9_pdest; \
        force U_IF_NAME.io_diffCommits_info_9_rfWen = RTL_PATH.io_diffCommits_info_9_rfWen; \
        force U_IF_NAME.io_diffCommits_info_9_fpWen = RTL_PATH.io_diffCommits_info_9_fpWen; \
        force U_IF_NAME.io_diffCommits_info_9_vecWen = RTL_PATH.io_diffCommits_info_9_vecWen; \
        force U_IF_NAME.io_diffCommits_info_9_v0Wen = RTL_PATH.io_diffCommits_info_9_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_9_vlWen = RTL_PATH.io_diffCommits_info_9_vlWen; \
        force U_IF_NAME.io_diffCommits_info_10_ldest = RTL_PATH.io_diffCommits_info_10_ldest; \
        force U_IF_NAME.io_diffCommits_info_10_pdest = RTL_PATH.io_diffCommits_info_10_pdest; \
        force U_IF_NAME.io_diffCommits_info_10_rfWen = RTL_PATH.io_diffCommits_info_10_rfWen; \
        force U_IF_NAME.io_diffCommits_info_10_fpWen = RTL_PATH.io_diffCommits_info_10_fpWen; \
        force U_IF_NAME.io_diffCommits_info_10_vecWen = RTL_PATH.io_diffCommits_info_10_vecWen; \
        force U_IF_NAME.io_diffCommits_info_10_v0Wen = RTL_PATH.io_diffCommits_info_10_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_10_vlWen = RTL_PATH.io_diffCommits_info_10_vlWen; \
        force U_IF_NAME.io_diffCommits_info_11_ldest = RTL_PATH.io_diffCommits_info_11_ldest; \
        force U_IF_NAME.io_diffCommits_info_11_pdest = RTL_PATH.io_diffCommits_info_11_pdest; \
        force U_IF_NAME.io_diffCommits_info_11_rfWen = RTL_PATH.io_diffCommits_info_11_rfWen; \
        force U_IF_NAME.io_diffCommits_info_11_fpWen = RTL_PATH.io_diffCommits_info_11_fpWen; \
        force U_IF_NAME.io_diffCommits_info_11_vecWen = RTL_PATH.io_diffCommits_info_11_vecWen; \
        force U_IF_NAME.io_diffCommits_info_11_v0Wen = RTL_PATH.io_diffCommits_info_11_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_11_vlWen = RTL_PATH.io_diffCommits_info_11_vlWen; \
        force U_IF_NAME.io_diffCommits_info_12_ldest = RTL_PATH.io_diffCommits_info_12_ldest; \
        force U_IF_NAME.io_diffCommits_info_12_pdest = RTL_PATH.io_diffCommits_info_12_pdest; \
        force U_IF_NAME.io_diffCommits_info_12_rfWen = RTL_PATH.io_diffCommits_info_12_rfWen; \
        force U_IF_NAME.io_diffCommits_info_12_fpWen = RTL_PATH.io_diffCommits_info_12_fpWen; \
        force U_IF_NAME.io_diffCommits_info_12_vecWen = RTL_PATH.io_diffCommits_info_12_vecWen; \
        force U_IF_NAME.io_diffCommits_info_12_v0Wen = RTL_PATH.io_diffCommits_info_12_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_12_vlWen = RTL_PATH.io_diffCommits_info_12_vlWen; \
        force U_IF_NAME.io_diffCommits_info_13_ldest = RTL_PATH.io_diffCommits_info_13_ldest; \
        force U_IF_NAME.io_diffCommits_info_13_pdest = RTL_PATH.io_diffCommits_info_13_pdest; \
        force U_IF_NAME.io_diffCommits_info_13_rfWen = RTL_PATH.io_diffCommits_info_13_rfWen; \
        force U_IF_NAME.io_diffCommits_info_13_fpWen = RTL_PATH.io_diffCommits_info_13_fpWen; \
        force U_IF_NAME.io_diffCommits_info_13_vecWen = RTL_PATH.io_diffCommits_info_13_vecWen; \
        force U_IF_NAME.io_diffCommits_info_13_v0Wen = RTL_PATH.io_diffCommits_info_13_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_13_vlWen = RTL_PATH.io_diffCommits_info_13_vlWen; \
        force U_IF_NAME.io_diffCommits_info_14_ldest = RTL_PATH.io_diffCommits_info_14_ldest; \
        force U_IF_NAME.io_diffCommits_info_14_pdest = RTL_PATH.io_diffCommits_info_14_pdest; \
        force U_IF_NAME.io_diffCommits_info_14_rfWen = RTL_PATH.io_diffCommits_info_14_rfWen; \
        force U_IF_NAME.io_diffCommits_info_14_fpWen = RTL_PATH.io_diffCommits_info_14_fpWen; \
        force U_IF_NAME.io_diffCommits_info_14_vecWen = RTL_PATH.io_diffCommits_info_14_vecWen; \
        force U_IF_NAME.io_diffCommits_info_14_v0Wen = RTL_PATH.io_diffCommits_info_14_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_14_vlWen = RTL_PATH.io_diffCommits_info_14_vlWen; \
        force U_IF_NAME.io_diffCommits_info_15_ldest = RTL_PATH.io_diffCommits_info_15_ldest; \
        force U_IF_NAME.io_diffCommits_info_15_pdest = RTL_PATH.io_diffCommits_info_15_pdest; \
        force U_IF_NAME.io_diffCommits_info_15_rfWen = RTL_PATH.io_diffCommits_info_15_rfWen; \
        force U_IF_NAME.io_diffCommits_info_15_fpWen = RTL_PATH.io_diffCommits_info_15_fpWen; \
        force U_IF_NAME.io_diffCommits_info_15_vecWen = RTL_PATH.io_diffCommits_info_15_vecWen; \
        force U_IF_NAME.io_diffCommits_info_15_v0Wen = RTL_PATH.io_diffCommits_info_15_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_15_vlWen = RTL_PATH.io_diffCommits_info_15_vlWen; \
        force U_IF_NAME.io_diffCommits_info_16_ldest = RTL_PATH.io_diffCommits_info_16_ldest; \
        force U_IF_NAME.io_diffCommits_info_16_pdest = RTL_PATH.io_diffCommits_info_16_pdest; \
        force U_IF_NAME.io_diffCommits_info_16_rfWen = RTL_PATH.io_diffCommits_info_16_rfWen; \
        force U_IF_NAME.io_diffCommits_info_16_fpWen = RTL_PATH.io_diffCommits_info_16_fpWen; \
        force U_IF_NAME.io_diffCommits_info_16_vecWen = RTL_PATH.io_diffCommits_info_16_vecWen; \
        force U_IF_NAME.io_diffCommits_info_16_v0Wen = RTL_PATH.io_diffCommits_info_16_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_16_vlWen = RTL_PATH.io_diffCommits_info_16_vlWen; \
        force U_IF_NAME.io_diffCommits_info_17_ldest = RTL_PATH.io_diffCommits_info_17_ldest; \
        force U_IF_NAME.io_diffCommits_info_17_pdest = RTL_PATH.io_diffCommits_info_17_pdest; \
        force U_IF_NAME.io_diffCommits_info_17_rfWen = RTL_PATH.io_diffCommits_info_17_rfWen; \
        force U_IF_NAME.io_diffCommits_info_17_fpWen = RTL_PATH.io_diffCommits_info_17_fpWen; \
        force U_IF_NAME.io_diffCommits_info_17_vecWen = RTL_PATH.io_diffCommits_info_17_vecWen; \
        force U_IF_NAME.io_diffCommits_info_17_v0Wen = RTL_PATH.io_diffCommits_info_17_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_17_vlWen = RTL_PATH.io_diffCommits_info_17_vlWen; \
        force U_IF_NAME.io_diffCommits_info_18_ldest = RTL_PATH.io_diffCommits_info_18_ldest; \
        force U_IF_NAME.io_diffCommits_info_18_pdest = RTL_PATH.io_diffCommits_info_18_pdest; \
        force U_IF_NAME.io_diffCommits_info_18_rfWen = RTL_PATH.io_diffCommits_info_18_rfWen; \
        force U_IF_NAME.io_diffCommits_info_18_fpWen = RTL_PATH.io_diffCommits_info_18_fpWen; \
        force U_IF_NAME.io_diffCommits_info_18_vecWen = RTL_PATH.io_diffCommits_info_18_vecWen; \
        force U_IF_NAME.io_diffCommits_info_18_v0Wen = RTL_PATH.io_diffCommits_info_18_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_18_vlWen = RTL_PATH.io_diffCommits_info_18_vlWen; \
        force U_IF_NAME.io_diffCommits_info_19_ldest = RTL_PATH.io_diffCommits_info_19_ldest; \
        force U_IF_NAME.io_diffCommits_info_19_pdest = RTL_PATH.io_diffCommits_info_19_pdest; \
        force U_IF_NAME.io_diffCommits_info_19_rfWen = RTL_PATH.io_diffCommits_info_19_rfWen; \
        force U_IF_NAME.io_diffCommits_info_19_fpWen = RTL_PATH.io_diffCommits_info_19_fpWen; \
        force U_IF_NAME.io_diffCommits_info_19_vecWen = RTL_PATH.io_diffCommits_info_19_vecWen; \
        force U_IF_NAME.io_diffCommits_info_19_v0Wen = RTL_PATH.io_diffCommits_info_19_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_19_vlWen = RTL_PATH.io_diffCommits_info_19_vlWen; \
        force U_IF_NAME.io_diffCommits_info_20_ldest = RTL_PATH.io_diffCommits_info_20_ldest; \
        force U_IF_NAME.io_diffCommits_info_20_pdest = RTL_PATH.io_diffCommits_info_20_pdest; \
        force U_IF_NAME.io_diffCommits_info_20_rfWen = RTL_PATH.io_diffCommits_info_20_rfWen; \
        force U_IF_NAME.io_diffCommits_info_20_fpWen = RTL_PATH.io_diffCommits_info_20_fpWen; \
        force U_IF_NAME.io_diffCommits_info_20_vecWen = RTL_PATH.io_diffCommits_info_20_vecWen; \
        force U_IF_NAME.io_diffCommits_info_20_v0Wen = RTL_PATH.io_diffCommits_info_20_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_20_vlWen = RTL_PATH.io_diffCommits_info_20_vlWen; \
        force U_IF_NAME.io_diffCommits_info_21_ldest = RTL_PATH.io_diffCommits_info_21_ldest; \
        force U_IF_NAME.io_diffCommits_info_21_pdest = RTL_PATH.io_diffCommits_info_21_pdest; \
        force U_IF_NAME.io_diffCommits_info_21_rfWen = RTL_PATH.io_diffCommits_info_21_rfWen; \
        force U_IF_NAME.io_diffCommits_info_21_fpWen = RTL_PATH.io_diffCommits_info_21_fpWen; \
        force U_IF_NAME.io_diffCommits_info_21_vecWen = RTL_PATH.io_diffCommits_info_21_vecWen; \
        force U_IF_NAME.io_diffCommits_info_21_v0Wen = RTL_PATH.io_diffCommits_info_21_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_21_vlWen = RTL_PATH.io_diffCommits_info_21_vlWen; \
        force U_IF_NAME.io_diffCommits_info_22_ldest = RTL_PATH.io_diffCommits_info_22_ldest; \
        force U_IF_NAME.io_diffCommits_info_22_pdest = RTL_PATH.io_diffCommits_info_22_pdest; \
        force U_IF_NAME.io_diffCommits_info_22_rfWen = RTL_PATH.io_diffCommits_info_22_rfWen; \
        force U_IF_NAME.io_diffCommits_info_22_fpWen = RTL_PATH.io_diffCommits_info_22_fpWen; \
        force U_IF_NAME.io_diffCommits_info_22_vecWen = RTL_PATH.io_diffCommits_info_22_vecWen; \
        force U_IF_NAME.io_diffCommits_info_22_v0Wen = RTL_PATH.io_diffCommits_info_22_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_22_vlWen = RTL_PATH.io_diffCommits_info_22_vlWen; \
        force U_IF_NAME.io_diffCommits_info_23_ldest = RTL_PATH.io_diffCommits_info_23_ldest; \
        force U_IF_NAME.io_diffCommits_info_23_pdest = RTL_PATH.io_diffCommits_info_23_pdest; \
        force U_IF_NAME.io_diffCommits_info_23_rfWen = RTL_PATH.io_diffCommits_info_23_rfWen; \
        force U_IF_NAME.io_diffCommits_info_23_fpWen = RTL_PATH.io_diffCommits_info_23_fpWen; \
        force U_IF_NAME.io_diffCommits_info_23_vecWen = RTL_PATH.io_diffCommits_info_23_vecWen; \
        force U_IF_NAME.io_diffCommits_info_23_v0Wen = RTL_PATH.io_diffCommits_info_23_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_23_vlWen = RTL_PATH.io_diffCommits_info_23_vlWen; \
        force U_IF_NAME.io_diffCommits_info_24_ldest = RTL_PATH.io_diffCommits_info_24_ldest; \
        force U_IF_NAME.io_diffCommits_info_24_pdest = RTL_PATH.io_diffCommits_info_24_pdest; \
        force U_IF_NAME.io_diffCommits_info_24_rfWen = RTL_PATH.io_diffCommits_info_24_rfWen; \
        force U_IF_NAME.io_diffCommits_info_24_fpWen = RTL_PATH.io_diffCommits_info_24_fpWen; \
        force U_IF_NAME.io_diffCommits_info_24_vecWen = RTL_PATH.io_diffCommits_info_24_vecWen; \
        force U_IF_NAME.io_diffCommits_info_24_v0Wen = RTL_PATH.io_diffCommits_info_24_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_24_vlWen = RTL_PATH.io_diffCommits_info_24_vlWen; \
        force U_IF_NAME.io_diffCommits_info_25_ldest = RTL_PATH.io_diffCommits_info_25_ldest; \
        force U_IF_NAME.io_diffCommits_info_25_pdest = RTL_PATH.io_diffCommits_info_25_pdest; \
        force U_IF_NAME.io_diffCommits_info_25_rfWen = RTL_PATH.io_diffCommits_info_25_rfWen; \
        force U_IF_NAME.io_diffCommits_info_25_fpWen = RTL_PATH.io_diffCommits_info_25_fpWen; \
        force U_IF_NAME.io_diffCommits_info_25_vecWen = RTL_PATH.io_diffCommits_info_25_vecWen; \
        force U_IF_NAME.io_diffCommits_info_25_v0Wen = RTL_PATH.io_diffCommits_info_25_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_25_vlWen = RTL_PATH.io_diffCommits_info_25_vlWen; \
        force U_IF_NAME.io_diffCommits_info_26_ldest = RTL_PATH.io_diffCommits_info_26_ldest; \
        force U_IF_NAME.io_diffCommits_info_26_pdest = RTL_PATH.io_diffCommits_info_26_pdest; \
        force U_IF_NAME.io_diffCommits_info_26_rfWen = RTL_PATH.io_diffCommits_info_26_rfWen; \
        force U_IF_NAME.io_diffCommits_info_26_fpWen = RTL_PATH.io_diffCommits_info_26_fpWen; \
        force U_IF_NAME.io_diffCommits_info_26_vecWen = RTL_PATH.io_diffCommits_info_26_vecWen; \
        force U_IF_NAME.io_diffCommits_info_26_v0Wen = RTL_PATH.io_diffCommits_info_26_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_26_vlWen = RTL_PATH.io_diffCommits_info_26_vlWen; \
        force U_IF_NAME.io_diffCommits_info_27_ldest = RTL_PATH.io_diffCommits_info_27_ldest; \
        force U_IF_NAME.io_diffCommits_info_27_pdest = RTL_PATH.io_diffCommits_info_27_pdest; \
        force U_IF_NAME.io_diffCommits_info_27_rfWen = RTL_PATH.io_diffCommits_info_27_rfWen; \
        force U_IF_NAME.io_diffCommits_info_27_fpWen = RTL_PATH.io_diffCommits_info_27_fpWen; \
        force U_IF_NAME.io_diffCommits_info_27_vecWen = RTL_PATH.io_diffCommits_info_27_vecWen; \
        force U_IF_NAME.io_diffCommits_info_27_v0Wen = RTL_PATH.io_diffCommits_info_27_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_27_vlWen = RTL_PATH.io_diffCommits_info_27_vlWen; \
        force U_IF_NAME.io_diffCommits_info_28_ldest = RTL_PATH.io_diffCommits_info_28_ldest; \
        force U_IF_NAME.io_diffCommits_info_28_pdest = RTL_PATH.io_diffCommits_info_28_pdest; \
        force U_IF_NAME.io_diffCommits_info_28_rfWen = RTL_PATH.io_diffCommits_info_28_rfWen; \
        force U_IF_NAME.io_diffCommits_info_28_fpWen = RTL_PATH.io_diffCommits_info_28_fpWen; \
        force U_IF_NAME.io_diffCommits_info_28_vecWen = RTL_PATH.io_diffCommits_info_28_vecWen; \
        force U_IF_NAME.io_diffCommits_info_28_v0Wen = RTL_PATH.io_diffCommits_info_28_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_28_vlWen = RTL_PATH.io_diffCommits_info_28_vlWen; \
        force U_IF_NAME.io_diffCommits_info_29_ldest = RTL_PATH.io_diffCommits_info_29_ldest; \
        force U_IF_NAME.io_diffCommits_info_29_pdest = RTL_PATH.io_diffCommits_info_29_pdest; \
        force U_IF_NAME.io_diffCommits_info_29_rfWen = RTL_PATH.io_diffCommits_info_29_rfWen; \
        force U_IF_NAME.io_diffCommits_info_29_fpWen = RTL_PATH.io_diffCommits_info_29_fpWen; \
        force U_IF_NAME.io_diffCommits_info_29_vecWen = RTL_PATH.io_diffCommits_info_29_vecWen; \
        force U_IF_NAME.io_diffCommits_info_29_v0Wen = RTL_PATH.io_diffCommits_info_29_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_29_vlWen = RTL_PATH.io_diffCommits_info_29_vlWen; \
        force U_IF_NAME.io_diffCommits_info_30_ldest = RTL_PATH.io_diffCommits_info_30_ldest; \
        force U_IF_NAME.io_diffCommits_info_30_pdest = RTL_PATH.io_diffCommits_info_30_pdest; \
        force U_IF_NAME.io_diffCommits_info_30_rfWen = RTL_PATH.io_diffCommits_info_30_rfWen; \
        force U_IF_NAME.io_diffCommits_info_30_fpWen = RTL_PATH.io_diffCommits_info_30_fpWen; \
        force U_IF_NAME.io_diffCommits_info_30_vecWen = RTL_PATH.io_diffCommits_info_30_vecWen; \
        force U_IF_NAME.io_diffCommits_info_30_v0Wen = RTL_PATH.io_diffCommits_info_30_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_30_vlWen = RTL_PATH.io_diffCommits_info_30_vlWen; \
        force U_IF_NAME.io_diffCommits_info_31_ldest = RTL_PATH.io_diffCommits_info_31_ldest; \
        force U_IF_NAME.io_diffCommits_info_31_pdest = RTL_PATH.io_diffCommits_info_31_pdest; \
        force U_IF_NAME.io_diffCommits_info_31_rfWen = RTL_PATH.io_diffCommits_info_31_rfWen; \
        force U_IF_NAME.io_diffCommits_info_31_fpWen = RTL_PATH.io_diffCommits_info_31_fpWen; \
        force U_IF_NAME.io_diffCommits_info_31_vecWen = RTL_PATH.io_diffCommits_info_31_vecWen; \
        force U_IF_NAME.io_diffCommits_info_31_v0Wen = RTL_PATH.io_diffCommits_info_31_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_31_vlWen = RTL_PATH.io_diffCommits_info_31_vlWen; \
        force U_IF_NAME.io_diffCommits_info_32_ldest = RTL_PATH.io_diffCommits_info_32_ldest; \
        force U_IF_NAME.io_diffCommits_info_32_pdest = RTL_PATH.io_diffCommits_info_32_pdest; \
        force U_IF_NAME.io_diffCommits_info_32_rfWen = RTL_PATH.io_diffCommits_info_32_rfWen; \
        force U_IF_NAME.io_diffCommits_info_32_fpWen = RTL_PATH.io_diffCommits_info_32_fpWen; \
        force U_IF_NAME.io_diffCommits_info_32_vecWen = RTL_PATH.io_diffCommits_info_32_vecWen; \
        force U_IF_NAME.io_diffCommits_info_32_v0Wen = RTL_PATH.io_diffCommits_info_32_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_32_vlWen = RTL_PATH.io_diffCommits_info_32_vlWen; \
        force U_IF_NAME.io_diffCommits_info_33_ldest = RTL_PATH.io_diffCommits_info_33_ldest; \
        force U_IF_NAME.io_diffCommits_info_33_pdest = RTL_PATH.io_diffCommits_info_33_pdest; \
        force U_IF_NAME.io_diffCommits_info_33_rfWen = RTL_PATH.io_diffCommits_info_33_rfWen; \
        force U_IF_NAME.io_diffCommits_info_33_fpWen = RTL_PATH.io_diffCommits_info_33_fpWen; \
        force U_IF_NAME.io_diffCommits_info_33_vecWen = RTL_PATH.io_diffCommits_info_33_vecWen; \
        force U_IF_NAME.io_diffCommits_info_33_v0Wen = RTL_PATH.io_diffCommits_info_33_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_33_vlWen = RTL_PATH.io_diffCommits_info_33_vlWen; \
        force U_IF_NAME.io_diffCommits_info_34_ldest = RTL_PATH.io_diffCommits_info_34_ldest; \
        force U_IF_NAME.io_diffCommits_info_34_pdest = RTL_PATH.io_diffCommits_info_34_pdest; \
        force U_IF_NAME.io_diffCommits_info_34_rfWen = RTL_PATH.io_diffCommits_info_34_rfWen; \
        force U_IF_NAME.io_diffCommits_info_34_fpWen = RTL_PATH.io_diffCommits_info_34_fpWen; \
        force U_IF_NAME.io_diffCommits_info_34_vecWen = RTL_PATH.io_diffCommits_info_34_vecWen; \
        force U_IF_NAME.io_diffCommits_info_34_v0Wen = RTL_PATH.io_diffCommits_info_34_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_34_vlWen = RTL_PATH.io_diffCommits_info_34_vlWen; \
        force U_IF_NAME.io_diffCommits_info_35_ldest = RTL_PATH.io_diffCommits_info_35_ldest; \
        force U_IF_NAME.io_diffCommits_info_35_pdest = RTL_PATH.io_diffCommits_info_35_pdest; \
        force U_IF_NAME.io_diffCommits_info_35_rfWen = RTL_PATH.io_diffCommits_info_35_rfWen; \
        force U_IF_NAME.io_diffCommits_info_35_fpWen = RTL_PATH.io_diffCommits_info_35_fpWen; \
        force U_IF_NAME.io_diffCommits_info_35_vecWen = RTL_PATH.io_diffCommits_info_35_vecWen; \
        force U_IF_NAME.io_diffCommits_info_35_v0Wen = RTL_PATH.io_diffCommits_info_35_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_35_vlWen = RTL_PATH.io_diffCommits_info_35_vlWen; \
        force U_IF_NAME.io_diffCommits_info_36_ldest = RTL_PATH.io_diffCommits_info_36_ldest; \
        force U_IF_NAME.io_diffCommits_info_36_pdest = RTL_PATH.io_diffCommits_info_36_pdest; \
        force U_IF_NAME.io_diffCommits_info_36_rfWen = RTL_PATH.io_diffCommits_info_36_rfWen; \
        force U_IF_NAME.io_diffCommits_info_36_fpWen = RTL_PATH.io_diffCommits_info_36_fpWen; \
        force U_IF_NAME.io_diffCommits_info_36_vecWen = RTL_PATH.io_diffCommits_info_36_vecWen; \
        force U_IF_NAME.io_diffCommits_info_36_v0Wen = RTL_PATH.io_diffCommits_info_36_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_36_vlWen = RTL_PATH.io_diffCommits_info_36_vlWen; \
        force U_IF_NAME.io_diffCommits_info_37_ldest = RTL_PATH.io_diffCommits_info_37_ldest; \
        force U_IF_NAME.io_diffCommits_info_37_pdest = RTL_PATH.io_diffCommits_info_37_pdest; \
        force U_IF_NAME.io_diffCommits_info_37_rfWen = RTL_PATH.io_diffCommits_info_37_rfWen; \
        force U_IF_NAME.io_diffCommits_info_37_fpWen = RTL_PATH.io_diffCommits_info_37_fpWen; \
        force U_IF_NAME.io_diffCommits_info_37_vecWen = RTL_PATH.io_diffCommits_info_37_vecWen; \
        force U_IF_NAME.io_diffCommits_info_37_v0Wen = RTL_PATH.io_diffCommits_info_37_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_37_vlWen = RTL_PATH.io_diffCommits_info_37_vlWen; \
        force U_IF_NAME.io_diffCommits_info_38_ldest = RTL_PATH.io_diffCommits_info_38_ldest; \
        force U_IF_NAME.io_diffCommits_info_38_pdest = RTL_PATH.io_diffCommits_info_38_pdest; \
        force U_IF_NAME.io_diffCommits_info_38_rfWen = RTL_PATH.io_diffCommits_info_38_rfWen; \
        force U_IF_NAME.io_diffCommits_info_38_fpWen = RTL_PATH.io_diffCommits_info_38_fpWen; \
        force U_IF_NAME.io_diffCommits_info_38_vecWen = RTL_PATH.io_diffCommits_info_38_vecWen; \
        force U_IF_NAME.io_diffCommits_info_38_v0Wen = RTL_PATH.io_diffCommits_info_38_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_38_vlWen = RTL_PATH.io_diffCommits_info_38_vlWen; \
        force U_IF_NAME.io_diffCommits_info_39_ldest = RTL_PATH.io_diffCommits_info_39_ldest; \
        force U_IF_NAME.io_diffCommits_info_39_pdest = RTL_PATH.io_diffCommits_info_39_pdest; \
        force U_IF_NAME.io_diffCommits_info_39_rfWen = RTL_PATH.io_diffCommits_info_39_rfWen; \
        force U_IF_NAME.io_diffCommits_info_39_fpWen = RTL_PATH.io_diffCommits_info_39_fpWen; \
        force U_IF_NAME.io_diffCommits_info_39_vecWen = RTL_PATH.io_diffCommits_info_39_vecWen; \
        force U_IF_NAME.io_diffCommits_info_39_v0Wen = RTL_PATH.io_diffCommits_info_39_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_39_vlWen = RTL_PATH.io_diffCommits_info_39_vlWen; \
        force U_IF_NAME.io_diffCommits_info_40_ldest = RTL_PATH.io_diffCommits_info_40_ldest; \
        force U_IF_NAME.io_diffCommits_info_40_pdest = RTL_PATH.io_diffCommits_info_40_pdest; \
        force U_IF_NAME.io_diffCommits_info_40_rfWen = RTL_PATH.io_diffCommits_info_40_rfWen; \
        force U_IF_NAME.io_diffCommits_info_40_fpWen = RTL_PATH.io_diffCommits_info_40_fpWen; \
        force U_IF_NAME.io_diffCommits_info_40_vecWen = RTL_PATH.io_diffCommits_info_40_vecWen; \
        force U_IF_NAME.io_diffCommits_info_40_v0Wen = RTL_PATH.io_diffCommits_info_40_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_40_vlWen = RTL_PATH.io_diffCommits_info_40_vlWen; \
        force U_IF_NAME.io_diffCommits_info_41_ldest = RTL_PATH.io_diffCommits_info_41_ldest; \
        force U_IF_NAME.io_diffCommits_info_41_pdest = RTL_PATH.io_diffCommits_info_41_pdest; \
        force U_IF_NAME.io_diffCommits_info_41_rfWen = RTL_PATH.io_diffCommits_info_41_rfWen; \
        force U_IF_NAME.io_diffCommits_info_41_fpWen = RTL_PATH.io_diffCommits_info_41_fpWen; \
        force U_IF_NAME.io_diffCommits_info_41_vecWen = RTL_PATH.io_diffCommits_info_41_vecWen; \
        force U_IF_NAME.io_diffCommits_info_41_v0Wen = RTL_PATH.io_diffCommits_info_41_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_41_vlWen = RTL_PATH.io_diffCommits_info_41_vlWen; \
        force U_IF_NAME.io_diffCommits_info_42_ldest = RTL_PATH.io_diffCommits_info_42_ldest; \
        force U_IF_NAME.io_diffCommits_info_42_pdest = RTL_PATH.io_diffCommits_info_42_pdest; \
        force U_IF_NAME.io_diffCommits_info_42_rfWen = RTL_PATH.io_diffCommits_info_42_rfWen; \
        force U_IF_NAME.io_diffCommits_info_42_fpWen = RTL_PATH.io_diffCommits_info_42_fpWen; \
        force U_IF_NAME.io_diffCommits_info_42_vecWen = RTL_PATH.io_diffCommits_info_42_vecWen; \
        force U_IF_NAME.io_diffCommits_info_42_v0Wen = RTL_PATH.io_diffCommits_info_42_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_42_vlWen = RTL_PATH.io_diffCommits_info_42_vlWen; \
        force U_IF_NAME.io_diffCommits_info_43_ldest = RTL_PATH.io_diffCommits_info_43_ldest; \
        force U_IF_NAME.io_diffCommits_info_43_pdest = RTL_PATH.io_diffCommits_info_43_pdest; \
        force U_IF_NAME.io_diffCommits_info_43_rfWen = RTL_PATH.io_diffCommits_info_43_rfWen; \
        force U_IF_NAME.io_diffCommits_info_43_fpWen = RTL_PATH.io_diffCommits_info_43_fpWen; \
        force U_IF_NAME.io_diffCommits_info_43_vecWen = RTL_PATH.io_diffCommits_info_43_vecWen; \
        force U_IF_NAME.io_diffCommits_info_43_v0Wen = RTL_PATH.io_diffCommits_info_43_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_43_vlWen = RTL_PATH.io_diffCommits_info_43_vlWen; \
        force U_IF_NAME.io_diffCommits_info_44_ldest = RTL_PATH.io_diffCommits_info_44_ldest; \
        force U_IF_NAME.io_diffCommits_info_44_pdest = RTL_PATH.io_diffCommits_info_44_pdest; \
        force U_IF_NAME.io_diffCommits_info_44_rfWen = RTL_PATH.io_diffCommits_info_44_rfWen; \
        force U_IF_NAME.io_diffCommits_info_44_fpWen = RTL_PATH.io_diffCommits_info_44_fpWen; \
        force U_IF_NAME.io_diffCommits_info_44_vecWen = RTL_PATH.io_diffCommits_info_44_vecWen; \
        force U_IF_NAME.io_diffCommits_info_44_v0Wen = RTL_PATH.io_diffCommits_info_44_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_44_vlWen = RTL_PATH.io_diffCommits_info_44_vlWen; \
        force U_IF_NAME.io_diffCommits_info_45_ldest = RTL_PATH.io_diffCommits_info_45_ldest; \
        force U_IF_NAME.io_diffCommits_info_45_pdest = RTL_PATH.io_diffCommits_info_45_pdest; \
        force U_IF_NAME.io_diffCommits_info_45_rfWen = RTL_PATH.io_diffCommits_info_45_rfWen; \
        force U_IF_NAME.io_diffCommits_info_45_fpWen = RTL_PATH.io_diffCommits_info_45_fpWen; \
        force U_IF_NAME.io_diffCommits_info_45_vecWen = RTL_PATH.io_diffCommits_info_45_vecWen; \
        force U_IF_NAME.io_diffCommits_info_45_v0Wen = RTL_PATH.io_diffCommits_info_45_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_45_vlWen = RTL_PATH.io_diffCommits_info_45_vlWen; \
        force U_IF_NAME.io_diffCommits_info_46_ldest = RTL_PATH.io_diffCommits_info_46_ldest; \
        force U_IF_NAME.io_diffCommits_info_46_pdest = RTL_PATH.io_diffCommits_info_46_pdest; \
        force U_IF_NAME.io_diffCommits_info_46_rfWen = RTL_PATH.io_diffCommits_info_46_rfWen; \
        force U_IF_NAME.io_diffCommits_info_46_fpWen = RTL_PATH.io_diffCommits_info_46_fpWen; \
        force U_IF_NAME.io_diffCommits_info_46_vecWen = RTL_PATH.io_diffCommits_info_46_vecWen; \
        force U_IF_NAME.io_diffCommits_info_46_v0Wen = RTL_PATH.io_diffCommits_info_46_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_46_vlWen = RTL_PATH.io_diffCommits_info_46_vlWen; \
        force U_IF_NAME.io_diffCommits_info_47_ldest = RTL_PATH.io_diffCommits_info_47_ldest; \
        force U_IF_NAME.io_diffCommits_info_47_pdest = RTL_PATH.io_diffCommits_info_47_pdest; \
        force U_IF_NAME.io_diffCommits_info_47_rfWen = RTL_PATH.io_diffCommits_info_47_rfWen; \
        force U_IF_NAME.io_diffCommits_info_47_fpWen = RTL_PATH.io_diffCommits_info_47_fpWen; \
        force U_IF_NAME.io_diffCommits_info_47_vecWen = RTL_PATH.io_diffCommits_info_47_vecWen; \
        force U_IF_NAME.io_diffCommits_info_47_v0Wen = RTL_PATH.io_diffCommits_info_47_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_47_vlWen = RTL_PATH.io_diffCommits_info_47_vlWen; \
        force U_IF_NAME.io_diffCommits_info_48_ldest = RTL_PATH.io_diffCommits_info_48_ldest; \
        force U_IF_NAME.io_diffCommits_info_48_pdest = RTL_PATH.io_diffCommits_info_48_pdest; \
        force U_IF_NAME.io_diffCommits_info_48_rfWen = RTL_PATH.io_diffCommits_info_48_rfWen; \
        force U_IF_NAME.io_diffCommits_info_48_fpWen = RTL_PATH.io_diffCommits_info_48_fpWen; \
        force U_IF_NAME.io_diffCommits_info_48_vecWen = RTL_PATH.io_diffCommits_info_48_vecWen; \
        force U_IF_NAME.io_diffCommits_info_48_v0Wen = RTL_PATH.io_diffCommits_info_48_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_48_vlWen = RTL_PATH.io_diffCommits_info_48_vlWen; \
        force U_IF_NAME.io_diffCommits_info_49_ldest = RTL_PATH.io_diffCommits_info_49_ldest; \
        force U_IF_NAME.io_diffCommits_info_49_pdest = RTL_PATH.io_diffCommits_info_49_pdest; \
        force U_IF_NAME.io_diffCommits_info_49_rfWen = RTL_PATH.io_diffCommits_info_49_rfWen; \
        force U_IF_NAME.io_diffCommits_info_49_fpWen = RTL_PATH.io_diffCommits_info_49_fpWen; \
        force U_IF_NAME.io_diffCommits_info_49_vecWen = RTL_PATH.io_diffCommits_info_49_vecWen; \
        force U_IF_NAME.io_diffCommits_info_49_v0Wen = RTL_PATH.io_diffCommits_info_49_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_49_vlWen = RTL_PATH.io_diffCommits_info_49_vlWen; \
        force U_IF_NAME.io_diffCommits_info_50_ldest = RTL_PATH.io_diffCommits_info_50_ldest; \
        force U_IF_NAME.io_diffCommits_info_50_pdest = RTL_PATH.io_diffCommits_info_50_pdest; \
        force U_IF_NAME.io_diffCommits_info_50_rfWen = RTL_PATH.io_diffCommits_info_50_rfWen; \
        force U_IF_NAME.io_diffCommits_info_50_fpWen = RTL_PATH.io_diffCommits_info_50_fpWen; \
        force U_IF_NAME.io_diffCommits_info_50_vecWen = RTL_PATH.io_diffCommits_info_50_vecWen; \
        force U_IF_NAME.io_diffCommits_info_50_v0Wen = RTL_PATH.io_diffCommits_info_50_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_50_vlWen = RTL_PATH.io_diffCommits_info_50_vlWen; \
        force U_IF_NAME.io_diffCommits_info_51_ldest = RTL_PATH.io_diffCommits_info_51_ldest; \
        force U_IF_NAME.io_diffCommits_info_51_pdest = RTL_PATH.io_diffCommits_info_51_pdest; \
        force U_IF_NAME.io_diffCommits_info_51_rfWen = RTL_PATH.io_diffCommits_info_51_rfWen; \
        force U_IF_NAME.io_diffCommits_info_51_fpWen = RTL_PATH.io_diffCommits_info_51_fpWen; \
        force U_IF_NAME.io_diffCommits_info_51_vecWen = RTL_PATH.io_diffCommits_info_51_vecWen; \
        force U_IF_NAME.io_diffCommits_info_51_v0Wen = RTL_PATH.io_diffCommits_info_51_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_51_vlWen = RTL_PATH.io_diffCommits_info_51_vlWen; \
        force U_IF_NAME.io_diffCommits_info_52_ldest = RTL_PATH.io_diffCommits_info_52_ldest; \
        force U_IF_NAME.io_diffCommits_info_52_pdest = RTL_PATH.io_diffCommits_info_52_pdest; \
        force U_IF_NAME.io_diffCommits_info_52_rfWen = RTL_PATH.io_diffCommits_info_52_rfWen; \
        force U_IF_NAME.io_diffCommits_info_52_fpWen = RTL_PATH.io_diffCommits_info_52_fpWen; \
        force U_IF_NAME.io_diffCommits_info_52_vecWen = RTL_PATH.io_diffCommits_info_52_vecWen; \
        force U_IF_NAME.io_diffCommits_info_52_v0Wen = RTL_PATH.io_diffCommits_info_52_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_52_vlWen = RTL_PATH.io_diffCommits_info_52_vlWen; \
        force U_IF_NAME.io_diffCommits_info_53_ldest = RTL_PATH.io_diffCommits_info_53_ldest; \
        force U_IF_NAME.io_diffCommits_info_53_pdest = RTL_PATH.io_diffCommits_info_53_pdest; \
        force U_IF_NAME.io_diffCommits_info_53_rfWen = RTL_PATH.io_diffCommits_info_53_rfWen; \
        force U_IF_NAME.io_diffCommits_info_53_fpWen = RTL_PATH.io_diffCommits_info_53_fpWen; \
        force U_IF_NAME.io_diffCommits_info_53_vecWen = RTL_PATH.io_diffCommits_info_53_vecWen; \
        force U_IF_NAME.io_diffCommits_info_53_v0Wen = RTL_PATH.io_diffCommits_info_53_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_53_vlWen = RTL_PATH.io_diffCommits_info_53_vlWen; \
        force U_IF_NAME.io_diffCommits_info_54_ldest = RTL_PATH.io_diffCommits_info_54_ldest; \
        force U_IF_NAME.io_diffCommits_info_54_pdest = RTL_PATH.io_diffCommits_info_54_pdest; \
        force U_IF_NAME.io_diffCommits_info_54_rfWen = RTL_PATH.io_diffCommits_info_54_rfWen; \
        force U_IF_NAME.io_diffCommits_info_54_fpWen = RTL_PATH.io_diffCommits_info_54_fpWen; \
        force U_IF_NAME.io_diffCommits_info_54_vecWen = RTL_PATH.io_diffCommits_info_54_vecWen; \
        force U_IF_NAME.io_diffCommits_info_54_v0Wen = RTL_PATH.io_diffCommits_info_54_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_54_vlWen = RTL_PATH.io_diffCommits_info_54_vlWen; \
        force U_IF_NAME.io_diffCommits_info_55_ldest = RTL_PATH.io_diffCommits_info_55_ldest; \
        force U_IF_NAME.io_diffCommits_info_55_pdest = RTL_PATH.io_diffCommits_info_55_pdest; \
        force U_IF_NAME.io_diffCommits_info_55_rfWen = RTL_PATH.io_diffCommits_info_55_rfWen; \
        force U_IF_NAME.io_diffCommits_info_55_fpWen = RTL_PATH.io_diffCommits_info_55_fpWen; \
        force U_IF_NAME.io_diffCommits_info_55_vecWen = RTL_PATH.io_diffCommits_info_55_vecWen; \
        force U_IF_NAME.io_diffCommits_info_55_v0Wen = RTL_PATH.io_diffCommits_info_55_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_55_vlWen = RTL_PATH.io_diffCommits_info_55_vlWen; \
        force U_IF_NAME.io_diffCommits_info_56_ldest = RTL_PATH.io_diffCommits_info_56_ldest; \
        force U_IF_NAME.io_diffCommits_info_56_pdest = RTL_PATH.io_diffCommits_info_56_pdest; \
        force U_IF_NAME.io_diffCommits_info_56_rfWen = RTL_PATH.io_diffCommits_info_56_rfWen; \
        force U_IF_NAME.io_diffCommits_info_56_fpWen = RTL_PATH.io_diffCommits_info_56_fpWen; \
        force U_IF_NAME.io_diffCommits_info_56_vecWen = RTL_PATH.io_diffCommits_info_56_vecWen; \
        force U_IF_NAME.io_diffCommits_info_56_v0Wen = RTL_PATH.io_diffCommits_info_56_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_56_vlWen = RTL_PATH.io_diffCommits_info_56_vlWen; \
        force U_IF_NAME.io_diffCommits_info_57_ldest = RTL_PATH.io_diffCommits_info_57_ldest; \
        force U_IF_NAME.io_diffCommits_info_57_pdest = RTL_PATH.io_diffCommits_info_57_pdest; \
        force U_IF_NAME.io_diffCommits_info_57_rfWen = RTL_PATH.io_diffCommits_info_57_rfWen; \
        force U_IF_NAME.io_diffCommits_info_57_fpWen = RTL_PATH.io_diffCommits_info_57_fpWen; \
        force U_IF_NAME.io_diffCommits_info_57_vecWen = RTL_PATH.io_diffCommits_info_57_vecWen; \
        force U_IF_NAME.io_diffCommits_info_57_v0Wen = RTL_PATH.io_diffCommits_info_57_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_57_vlWen = RTL_PATH.io_diffCommits_info_57_vlWen; \
        force U_IF_NAME.io_diffCommits_info_58_ldest = RTL_PATH.io_diffCommits_info_58_ldest; \
        force U_IF_NAME.io_diffCommits_info_58_pdest = RTL_PATH.io_diffCommits_info_58_pdest; \
        force U_IF_NAME.io_diffCommits_info_58_rfWen = RTL_PATH.io_diffCommits_info_58_rfWen; \
        force U_IF_NAME.io_diffCommits_info_58_fpWen = RTL_PATH.io_diffCommits_info_58_fpWen; \
        force U_IF_NAME.io_diffCommits_info_58_vecWen = RTL_PATH.io_diffCommits_info_58_vecWen; \
        force U_IF_NAME.io_diffCommits_info_58_v0Wen = RTL_PATH.io_diffCommits_info_58_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_58_vlWen = RTL_PATH.io_diffCommits_info_58_vlWen; \
        force U_IF_NAME.io_diffCommits_info_59_ldest = RTL_PATH.io_diffCommits_info_59_ldest; \
        force U_IF_NAME.io_diffCommits_info_59_pdest = RTL_PATH.io_diffCommits_info_59_pdest; \
        force U_IF_NAME.io_diffCommits_info_59_rfWen = RTL_PATH.io_diffCommits_info_59_rfWen; \
        force U_IF_NAME.io_diffCommits_info_59_fpWen = RTL_PATH.io_diffCommits_info_59_fpWen; \
        force U_IF_NAME.io_diffCommits_info_59_vecWen = RTL_PATH.io_diffCommits_info_59_vecWen; \
        force U_IF_NAME.io_diffCommits_info_59_v0Wen = RTL_PATH.io_diffCommits_info_59_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_59_vlWen = RTL_PATH.io_diffCommits_info_59_vlWen; \
        force U_IF_NAME.io_diffCommits_info_60_ldest = RTL_PATH.io_diffCommits_info_60_ldest; \
        force U_IF_NAME.io_diffCommits_info_60_pdest = RTL_PATH.io_diffCommits_info_60_pdest; \
        force U_IF_NAME.io_diffCommits_info_60_rfWen = RTL_PATH.io_diffCommits_info_60_rfWen; \
        force U_IF_NAME.io_diffCommits_info_60_fpWen = RTL_PATH.io_diffCommits_info_60_fpWen; \
        force U_IF_NAME.io_diffCommits_info_60_vecWen = RTL_PATH.io_diffCommits_info_60_vecWen; \
        force U_IF_NAME.io_diffCommits_info_60_v0Wen = RTL_PATH.io_diffCommits_info_60_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_60_vlWen = RTL_PATH.io_diffCommits_info_60_vlWen; \
        force U_IF_NAME.io_diffCommits_info_61_ldest = RTL_PATH.io_diffCommits_info_61_ldest; \
        force U_IF_NAME.io_diffCommits_info_61_pdest = RTL_PATH.io_diffCommits_info_61_pdest; \
        force U_IF_NAME.io_diffCommits_info_61_rfWen = RTL_PATH.io_diffCommits_info_61_rfWen; \
        force U_IF_NAME.io_diffCommits_info_61_fpWen = RTL_PATH.io_diffCommits_info_61_fpWen; \
        force U_IF_NAME.io_diffCommits_info_61_vecWen = RTL_PATH.io_diffCommits_info_61_vecWen; \
        force U_IF_NAME.io_diffCommits_info_61_v0Wen = RTL_PATH.io_diffCommits_info_61_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_61_vlWen = RTL_PATH.io_diffCommits_info_61_vlWen; \
        force U_IF_NAME.io_diffCommits_info_62_ldest = RTL_PATH.io_diffCommits_info_62_ldest; \
        force U_IF_NAME.io_diffCommits_info_62_pdest = RTL_PATH.io_diffCommits_info_62_pdest; \
        force U_IF_NAME.io_diffCommits_info_62_rfWen = RTL_PATH.io_diffCommits_info_62_rfWen; \
        force U_IF_NAME.io_diffCommits_info_62_fpWen = RTL_PATH.io_diffCommits_info_62_fpWen; \
        force U_IF_NAME.io_diffCommits_info_62_vecWen = RTL_PATH.io_diffCommits_info_62_vecWen; \
        force U_IF_NAME.io_diffCommits_info_62_v0Wen = RTL_PATH.io_diffCommits_info_62_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_62_vlWen = RTL_PATH.io_diffCommits_info_62_vlWen; \
        force U_IF_NAME.io_diffCommits_info_63_ldest = RTL_PATH.io_diffCommits_info_63_ldest; \
        force U_IF_NAME.io_diffCommits_info_63_pdest = RTL_PATH.io_diffCommits_info_63_pdest; \
        force U_IF_NAME.io_diffCommits_info_63_rfWen = RTL_PATH.io_diffCommits_info_63_rfWen; \
        force U_IF_NAME.io_diffCommits_info_63_fpWen = RTL_PATH.io_diffCommits_info_63_fpWen; \
        force U_IF_NAME.io_diffCommits_info_63_vecWen = RTL_PATH.io_diffCommits_info_63_vecWen; \
        force U_IF_NAME.io_diffCommits_info_63_v0Wen = RTL_PATH.io_diffCommits_info_63_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_63_vlWen = RTL_PATH.io_diffCommits_info_63_vlWen; \
        force U_IF_NAME.io_diffCommits_info_64_ldest = RTL_PATH.io_diffCommits_info_64_ldest; \
        force U_IF_NAME.io_diffCommits_info_64_pdest = RTL_PATH.io_diffCommits_info_64_pdest; \
        force U_IF_NAME.io_diffCommits_info_64_rfWen = RTL_PATH.io_diffCommits_info_64_rfWen; \
        force U_IF_NAME.io_diffCommits_info_64_fpWen = RTL_PATH.io_diffCommits_info_64_fpWen; \
        force U_IF_NAME.io_diffCommits_info_64_vecWen = RTL_PATH.io_diffCommits_info_64_vecWen; \
        force U_IF_NAME.io_diffCommits_info_64_v0Wen = RTL_PATH.io_diffCommits_info_64_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_64_vlWen = RTL_PATH.io_diffCommits_info_64_vlWen; \
        force U_IF_NAME.io_diffCommits_info_65_ldest = RTL_PATH.io_diffCommits_info_65_ldest; \
        force U_IF_NAME.io_diffCommits_info_65_pdest = RTL_PATH.io_diffCommits_info_65_pdest; \
        force U_IF_NAME.io_diffCommits_info_65_rfWen = RTL_PATH.io_diffCommits_info_65_rfWen; \
        force U_IF_NAME.io_diffCommits_info_65_fpWen = RTL_PATH.io_diffCommits_info_65_fpWen; \
        force U_IF_NAME.io_diffCommits_info_65_vecWen = RTL_PATH.io_diffCommits_info_65_vecWen; \
        force U_IF_NAME.io_diffCommits_info_65_v0Wen = RTL_PATH.io_diffCommits_info_65_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_65_vlWen = RTL_PATH.io_diffCommits_info_65_vlWen; \
        force U_IF_NAME.io_diffCommits_info_66_ldest = RTL_PATH.io_diffCommits_info_66_ldest; \
        force U_IF_NAME.io_diffCommits_info_66_pdest = RTL_PATH.io_diffCommits_info_66_pdest; \
        force U_IF_NAME.io_diffCommits_info_66_rfWen = RTL_PATH.io_diffCommits_info_66_rfWen; \
        force U_IF_NAME.io_diffCommits_info_66_fpWen = RTL_PATH.io_diffCommits_info_66_fpWen; \
        force U_IF_NAME.io_diffCommits_info_66_vecWen = RTL_PATH.io_diffCommits_info_66_vecWen; \
        force U_IF_NAME.io_diffCommits_info_66_v0Wen = RTL_PATH.io_diffCommits_info_66_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_66_vlWen = RTL_PATH.io_diffCommits_info_66_vlWen; \
        force U_IF_NAME.io_diffCommits_info_67_ldest = RTL_PATH.io_diffCommits_info_67_ldest; \
        force U_IF_NAME.io_diffCommits_info_67_pdest = RTL_PATH.io_diffCommits_info_67_pdest; \
        force U_IF_NAME.io_diffCommits_info_67_rfWen = RTL_PATH.io_diffCommits_info_67_rfWen; \
        force U_IF_NAME.io_diffCommits_info_67_fpWen = RTL_PATH.io_diffCommits_info_67_fpWen; \
        force U_IF_NAME.io_diffCommits_info_67_vecWen = RTL_PATH.io_diffCommits_info_67_vecWen; \
        force U_IF_NAME.io_diffCommits_info_67_v0Wen = RTL_PATH.io_diffCommits_info_67_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_67_vlWen = RTL_PATH.io_diffCommits_info_67_vlWen; \
        force U_IF_NAME.io_diffCommits_info_68_ldest = RTL_PATH.io_diffCommits_info_68_ldest; \
        force U_IF_NAME.io_diffCommits_info_68_pdest = RTL_PATH.io_diffCommits_info_68_pdest; \
        force U_IF_NAME.io_diffCommits_info_68_rfWen = RTL_PATH.io_diffCommits_info_68_rfWen; \
        force U_IF_NAME.io_diffCommits_info_68_fpWen = RTL_PATH.io_diffCommits_info_68_fpWen; \
        force U_IF_NAME.io_diffCommits_info_68_vecWen = RTL_PATH.io_diffCommits_info_68_vecWen; \
        force U_IF_NAME.io_diffCommits_info_68_v0Wen = RTL_PATH.io_diffCommits_info_68_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_68_vlWen = RTL_PATH.io_diffCommits_info_68_vlWen; \
        force U_IF_NAME.io_diffCommits_info_69_ldest = RTL_PATH.io_diffCommits_info_69_ldest; \
        force U_IF_NAME.io_diffCommits_info_69_pdest = RTL_PATH.io_diffCommits_info_69_pdest; \
        force U_IF_NAME.io_diffCommits_info_69_rfWen = RTL_PATH.io_diffCommits_info_69_rfWen; \
        force U_IF_NAME.io_diffCommits_info_69_fpWen = RTL_PATH.io_diffCommits_info_69_fpWen; \
        force U_IF_NAME.io_diffCommits_info_69_vecWen = RTL_PATH.io_diffCommits_info_69_vecWen; \
        force U_IF_NAME.io_diffCommits_info_69_v0Wen = RTL_PATH.io_diffCommits_info_69_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_69_vlWen = RTL_PATH.io_diffCommits_info_69_vlWen; \
        force U_IF_NAME.io_diffCommits_info_70_ldest = RTL_PATH.io_diffCommits_info_70_ldest; \
        force U_IF_NAME.io_diffCommits_info_70_pdest = RTL_PATH.io_diffCommits_info_70_pdest; \
        force U_IF_NAME.io_diffCommits_info_70_rfWen = RTL_PATH.io_diffCommits_info_70_rfWen; \
        force U_IF_NAME.io_diffCommits_info_70_fpWen = RTL_PATH.io_diffCommits_info_70_fpWen; \
        force U_IF_NAME.io_diffCommits_info_70_vecWen = RTL_PATH.io_diffCommits_info_70_vecWen; \
        force U_IF_NAME.io_diffCommits_info_70_v0Wen = RTL_PATH.io_diffCommits_info_70_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_70_vlWen = RTL_PATH.io_diffCommits_info_70_vlWen; \
        force U_IF_NAME.io_diffCommits_info_71_ldest = RTL_PATH.io_diffCommits_info_71_ldest; \
        force U_IF_NAME.io_diffCommits_info_71_pdest = RTL_PATH.io_diffCommits_info_71_pdest; \
        force U_IF_NAME.io_diffCommits_info_71_rfWen = RTL_PATH.io_diffCommits_info_71_rfWen; \
        force U_IF_NAME.io_diffCommits_info_71_fpWen = RTL_PATH.io_diffCommits_info_71_fpWen; \
        force U_IF_NAME.io_diffCommits_info_71_vecWen = RTL_PATH.io_diffCommits_info_71_vecWen; \
        force U_IF_NAME.io_diffCommits_info_71_v0Wen = RTL_PATH.io_diffCommits_info_71_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_71_vlWen = RTL_PATH.io_diffCommits_info_71_vlWen; \
        force U_IF_NAME.io_diffCommits_info_72_ldest = RTL_PATH.io_diffCommits_info_72_ldest; \
        force U_IF_NAME.io_diffCommits_info_72_pdest = RTL_PATH.io_diffCommits_info_72_pdest; \
        force U_IF_NAME.io_diffCommits_info_72_rfWen = RTL_PATH.io_diffCommits_info_72_rfWen; \
        force U_IF_NAME.io_diffCommits_info_72_fpWen = RTL_PATH.io_diffCommits_info_72_fpWen; \
        force U_IF_NAME.io_diffCommits_info_72_vecWen = RTL_PATH.io_diffCommits_info_72_vecWen; \
        force U_IF_NAME.io_diffCommits_info_72_v0Wen = RTL_PATH.io_diffCommits_info_72_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_72_vlWen = RTL_PATH.io_diffCommits_info_72_vlWen; \
        force U_IF_NAME.io_diffCommits_info_73_ldest = RTL_PATH.io_diffCommits_info_73_ldest; \
        force U_IF_NAME.io_diffCommits_info_73_pdest = RTL_PATH.io_diffCommits_info_73_pdest; \
        force U_IF_NAME.io_diffCommits_info_73_rfWen = RTL_PATH.io_diffCommits_info_73_rfWen; \
        force U_IF_NAME.io_diffCommits_info_73_fpWen = RTL_PATH.io_diffCommits_info_73_fpWen; \
        force U_IF_NAME.io_diffCommits_info_73_vecWen = RTL_PATH.io_diffCommits_info_73_vecWen; \
        force U_IF_NAME.io_diffCommits_info_73_v0Wen = RTL_PATH.io_diffCommits_info_73_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_73_vlWen = RTL_PATH.io_diffCommits_info_73_vlWen; \
        force U_IF_NAME.io_diffCommits_info_74_ldest = RTL_PATH.io_diffCommits_info_74_ldest; \
        force U_IF_NAME.io_diffCommits_info_74_pdest = RTL_PATH.io_diffCommits_info_74_pdest; \
        force U_IF_NAME.io_diffCommits_info_74_rfWen = RTL_PATH.io_diffCommits_info_74_rfWen; \
        force U_IF_NAME.io_diffCommits_info_74_fpWen = RTL_PATH.io_diffCommits_info_74_fpWen; \
        force U_IF_NAME.io_diffCommits_info_74_vecWen = RTL_PATH.io_diffCommits_info_74_vecWen; \
        force U_IF_NAME.io_diffCommits_info_74_v0Wen = RTL_PATH.io_diffCommits_info_74_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_74_vlWen = RTL_PATH.io_diffCommits_info_74_vlWen; \
        force U_IF_NAME.io_diffCommits_info_75_ldest = RTL_PATH.io_diffCommits_info_75_ldest; \
        force U_IF_NAME.io_diffCommits_info_75_pdest = RTL_PATH.io_diffCommits_info_75_pdest; \
        force U_IF_NAME.io_diffCommits_info_75_rfWen = RTL_PATH.io_diffCommits_info_75_rfWen; \
        force U_IF_NAME.io_diffCommits_info_75_fpWen = RTL_PATH.io_diffCommits_info_75_fpWen; \
        force U_IF_NAME.io_diffCommits_info_75_vecWen = RTL_PATH.io_diffCommits_info_75_vecWen; \
        force U_IF_NAME.io_diffCommits_info_75_v0Wen = RTL_PATH.io_diffCommits_info_75_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_75_vlWen = RTL_PATH.io_diffCommits_info_75_vlWen; \
        force U_IF_NAME.io_diffCommits_info_76_ldest = RTL_PATH.io_diffCommits_info_76_ldest; \
        force U_IF_NAME.io_diffCommits_info_76_pdest = RTL_PATH.io_diffCommits_info_76_pdest; \
        force U_IF_NAME.io_diffCommits_info_76_rfWen = RTL_PATH.io_diffCommits_info_76_rfWen; \
        force U_IF_NAME.io_diffCommits_info_76_fpWen = RTL_PATH.io_diffCommits_info_76_fpWen; \
        force U_IF_NAME.io_diffCommits_info_76_vecWen = RTL_PATH.io_diffCommits_info_76_vecWen; \
        force U_IF_NAME.io_diffCommits_info_76_v0Wen = RTL_PATH.io_diffCommits_info_76_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_76_vlWen = RTL_PATH.io_diffCommits_info_76_vlWen; \
        force U_IF_NAME.io_diffCommits_info_77_ldest = RTL_PATH.io_diffCommits_info_77_ldest; \
        force U_IF_NAME.io_diffCommits_info_77_pdest = RTL_PATH.io_diffCommits_info_77_pdest; \
        force U_IF_NAME.io_diffCommits_info_77_rfWen = RTL_PATH.io_diffCommits_info_77_rfWen; \
        force U_IF_NAME.io_diffCommits_info_77_fpWen = RTL_PATH.io_diffCommits_info_77_fpWen; \
        force U_IF_NAME.io_diffCommits_info_77_vecWen = RTL_PATH.io_diffCommits_info_77_vecWen; \
        force U_IF_NAME.io_diffCommits_info_77_v0Wen = RTL_PATH.io_diffCommits_info_77_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_77_vlWen = RTL_PATH.io_diffCommits_info_77_vlWen; \
        force U_IF_NAME.io_diffCommits_info_78_ldest = RTL_PATH.io_diffCommits_info_78_ldest; \
        force U_IF_NAME.io_diffCommits_info_78_pdest = RTL_PATH.io_diffCommits_info_78_pdest; \
        force U_IF_NAME.io_diffCommits_info_78_rfWen = RTL_PATH.io_diffCommits_info_78_rfWen; \
        force U_IF_NAME.io_diffCommits_info_78_fpWen = RTL_PATH.io_diffCommits_info_78_fpWen; \
        force U_IF_NAME.io_diffCommits_info_78_vecWen = RTL_PATH.io_diffCommits_info_78_vecWen; \
        force U_IF_NAME.io_diffCommits_info_78_v0Wen = RTL_PATH.io_diffCommits_info_78_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_78_vlWen = RTL_PATH.io_diffCommits_info_78_vlWen; \
        force U_IF_NAME.io_diffCommits_info_79_ldest = RTL_PATH.io_diffCommits_info_79_ldest; \
        force U_IF_NAME.io_diffCommits_info_79_pdest = RTL_PATH.io_diffCommits_info_79_pdest; \
        force U_IF_NAME.io_diffCommits_info_79_rfWen = RTL_PATH.io_diffCommits_info_79_rfWen; \
        force U_IF_NAME.io_diffCommits_info_79_fpWen = RTL_PATH.io_diffCommits_info_79_fpWen; \
        force U_IF_NAME.io_diffCommits_info_79_vecWen = RTL_PATH.io_diffCommits_info_79_vecWen; \
        force U_IF_NAME.io_diffCommits_info_79_v0Wen = RTL_PATH.io_diffCommits_info_79_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_79_vlWen = RTL_PATH.io_diffCommits_info_79_vlWen; \
        force U_IF_NAME.io_diffCommits_info_80_ldest = RTL_PATH.io_diffCommits_info_80_ldest; \
        force U_IF_NAME.io_diffCommits_info_80_pdest = RTL_PATH.io_diffCommits_info_80_pdest; \
        force U_IF_NAME.io_diffCommits_info_80_rfWen = RTL_PATH.io_diffCommits_info_80_rfWen; \
        force U_IF_NAME.io_diffCommits_info_80_fpWen = RTL_PATH.io_diffCommits_info_80_fpWen; \
        force U_IF_NAME.io_diffCommits_info_80_vecWen = RTL_PATH.io_diffCommits_info_80_vecWen; \
        force U_IF_NAME.io_diffCommits_info_80_v0Wen = RTL_PATH.io_diffCommits_info_80_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_80_vlWen = RTL_PATH.io_diffCommits_info_80_vlWen; \
        force U_IF_NAME.io_diffCommits_info_81_ldest = RTL_PATH.io_diffCommits_info_81_ldest; \
        force U_IF_NAME.io_diffCommits_info_81_pdest = RTL_PATH.io_diffCommits_info_81_pdest; \
        force U_IF_NAME.io_diffCommits_info_81_rfWen = RTL_PATH.io_diffCommits_info_81_rfWen; \
        force U_IF_NAME.io_diffCommits_info_81_fpWen = RTL_PATH.io_diffCommits_info_81_fpWen; \
        force U_IF_NAME.io_diffCommits_info_81_vecWen = RTL_PATH.io_diffCommits_info_81_vecWen; \
        force U_IF_NAME.io_diffCommits_info_81_v0Wen = RTL_PATH.io_diffCommits_info_81_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_81_vlWen = RTL_PATH.io_diffCommits_info_81_vlWen; \
        force U_IF_NAME.io_diffCommits_info_82_ldest = RTL_PATH.io_diffCommits_info_82_ldest; \
        force U_IF_NAME.io_diffCommits_info_82_pdest = RTL_PATH.io_diffCommits_info_82_pdest; \
        force U_IF_NAME.io_diffCommits_info_82_rfWen = RTL_PATH.io_diffCommits_info_82_rfWen; \
        force U_IF_NAME.io_diffCommits_info_82_fpWen = RTL_PATH.io_diffCommits_info_82_fpWen; \
        force U_IF_NAME.io_diffCommits_info_82_vecWen = RTL_PATH.io_diffCommits_info_82_vecWen; \
        force U_IF_NAME.io_diffCommits_info_82_v0Wen = RTL_PATH.io_diffCommits_info_82_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_82_vlWen = RTL_PATH.io_diffCommits_info_82_vlWen; \
        force U_IF_NAME.io_diffCommits_info_83_ldest = RTL_PATH.io_diffCommits_info_83_ldest; \
        force U_IF_NAME.io_diffCommits_info_83_pdest = RTL_PATH.io_diffCommits_info_83_pdest; \
        force U_IF_NAME.io_diffCommits_info_83_rfWen = RTL_PATH.io_diffCommits_info_83_rfWen; \
        force U_IF_NAME.io_diffCommits_info_83_fpWen = RTL_PATH.io_diffCommits_info_83_fpWen; \
        force U_IF_NAME.io_diffCommits_info_83_vecWen = RTL_PATH.io_diffCommits_info_83_vecWen; \
        force U_IF_NAME.io_diffCommits_info_83_v0Wen = RTL_PATH.io_diffCommits_info_83_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_83_vlWen = RTL_PATH.io_diffCommits_info_83_vlWen; \
        force U_IF_NAME.io_diffCommits_info_84_ldest = RTL_PATH.io_diffCommits_info_84_ldest; \
        force U_IF_NAME.io_diffCommits_info_84_pdest = RTL_PATH.io_diffCommits_info_84_pdest; \
        force U_IF_NAME.io_diffCommits_info_84_rfWen = RTL_PATH.io_diffCommits_info_84_rfWen; \
        force U_IF_NAME.io_diffCommits_info_84_fpWen = RTL_PATH.io_diffCommits_info_84_fpWen; \
        force U_IF_NAME.io_diffCommits_info_84_vecWen = RTL_PATH.io_diffCommits_info_84_vecWen; \
        force U_IF_NAME.io_diffCommits_info_84_v0Wen = RTL_PATH.io_diffCommits_info_84_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_84_vlWen = RTL_PATH.io_diffCommits_info_84_vlWen; \
        force U_IF_NAME.io_diffCommits_info_85_ldest = RTL_PATH.io_diffCommits_info_85_ldest; \
        force U_IF_NAME.io_diffCommits_info_85_pdest = RTL_PATH.io_diffCommits_info_85_pdest; \
        force U_IF_NAME.io_diffCommits_info_85_rfWen = RTL_PATH.io_diffCommits_info_85_rfWen; \
        force U_IF_NAME.io_diffCommits_info_85_fpWen = RTL_PATH.io_diffCommits_info_85_fpWen; \
        force U_IF_NAME.io_diffCommits_info_85_vecWen = RTL_PATH.io_diffCommits_info_85_vecWen; \
        force U_IF_NAME.io_diffCommits_info_85_v0Wen = RTL_PATH.io_diffCommits_info_85_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_85_vlWen = RTL_PATH.io_diffCommits_info_85_vlWen; \
        force U_IF_NAME.io_diffCommits_info_86_ldest = RTL_PATH.io_diffCommits_info_86_ldest; \
        force U_IF_NAME.io_diffCommits_info_86_pdest = RTL_PATH.io_diffCommits_info_86_pdest; \
        force U_IF_NAME.io_diffCommits_info_86_rfWen = RTL_PATH.io_diffCommits_info_86_rfWen; \
        force U_IF_NAME.io_diffCommits_info_86_fpWen = RTL_PATH.io_diffCommits_info_86_fpWen; \
        force U_IF_NAME.io_diffCommits_info_86_vecWen = RTL_PATH.io_diffCommits_info_86_vecWen; \
        force U_IF_NAME.io_diffCommits_info_86_v0Wen = RTL_PATH.io_diffCommits_info_86_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_86_vlWen = RTL_PATH.io_diffCommits_info_86_vlWen; \
        force U_IF_NAME.io_diffCommits_info_87_ldest = RTL_PATH.io_diffCommits_info_87_ldest; \
        force U_IF_NAME.io_diffCommits_info_87_pdest = RTL_PATH.io_diffCommits_info_87_pdest; \
        force U_IF_NAME.io_diffCommits_info_87_rfWen = RTL_PATH.io_diffCommits_info_87_rfWen; \
        force U_IF_NAME.io_diffCommits_info_87_fpWen = RTL_PATH.io_diffCommits_info_87_fpWen; \
        force U_IF_NAME.io_diffCommits_info_87_vecWen = RTL_PATH.io_diffCommits_info_87_vecWen; \
        force U_IF_NAME.io_diffCommits_info_87_v0Wen = RTL_PATH.io_diffCommits_info_87_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_87_vlWen = RTL_PATH.io_diffCommits_info_87_vlWen; \
        force U_IF_NAME.io_diffCommits_info_88_ldest = RTL_PATH.io_diffCommits_info_88_ldest; \
        force U_IF_NAME.io_diffCommits_info_88_pdest = RTL_PATH.io_diffCommits_info_88_pdest; \
        force U_IF_NAME.io_diffCommits_info_88_rfWen = RTL_PATH.io_diffCommits_info_88_rfWen; \
        force U_IF_NAME.io_diffCommits_info_88_fpWen = RTL_PATH.io_diffCommits_info_88_fpWen; \
        force U_IF_NAME.io_diffCommits_info_88_vecWen = RTL_PATH.io_diffCommits_info_88_vecWen; \
        force U_IF_NAME.io_diffCommits_info_88_v0Wen = RTL_PATH.io_diffCommits_info_88_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_88_vlWen = RTL_PATH.io_diffCommits_info_88_vlWen; \
        force U_IF_NAME.io_diffCommits_info_89_ldest = RTL_PATH.io_diffCommits_info_89_ldest; \
        force U_IF_NAME.io_diffCommits_info_89_pdest = RTL_PATH.io_diffCommits_info_89_pdest; \
        force U_IF_NAME.io_diffCommits_info_89_rfWen = RTL_PATH.io_diffCommits_info_89_rfWen; \
        force U_IF_NAME.io_diffCommits_info_89_fpWen = RTL_PATH.io_diffCommits_info_89_fpWen; \
        force U_IF_NAME.io_diffCommits_info_89_vecWen = RTL_PATH.io_diffCommits_info_89_vecWen; \
        force U_IF_NAME.io_diffCommits_info_89_v0Wen = RTL_PATH.io_diffCommits_info_89_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_89_vlWen = RTL_PATH.io_diffCommits_info_89_vlWen; \
        force U_IF_NAME.io_diffCommits_info_90_ldest = RTL_PATH.io_diffCommits_info_90_ldest; \
        force U_IF_NAME.io_diffCommits_info_90_pdest = RTL_PATH.io_diffCommits_info_90_pdest; \
        force U_IF_NAME.io_diffCommits_info_90_rfWen = RTL_PATH.io_diffCommits_info_90_rfWen; \
        force U_IF_NAME.io_diffCommits_info_90_fpWen = RTL_PATH.io_diffCommits_info_90_fpWen; \
        force U_IF_NAME.io_diffCommits_info_90_vecWen = RTL_PATH.io_diffCommits_info_90_vecWen; \
        force U_IF_NAME.io_diffCommits_info_90_v0Wen = RTL_PATH.io_diffCommits_info_90_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_90_vlWen = RTL_PATH.io_diffCommits_info_90_vlWen; \
        force U_IF_NAME.io_diffCommits_info_91_ldest = RTL_PATH.io_diffCommits_info_91_ldest; \
        force U_IF_NAME.io_diffCommits_info_91_pdest = RTL_PATH.io_diffCommits_info_91_pdest; \
        force U_IF_NAME.io_diffCommits_info_91_rfWen = RTL_PATH.io_diffCommits_info_91_rfWen; \
        force U_IF_NAME.io_diffCommits_info_91_fpWen = RTL_PATH.io_diffCommits_info_91_fpWen; \
        force U_IF_NAME.io_diffCommits_info_91_vecWen = RTL_PATH.io_diffCommits_info_91_vecWen; \
        force U_IF_NAME.io_diffCommits_info_91_v0Wen = RTL_PATH.io_diffCommits_info_91_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_91_vlWen = RTL_PATH.io_diffCommits_info_91_vlWen; \
        force U_IF_NAME.io_diffCommits_info_92_ldest = RTL_PATH.io_diffCommits_info_92_ldest; \
        force U_IF_NAME.io_diffCommits_info_92_pdest = RTL_PATH.io_diffCommits_info_92_pdest; \
        force U_IF_NAME.io_diffCommits_info_92_rfWen = RTL_PATH.io_diffCommits_info_92_rfWen; \
        force U_IF_NAME.io_diffCommits_info_92_fpWen = RTL_PATH.io_diffCommits_info_92_fpWen; \
        force U_IF_NAME.io_diffCommits_info_92_vecWen = RTL_PATH.io_diffCommits_info_92_vecWen; \
        force U_IF_NAME.io_diffCommits_info_92_v0Wen = RTL_PATH.io_diffCommits_info_92_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_92_vlWen = RTL_PATH.io_diffCommits_info_92_vlWen; \
        force U_IF_NAME.io_diffCommits_info_93_ldest = RTL_PATH.io_diffCommits_info_93_ldest; \
        force U_IF_NAME.io_diffCommits_info_93_pdest = RTL_PATH.io_diffCommits_info_93_pdest; \
        force U_IF_NAME.io_diffCommits_info_93_rfWen = RTL_PATH.io_diffCommits_info_93_rfWen; \
        force U_IF_NAME.io_diffCommits_info_93_fpWen = RTL_PATH.io_diffCommits_info_93_fpWen; \
        force U_IF_NAME.io_diffCommits_info_93_vecWen = RTL_PATH.io_diffCommits_info_93_vecWen; \
        force U_IF_NAME.io_diffCommits_info_93_v0Wen = RTL_PATH.io_diffCommits_info_93_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_93_vlWen = RTL_PATH.io_diffCommits_info_93_vlWen; \
        force U_IF_NAME.io_diffCommits_info_94_ldest = RTL_PATH.io_diffCommits_info_94_ldest; \
        force U_IF_NAME.io_diffCommits_info_94_pdest = RTL_PATH.io_diffCommits_info_94_pdest; \
        force U_IF_NAME.io_diffCommits_info_94_rfWen = RTL_PATH.io_diffCommits_info_94_rfWen; \
        force U_IF_NAME.io_diffCommits_info_94_fpWen = RTL_PATH.io_diffCommits_info_94_fpWen; \
        force U_IF_NAME.io_diffCommits_info_94_vecWen = RTL_PATH.io_diffCommits_info_94_vecWen; \
        force U_IF_NAME.io_diffCommits_info_94_v0Wen = RTL_PATH.io_diffCommits_info_94_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_94_vlWen = RTL_PATH.io_diffCommits_info_94_vlWen; \
        force U_IF_NAME.io_diffCommits_info_95_ldest = RTL_PATH.io_diffCommits_info_95_ldest; \
        force U_IF_NAME.io_diffCommits_info_95_pdest = RTL_PATH.io_diffCommits_info_95_pdest; \
        force U_IF_NAME.io_diffCommits_info_95_rfWen = RTL_PATH.io_diffCommits_info_95_rfWen; \
        force U_IF_NAME.io_diffCommits_info_95_fpWen = RTL_PATH.io_diffCommits_info_95_fpWen; \
        force U_IF_NAME.io_diffCommits_info_95_vecWen = RTL_PATH.io_diffCommits_info_95_vecWen; \
        force U_IF_NAME.io_diffCommits_info_95_v0Wen = RTL_PATH.io_diffCommits_info_95_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_95_vlWen = RTL_PATH.io_diffCommits_info_95_vlWen; \
        force U_IF_NAME.io_diffCommits_info_96_ldest = RTL_PATH.io_diffCommits_info_96_ldest; \
        force U_IF_NAME.io_diffCommits_info_96_pdest = RTL_PATH.io_diffCommits_info_96_pdest; \
        force U_IF_NAME.io_diffCommits_info_96_rfWen = RTL_PATH.io_diffCommits_info_96_rfWen; \
        force U_IF_NAME.io_diffCommits_info_96_fpWen = RTL_PATH.io_diffCommits_info_96_fpWen; \
        force U_IF_NAME.io_diffCommits_info_96_vecWen = RTL_PATH.io_diffCommits_info_96_vecWen; \
        force U_IF_NAME.io_diffCommits_info_96_v0Wen = RTL_PATH.io_diffCommits_info_96_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_96_vlWen = RTL_PATH.io_diffCommits_info_96_vlWen; \
        force U_IF_NAME.io_diffCommits_info_97_ldest = RTL_PATH.io_diffCommits_info_97_ldest; \
        force U_IF_NAME.io_diffCommits_info_97_pdest = RTL_PATH.io_diffCommits_info_97_pdest; \
        force U_IF_NAME.io_diffCommits_info_97_rfWen = RTL_PATH.io_diffCommits_info_97_rfWen; \
        force U_IF_NAME.io_diffCommits_info_97_fpWen = RTL_PATH.io_diffCommits_info_97_fpWen; \
        force U_IF_NAME.io_diffCommits_info_97_vecWen = RTL_PATH.io_diffCommits_info_97_vecWen; \
        force U_IF_NAME.io_diffCommits_info_97_v0Wen = RTL_PATH.io_diffCommits_info_97_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_97_vlWen = RTL_PATH.io_diffCommits_info_97_vlWen; \
        force U_IF_NAME.io_diffCommits_info_98_ldest = RTL_PATH.io_diffCommits_info_98_ldest; \
        force U_IF_NAME.io_diffCommits_info_98_pdest = RTL_PATH.io_diffCommits_info_98_pdest; \
        force U_IF_NAME.io_diffCommits_info_98_rfWen = RTL_PATH.io_diffCommits_info_98_rfWen; \
        force U_IF_NAME.io_diffCommits_info_98_fpWen = RTL_PATH.io_diffCommits_info_98_fpWen; \
        force U_IF_NAME.io_diffCommits_info_98_vecWen = RTL_PATH.io_diffCommits_info_98_vecWen; \
        force U_IF_NAME.io_diffCommits_info_98_v0Wen = RTL_PATH.io_diffCommits_info_98_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_98_vlWen = RTL_PATH.io_diffCommits_info_98_vlWen; \
        force U_IF_NAME.io_diffCommits_info_99_ldest = RTL_PATH.io_diffCommits_info_99_ldest; \
        force U_IF_NAME.io_diffCommits_info_99_pdest = RTL_PATH.io_diffCommits_info_99_pdest; \
        force U_IF_NAME.io_diffCommits_info_99_rfWen = RTL_PATH.io_diffCommits_info_99_rfWen; \
        force U_IF_NAME.io_diffCommits_info_99_fpWen = RTL_PATH.io_diffCommits_info_99_fpWen; \
        force U_IF_NAME.io_diffCommits_info_99_vecWen = RTL_PATH.io_diffCommits_info_99_vecWen; \
        force U_IF_NAME.io_diffCommits_info_99_v0Wen = RTL_PATH.io_diffCommits_info_99_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_99_vlWen = RTL_PATH.io_diffCommits_info_99_vlWen; \
        force U_IF_NAME.io_diffCommits_info_100_ldest = RTL_PATH.io_diffCommits_info_100_ldest; \
        force U_IF_NAME.io_diffCommits_info_100_pdest = RTL_PATH.io_diffCommits_info_100_pdest; \
        force U_IF_NAME.io_diffCommits_info_100_rfWen = RTL_PATH.io_diffCommits_info_100_rfWen; \
        force U_IF_NAME.io_diffCommits_info_100_fpWen = RTL_PATH.io_diffCommits_info_100_fpWen; \
        force U_IF_NAME.io_diffCommits_info_100_vecWen = RTL_PATH.io_diffCommits_info_100_vecWen; \
        force U_IF_NAME.io_diffCommits_info_100_v0Wen = RTL_PATH.io_diffCommits_info_100_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_100_vlWen = RTL_PATH.io_diffCommits_info_100_vlWen; \
        force U_IF_NAME.io_diffCommits_info_101_ldest = RTL_PATH.io_diffCommits_info_101_ldest; \
        force U_IF_NAME.io_diffCommits_info_101_pdest = RTL_PATH.io_diffCommits_info_101_pdest; \
        force U_IF_NAME.io_diffCommits_info_101_rfWen = RTL_PATH.io_diffCommits_info_101_rfWen; \
        force U_IF_NAME.io_diffCommits_info_101_fpWen = RTL_PATH.io_diffCommits_info_101_fpWen; \
        force U_IF_NAME.io_diffCommits_info_101_vecWen = RTL_PATH.io_diffCommits_info_101_vecWen; \
        force U_IF_NAME.io_diffCommits_info_101_v0Wen = RTL_PATH.io_diffCommits_info_101_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_101_vlWen = RTL_PATH.io_diffCommits_info_101_vlWen; \
        force U_IF_NAME.io_diffCommits_info_102_ldest = RTL_PATH.io_diffCommits_info_102_ldest; \
        force U_IF_NAME.io_diffCommits_info_102_pdest = RTL_PATH.io_diffCommits_info_102_pdest; \
        force U_IF_NAME.io_diffCommits_info_102_rfWen = RTL_PATH.io_diffCommits_info_102_rfWen; \
        force U_IF_NAME.io_diffCommits_info_102_fpWen = RTL_PATH.io_diffCommits_info_102_fpWen; \
        force U_IF_NAME.io_diffCommits_info_102_vecWen = RTL_PATH.io_diffCommits_info_102_vecWen; \
        force U_IF_NAME.io_diffCommits_info_102_v0Wen = RTL_PATH.io_diffCommits_info_102_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_102_vlWen = RTL_PATH.io_diffCommits_info_102_vlWen; \
        force U_IF_NAME.io_diffCommits_info_103_ldest = RTL_PATH.io_diffCommits_info_103_ldest; \
        force U_IF_NAME.io_diffCommits_info_103_pdest = RTL_PATH.io_diffCommits_info_103_pdest; \
        force U_IF_NAME.io_diffCommits_info_103_rfWen = RTL_PATH.io_diffCommits_info_103_rfWen; \
        force U_IF_NAME.io_diffCommits_info_103_fpWen = RTL_PATH.io_diffCommits_info_103_fpWen; \
        force U_IF_NAME.io_diffCommits_info_103_vecWen = RTL_PATH.io_diffCommits_info_103_vecWen; \
        force U_IF_NAME.io_diffCommits_info_103_v0Wen = RTL_PATH.io_diffCommits_info_103_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_103_vlWen = RTL_PATH.io_diffCommits_info_103_vlWen; \
        force U_IF_NAME.io_diffCommits_info_104_ldest = RTL_PATH.io_diffCommits_info_104_ldest; \
        force U_IF_NAME.io_diffCommits_info_104_pdest = RTL_PATH.io_diffCommits_info_104_pdest; \
        force U_IF_NAME.io_diffCommits_info_104_rfWen = RTL_PATH.io_diffCommits_info_104_rfWen; \
        force U_IF_NAME.io_diffCommits_info_104_fpWen = RTL_PATH.io_diffCommits_info_104_fpWen; \
        force U_IF_NAME.io_diffCommits_info_104_vecWen = RTL_PATH.io_diffCommits_info_104_vecWen; \
        force U_IF_NAME.io_diffCommits_info_104_v0Wen = RTL_PATH.io_diffCommits_info_104_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_104_vlWen = RTL_PATH.io_diffCommits_info_104_vlWen; \
        force U_IF_NAME.io_diffCommits_info_105_ldest = RTL_PATH.io_diffCommits_info_105_ldest; \
        force U_IF_NAME.io_diffCommits_info_105_pdest = RTL_PATH.io_diffCommits_info_105_pdest; \
        force U_IF_NAME.io_diffCommits_info_105_rfWen = RTL_PATH.io_diffCommits_info_105_rfWen; \
        force U_IF_NAME.io_diffCommits_info_105_fpWen = RTL_PATH.io_diffCommits_info_105_fpWen; \
        force U_IF_NAME.io_diffCommits_info_105_vecWen = RTL_PATH.io_diffCommits_info_105_vecWen; \
        force U_IF_NAME.io_diffCommits_info_105_v0Wen = RTL_PATH.io_diffCommits_info_105_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_105_vlWen = RTL_PATH.io_diffCommits_info_105_vlWen; \
        force U_IF_NAME.io_diffCommits_info_106_ldest = RTL_PATH.io_diffCommits_info_106_ldest; \
        force U_IF_NAME.io_diffCommits_info_106_pdest = RTL_PATH.io_diffCommits_info_106_pdest; \
        force U_IF_NAME.io_diffCommits_info_106_rfWen = RTL_PATH.io_diffCommits_info_106_rfWen; \
        force U_IF_NAME.io_diffCommits_info_106_fpWen = RTL_PATH.io_diffCommits_info_106_fpWen; \
        force U_IF_NAME.io_diffCommits_info_106_vecWen = RTL_PATH.io_diffCommits_info_106_vecWen; \
        force U_IF_NAME.io_diffCommits_info_106_v0Wen = RTL_PATH.io_diffCommits_info_106_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_106_vlWen = RTL_PATH.io_diffCommits_info_106_vlWen; \
        force U_IF_NAME.io_diffCommits_info_107_ldest = RTL_PATH.io_diffCommits_info_107_ldest; \
        force U_IF_NAME.io_diffCommits_info_107_pdest = RTL_PATH.io_diffCommits_info_107_pdest; \
        force U_IF_NAME.io_diffCommits_info_107_rfWen = RTL_PATH.io_diffCommits_info_107_rfWen; \
        force U_IF_NAME.io_diffCommits_info_107_fpWen = RTL_PATH.io_diffCommits_info_107_fpWen; \
        force U_IF_NAME.io_diffCommits_info_107_vecWen = RTL_PATH.io_diffCommits_info_107_vecWen; \
        force U_IF_NAME.io_diffCommits_info_107_v0Wen = RTL_PATH.io_diffCommits_info_107_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_107_vlWen = RTL_PATH.io_diffCommits_info_107_vlWen; \
        force U_IF_NAME.io_diffCommits_info_108_ldest = RTL_PATH.io_diffCommits_info_108_ldest; \
        force U_IF_NAME.io_diffCommits_info_108_pdest = RTL_PATH.io_diffCommits_info_108_pdest; \
        force U_IF_NAME.io_diffCommits_info_108_rfWen = RTL_PATH.io_diffCommits_info_108_rfWen; \
        force U_IF_NAME.io_diffCommits_info_108_fpWen = RTL_PATH.io_diffCommits_info_108_fpWen; \
        force U_IF_NAME.io_diffCommits_info_108_vecWen = RTL_PATH.io_diffCommits_info_108_vecWen; \
        force U_IF_NAME.io_diffCommits_info_108_v0Wen = RTL_PATH.io_diffCommits_info_108_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_108_vlWen = RTL_PATH.io_diffCommits_info_108_vlWen; \
        force U_IF_NAME.io_diffCommits_info_109_ldest = RTL_PATH.io_diffCommits_info_109_ldest; \
        force U_IF_NAME.io_diffCommits_info_109_pdest = RTL_PATH.io_diffCommits_info_109_pdest; \
        force U_IF_NAME.io_diffCommits_info_109_rfWen = RTL_PATH.io_diffCommits_info_109_rfWen; \
        force U_IF_NAME.io_diffCommits_info_109_fpWen = RTL_PATH.io_diffCommits_info_109_fpWen; \
        force U_IF_NAME.io_diffCommits_info_109_vecWen = RTL_PATH.io_diffCommits_info_109_vecWen; \
        force U_IF_NAME.io_diffCommits_info_109_v0Wen = RTL_PATH.io_diffCommits_info_109_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_109_vlWen = RTL_PATH.io_diffCommits_info_109_vlWen; \
        force U_IF_NAME.io_diffCommits_info_110_ldest = RTL_PATH.io_diffCommits_info_110_ldest; \
        force U_IF_NAME.io_diffCommits_info_110_pdest = RTL_PATH.io_diffCommits_info_110_pdest; \
        force U_IF_NAME.io_diffCommits_info_110_rfWen = RTL_PATH.io_diffCommits_info_110_rfWen; \
        force U_IF_NAME.io_diffCommits_info_110_fpWen = RTL_PATH.io_diffCommits_info_110_fpWen; \
        force U_IF_NAME.io_diffCommits_info_110_vecWen = RTL_PATH.io_diffCommits_info_110_vecWen; \
        force U_IF_NAME.io_diffCommits_info_110_v0Wen = RTL_PATH.io_diffCommits_info_110_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_110_vlWen = RTL_PATH.io_diffCommits_info_110_vlWen; \
        force U_IF_NAME.io_diffCommits_info_111_ldest = RTL_PATH.io_diffCommits_info_111_ldest; \
        force U_IF_NAME.io_diffCommits_info_111_pdest = RTL_PATH.io_diffCommits_info_111_pdest; \
        force U_IF_NAME.io_diffCommits_info_111_rfWen = RTL_PATH.io_diffCommits_info_111_rfWen; \
        force U_IF_NAME.io_diffCommits_info_111_fpWen = RTL_PATH.io_diffCommits_info_111_fpWen; \
        force U_IF_NAME.io_diffCommits_info_111_vecWen = RTL_PATH.io_diffCommits_info_111_vecWen; \
        force U_IF_NAME.io_diffCommits_info_111_v0Wen = RTL_PATH.io_diffCommits_info_111_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_111_vlWen = RTL_PATH.io_diffCommits_info_111_vlWen; \
        force U_IF_NAME.io_diffCommits_info_112_ldest = RTL_PATH.io_diffCommits_info_112_ldest; \
        force U_IF_NAME.io_diffCommits_info_112_pdest = RTL_PATH.io_diffCommits_info_112_pdest; \
        force U_IF_NAME.io_diffCommits_info_112_rfWen = RTL_PATH.io_diffCommits_info_112_rfWen; \
        force U_IF_NAME.io_diffCommits_info_112_fpWen = RTL_PATH.io_diffCommits_info_112_fpWen; \
        force U_IF_NAME.io_diffCommits_info_112_vecWen = RTL_PATH.io_diffCommits_info_112_vecWen; \
        force U_IF_NAME.io_diffCommits_info_112_v0Wen = RTL_PATH.io_diffCommits_info_112_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_112_vlWen = RTL_PATH.io_diffCommits_info_112_vlWen; \
        force U_IF_NAME.io_diffCommits_info_113_ldest = RTL_PATH.io_diffCommits_info_113_ldest; \
        force U_IF_NAME.io_diffCommits_info_113_pdest = RTL_PATH.io_diffCommits_info_113_pdest; \
        force U_IF_NAME.io_diffCommits_info_113_rfWen = RTL_PATH.io_diffCommits_info_113_rfWen; \
        force U_IF_NAME.io_diffCommits_info_113_fpWen = RTL_PATH.io_diffCommits_info_113_fpWen; \
        force U_IF_NAME.io_diffCommits_info_113_vecWen = RTL_PATH.io_diffCommits_info_113_vecWen; \
        force U_IF_NAME.io_diffCommits_info_113_v0Wen = RTL_PATH.io_diffCommits_info_113_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_113_vlWen = RTL_PATH.io_diffCommits_info_113_vlWen; \
        force U_IF_NAME.io_diffCommits_info_114_ldest = RTL_PATH.io_diffCommits_info_114_ldest; \
        force U_IF_NAME.io_diffCommits_info_114_pdest = RTL_PATH.io_diffCommits_info_114_pdest; \
        force U_IF_NAME.io_diffCommits_info_114_rfWen = RTL_PATH.io_diffCommits_info_114_rfWen; \
        force U_IF_NAME.io_diffCommits_info_114_fpWen = RTL_PATH.io_diffCommits_info_114_fpWen; \
        force U_IF_NAME.io_diffCommits_info_114_vecWen = RTL_PATH.io_diffCommits_info_114_vecWen; \
        force U_IF_NAME.io_diffCommits_info_114_v0Wen = RTL_PATH.io_diffCommits_info_114_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_114_vlWen = RTL_PATH.io_diffCommits_info_114_vlWen; \
        force U_IF_NAME.io_diffCommits_info_115_ldest = RTL_PATH.io_diffCommits_info_115_ldest; \
        force U_IF_NAME.io_diffCommits_info_115_pdest = RTL_PATH.io_diffCommits_info_115_pdest; \
        force U_IF_NAME.io_diffCommits_info_115_rfWen = RTL_PATH.io_diffCommits_info_115_rfWen; \
        force U_IF_NAME.io_diffCommits_info_115_fpWen = RTL_PATH.io_diffCommits_info_115_fpWen; \
        force U_IF_NAME.io_diffCommits_info_115_vecWen = RTL_PATH.io_diffCommits_info_115_vecWen; \
        force U_IF_NAME.io_diffCommits_info_115_v0Wen = RTL_PATH.io_diffCommits_info_115_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_115_vlWen = RTL_PATH.io_diffCommits_info_115_vlWen; \
        force U_IF_NAME.io_diffCommits_info_116_ldest = RTL_PATH.io_diffCommits_info_116_ldest; \
        force U_IF_NAME.io_diffCommits_info_116_pdest = RTL_PATH.io_diffCommits_info_116_pdest; \
        force U_IF_NAME.io_diffCommits_info_116_rfWen = RTL_PATH.io_diffCommits_info_116_rfWen; \
        force U_IF_NAME.io_diffCommits_info_116_fpWen = RTL_PATH.io_diffCommits_info_116_fpWen; \
        force U_IF_NAME.io_diffCommits_info_116_vecWen = RTL_PATH.io_diffCommits_info_116_vecWen; \
        force U_IF_NAME.io_diffCommits_info_116_v0Wen = RTL_PATH.io_diffCommits_info_116_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_116_vlWen = RTL_PATH.io_diffCommits_info_116_vlWen; \
        force U_IF_NAME.io_diffCommits_info_117_ldest = RTL_PATH.io_diffCommits_info_117_ldest; \
        force U_IF_NAME.io_diffCommits_info_117_pdest = RTL_PATH.io_diffCommits_info_117_pdest; \
        force U_IF_NAME.io_diffCommits_info_117_rfWen = RTL_PATH.io_diffCommits_info_117_rfWen; \
        force U_IF_NAME.io_diffCommits_info_117_fpWen = RTL_PATH.io_diffCommits_info_117_fpWen; \
        force U_IF_NAME.io_diffCommits_info_117_vecWen = RTL_PATH.io_diffCommits_info_117_vecWen; \
        force U_IF_NAME.io_diffCommits_info_117_v0Wen = RTL_PATH.io_diffCommits_info_117_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_117_vlWen = RTL_PATH.io_diffCommits_info_117_vlWen; \
        force U_IF_NAME.io_diffCommits_info_118_ldest = RTL_PATH.io_diffCommits_info_118_ldest; \
        force U_IF_NAME.io_diffCommits_info_118_pdest = RTL_PATH.io_diffCommits_info_118_pdest; \
        force U_IF_NAME.io_diffCommits_info_118_rfWen = RTL_PATH.io_diffCommits_info_118_rfWen; \
        force U_IF_NAME.io_diffCommits_info_118_fpWen = RTL_PATH.io_diffCommits_info_118_fpWen; \
        force U_IF_NAME.io_diffCommits_info_118_vecWen = RTL_PATH.io_diffCommits_info_118_vecWen; \
        force U_IF_NAME.io_diffCommits_info_118_v0Wen = RTL_PATH.io_diffCommits_info_118_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_118_vlWen = RTL_PATH.io_diffCommits_info_118_vlWen; \
        force U_IF_NAME.io_diffCommits_info_119_ldest = RTL_PATH.io_diffCommits_info_119_ldest; \
        force U_IF_NAME.io_diffCommits_info_119_pdest = RTL_PATH.io_diffCommits_info_119_pdest; \
        force U_IF_NAME.io_diffCommits_info_119_rfWen = RTL_PATH.io_diffCommits_info_119_rfWen; \
        force U_IF_NAME.io_diffCommits_info_119_fpWen = RTL_PATH.io_diffCommits_info_119_fpWen; \
        force U_IF_NAME.io_diffCommits_info_119_vecWen = RTL_PATH.io_diffCommits_info_119_vecWen; \
        force U_IF_NAME.io_diffCommits_info_119_v0Wen = RTL_PATH.io_diffCommits_info_119_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_119_vlWen = RTL_PATH.io_diffCommits_info_119_vlWen; \
        force U_IF_NAME.io_diffCommits_info_120_ldest = RTL_PATH.io_diffCommits_info_120_ldest; \
        force U_IF_NAME.io_diffCommits_info_120_pdest = RTL_PATH.io_diffCommits_info_120_pdest; \
        force U_IF_NAME.io_diffCommits_info_120_rfWen = RTL_PATH.io_diffCommits_info_120_rfWen; \
        force U_IF_NAME.io_diffCommits_info_120_fpWen = RTL_PATH.io_diffCommits_info_120_fpWen; \
        force U_IF_NAME.io_diffCommits_info_120_vecWen = RTL_PATH.io_diffCommits_info_120_vecWen; \
        force U_IF_NAME.io_diffCommits_info_120_v0Wen = RTL_PATH.io_diffCommits_info_120_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_120_vlWen = RTL_PATH.io_diffCommits_info_120_vlWen; \
        force U_IF_NAME.io_diffCommits_info_121_ldest = RTL_PATH.io_diffCommits_info_121_ldest; \
        force U_IF_NAME.io_diffCommits_info_121_pdest = RTL_PATH.io_diffCommits_info_121_pdest; \
        force U_IF_NAME.io_diffCommits_info_121_rfWen = RTL_PATH.io_diffCommits_info_121_rfWen; \
        force U_IF_NAME.io_diffCommits_info_121_fpWen = RTL_PATH.io_diffCommits_info_121_fpWen; \
        force U_IF_NAME.io_diffCommits_info_121_vecWen = RTL_PATH.io_diffCommits_info_121_vecWen; \
        force U_IF_NAME.io_diffCommits_info_121_v0Wen = RTL_PATH.io_diffCommits_info_121_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_121_vlWen = RTL_PATH.io_diffCommits_info_121_vlWen; \
        force U_IF_NAME.io_diffCommits_info_122_ldest = RTL_PATH.io_diffCommits_info_122_ldest; \
        force U_IF_NAME.io_diffCommits_info_122_pdest = RTL_PATH.io_diffCommits_info_122_pdest; \
        force U_IF_NAME.io_diffCommits_info_122_rfWen = RTL_PATH.io_diffCommits_info_122_rfWen; \
        force U_IF_NAME.io_diffCommits_info_122_fpWen = RTL_PATH.io_diffCommits_info_122_fpWen; \
        force U_IF_NAME.io_diffCommits_info_122_vecWen = RTL_PATH.io_diffCommits_info_122_vecWen; \
        force U_IF_NAME.io_diffCommits_info_122_v0Wen = RTL_PATH.io_diffCommits_info_122_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_122_vlWen = RTL_PATH.io_diffCommits_info_122_vlWen; \
        force U_IF_NAME.io_diffCommits_info_123_ldest = RTL_PATH.io_diffCommits_info_123_ldest; \
        force U_IF_NAME.io_diffCommits_info_123_pdest = RTL_PATH.io_diffCommits_info_123_pdest; \
        force U_IF_NAME.io_diffCommits_info_123_rfWen = RTL_PATH.io_diffCommits_info_123_rfWen; \
        force U_IF_NAME.io_diffCommits_info_123_fpWen = RTL_PATH.io_diffCommits_info_123_fpWen; \
        force U_IF_NAME.io_diffCommits_info_123_vecWen = RTL_PATH.io_diffCommits_info_123_vecWen; \
        force U_IF_NAME.io_diffCommits_info_123_v0Wen = RTL_PATH.io_diffCommits_info_123_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_123_vlWen = RTL_PATH.io_diffCommits_info_123_vlWen; \
        force U_IF_NAME.io_diffCommits_info_124_ldest = RTL_PATH.io_diffCommits_info_124_ldest; \
        force U_IF_NAME.io_diffCommits_info_124_pdest = RTL_PATH.io_diffCommits_info_124_pdest; \
        force U_IF_NAME.io_diffCommits_info_124_rfWen = RTL_PATH.io_diffCommits_info_124_rfWen; \
        force U_IF_NAME.io_diffCommits_info_124_fpWen = RTL_PATH.io_diffCommits_info_124_fpWen; \
        force U_IF_NAME.io_diffCommits_info_124_vecWen = RTL_PATH.io_diffCommits_info_124_vecWen; \
        force U_IF_NAME.io_diffCommits_info_124_v0Wen = RTL_PATH.io_diffCommits_info_124_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_124_vlWen = RTL_PATH.io_diffCommits_info_124_vlWen; \
        force U_IF_NAME.io_diffCommits_info_125_ldest = RTL_PATH.io_diffCommits_info_125_ldest; \
        force U_IF_NAME.io_diffCommits_info_125_pdest = RTL_PATH.io_diffCommits_info_125_pdest; \
        force U_IF_NAME.io_diffCommits_info_125_rfWen = RTL_PATH.io_diffCommits_info_125_rfWen; \
        force U_IF_NAME.io_diffCommits_info_125_fpWen = RTL_PATH.io_diffCommits_info_125_fpWen; \
        force U_IF_NAME.io_diffCommits_info_125_vecWen = RTL_PATH.io_diffCommits_info_125_vecWen; \
        force U_IF_NAME.io_diffCommits_info_125_v0Wen = RTL_PATH.io_diffCommits_info_125_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_125_vlWen = RTL_PATH.io_diffCommits_info_125_vlWen; \
        force U_IF_NAME.io_diffCommits_info_126_ldest = RTL_PATH.io_diffCommits_info_126_ldest; \
        force U_IF_NAME.io_diffCommits_info_126_pdest = RTL_PATH.io_diffCommits_info_126_pdest; \
        force U_IF_NAME.io_diffCommits_info_126_rfWen = RTL_PATH.io_diffCommits_info_126_rfWen; \
        force U_IF_NAME.io_diffCommits_info_126_fpWen = RTL_PATH.io_diffCommits_info_126_fpWen; \
        force U_IF_NAME.io_diffCommits_info_126_vecWen = RTL_PATH.io_diffCommits_info_126_vecWen; \
        force U_IF_NAME.io_diffCommits_info_126_v0Wen = RTL_PATH.io_diffCommits_info_126_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_126_vlWen = RTL_PATH.io_diffCommits_info_126_vlWen; \
        force U_IF_NAME.io_diffCommits_info_127_ldest = RTL_PATH.io_diffCommits_info_127_ldest; \
        force U_IF_NAME.io_diffCommits_info_127_pdest = RTL_PATH.io_diffCommits_info_127_pdest; \
        force U_IF_NAME.io_diffCommits_info_127_rfWen = RTL_PATH.io_diffCommits_info_127_rfWen; \
        force U_IF_NAME.io_diffCommits_info_127_fpWen = RTL_PATH.io_diffCommits_info_127_fpWen; \
        force U_IF_NAME.io_diffCommits_info_127_vecWen = RTL_PATH.io_diffCommits_info_127_vecWen; \
        force U_IF_NAME.io_diffCommits_info_127_v0Wen = RTL_PATH.io_diffCommits_info_127_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_127_vlWen = RTL_PATH.io_diffCommits_info_127_vlWen; \
        force U_IF_NAME.io_diffCommits_info_128_ldest = RTL_PATH.io_diffCommits_info_128_ldest; \
        force U_IF_NAME.io_diffCommits_info_128_pdest = RTL_PATH.io_diffCommits_info_128_pdest; \
        force U_IF_NAME.io_diffCommits_info_128_rfWen = RTL_PATH.io_diffCommits_info_128_rfWen; \
        force U_IF_NAME.io_diffCommits_info_128_fpWen = RTL_PATH.io_diffCommits_info_128_fpWen; \
        force U_IF_NAME.io_diffCommits_info_128_vecWen = RTL_PATH.io_diffCommits_info_128_vecWen; \
        force U_IF_NAME.io_diffCommits_info_128_v0Wen = RTL_PATH.io_diffCommits_info_128_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_128_vlWen = RTL_PATH.io_diffCommits_info_128_vlWen; \
        force U_IF_NAME.io_diffCommits_info_129_ldest = RTL_PATH.io_diffCommits_info_129_ldest; \
        force U_IF_NAME.io_diffCommits_info_129_pdest = RTL_PATH.io_diffCommits_info_129_pdest; \
        force U_IF_NAME.io_diffCommits_info_129_rfWen = RTL_PATH.io_diffCommits_info_129_rfWen; \
        force U_IF_NAME.io_diffCommits_info_129_fpWen = RTL_PATH.io_diffCommits_info_129_fpWen; \
        force U_IF_NAME.io_diffCommits_info_129_vecWen = RTL_PATH.io_diffCommits_info_129_vecWen; \
        force U_IF_NAME.io_diffCommits_info_129_v0Wen = RTL_PATH.io_diffCommits_info_129_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_129_vlWen = RTL_PATH.io_diffCommits_info_129_vlWen; \
        force U_IF_NAME.io_diffCommits_info_130_ldest = RTL_PATH.io_diffCommits_info_130_ldest; \
        force U_IF_NAME.io_diffCommits_info_130_pdest = RTL_PATH.io_diffCommits_info_130_pdest; \
        force U_IF_NAME.io_diffCommits_info_130_rfWen = RTL_PATH.io_diffCommits_info_130_rfWen; \
        force U_IF_NAME.io_diffCommits_info_130_fpWen = RTL_PATH.io_diffCommits_info_130_fpWen; \
        force U_IF_NAME.io_diffCommits_info_130_vecWen = RTL_PATH.io_diffCommits_info_130_vecWen; \
        force U_IF_NAME.io_diffCommits_info_130_v0Wen = RTL_PATH.io_diffCommits_info_130_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_130_vlWen = RTL_PATH.io_diffCommits_info_130_vlWen; \
        force U_IF_NAME.io_diffCommits_info_131_ldest = RTL_PATH.io_diffCommits_info_131_ldest; \
        force U_IF_NAME.io_diffCommits_info_131_pdest = RTL_PATH.io_diffCommits_info_131_pdest; \
        force U_IF_NAME.io_diffCommits_info_131_rfWen = RTL_PATH.io_diffCommits_info_131_rfWen; \
        force U_IF_NAME.io_diffCommits_info_131_fpWen = RTL_PATH.io_diffCommits_info_131_fpWen; \
        force U_IF_NAME.io_diffCommits_info_131_vecWen = RTL_PATH.io_diffCommits_info_131_vecWen; \
        force U_IF_NAME.io_diffCommits_info_131_v0Wen = RTL_PATH.io_diffCommits_info_131_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_131_vlWen = RTL_PATH.io_diffCommits_info_131_vlWen; \
        force U_IF_NAME.io_diffCommits_info_132_ldest = RTL_PATH.io_diffCommits_info_132_ldest; \
        force U_IF_NAME.io_diffCommits_info_132_pdest = RTL_PATH.io_diffCommits_info_132_pdest; \
        force U_IF_NAME.io_diffCommits_info_132_rfWen = RTL_PATH.io_diffCommits_info_132_rfWen; \
        force U_IF_NAME.io_diffCommits_info_132_fpWen = RTL_PATH.io_diffCommits_info_132_fpWen; \
        force U_IF_NAME.io_diffCommits_info_132_vecWen = RTL_PATH.io_diffCommits_info_132_vecWen; \
        force U_IF_NAME.io_diffCommits_info_132_v0Wen = RTL_PATH.io_diffCommits_info_132_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_132_vlWen = RTL_PATH.io_diffCommits_info_132_vlWen; \
        force U_IF_NAME.io_diffCommits_info_133_ldest = RTL_PATH.io_diffCommits_info_133_ldest; \
        force U_IF_NAME.io_diffCommits_info_133_pdest = RTL_PATH.io_diffCommits_info_133_pdest; \
        force U_IF_NAME.io_diffCommits_info_133_rfWen = RTL_PATH.io_diffCommits_info_133_rfWen; \
        force U_IF_NAME.io_diffCommits_info_133_fpWen = RTL_PATH.io_diffCommits_info_133_fpWen; \
        force U_IF_NAME.io_diffCommits_info_133_vecWen = RTL_PATH.io_diffCommits_info_133_vecWen; \
        force U_IF_NAME.io_diffCommits_info_133_v0Wen = RTL_PATH.io_diffCommits_info_133_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_133_vlWen = RTL_PATH.io_diffCommits_info_133_vlWen; \
        force U_IF_NAME.io_diffCommits_info_134_ldest = RTL_PATH.io_diffCommits_info_134_ldest; \
        force U_IF_NAME.io_diffCommits_info_134_pdest = RTL_PATH.io_diffCommits_info_134_pdest; \
        force U_IF_NAME.io_diffCommits_info_134_rfWen = RTL_PATH.io_diffCommits_info_134_rfWen; \
        force U_IF_NAME.io_diffCommits_info_134_fpWen = RTL_PATH.io_diffCommits_info_134_fpWen; \
        force U_IF_NAME.io_diffCommits_info_134_vecWen = RTL_PATH.io_diffCommits_info_134_vecWen; \
        force U_IF_NAME.io_diffCommits_info_134_v0Wen = RTL_PATH.io_diffCommits_info_134_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_134_vlWen = RTL_PATH.io_diffCommits_info_134_vlWen; \
        force U_IF_NAME.io_diffCommits_info_135_ldest = RTL_PATH.io_diffCommits_info_135_ldest; \
        force U_IF_NAME.io_diffCommits_info_135_pdest = RTL_PATH.io_diffCommits_info_135_pdest; \
        force U_IF_NAME.io_diffCommits_info_135_rfWen = RTL_PATH.io_diffCommits_info_135_rfWen; \
        force U_IF_NAME.io_diffCommits_info_135_fpWen = RTL_PATH.io_diffCommits_info_135_fpWen; \
        force U_IF_NAME.io_diffCommits_info_135_vecWen = RTL_PATH.io_diffCommits_info_135_vecWen; \
        force U_IF_NAME.io_diffCommits_info_135_v0Wen = RTL_PATH.io_diffCommits_info_135_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_135_vlWen = RTL_PATH.io_diffCommits_info_135_vlWen; \
        force U_IF_NAME.io_diffCommits_info_136_ldest = RTL_PATH.io_diffCommits_info_136_ldest; \
        force U_IF_NAME.io_diffCommits_info_136_pdest = RTL_PATH.io_diffCommits_info_136_pdest; \
        force U_IF_NAME.io_diffCommits_info_136_rfWen = RTL_PATH.io_diffCommits_info_136_rfWen; \
        force U_IF_NAME.io_diffCommits_info_136_fpWen = RTL_PATH.io_diffCommits_info_136_fpWen; \
        force U_IF_NAME.io_diffCommits_info_136_vecWen = RTL_PATH.io_diffCommits_info_136_vecWen; \
        force U_IF_NAME.io_diffCommits_info_136_v0Wen = RTL_PATH.io_diffCommits_info_136_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_136_vlWen = RTL_PATH.io_diffCommits_info_136_vlWen; \
        force U_IF_NAME.io_diffCommits_info_137_ldest = RTL_PATH.io_diffCommits_info_137_ldest; \
        force U_IF_NAME.io_diffCommits_info_137_pdest = RTL_PATH.io_diffCommits_info_137_pdest; \
        force U_IF_NAME.io_diffCommits_info_137_rfWen = RTL_PATH.io_diffCommits_info_137_rfWen; \
        force U_IF_NAME.io_diffCommits_info_137_fpWen = RTL_PATH.io_diffCommits_info_137_fpWen; \
        force U_IF_NAME.io_diffCommits_info_137_vecWen = RTL_PATH.io_diffCommits_info_137_vecWen; \
        force U_IF_NAME.io_diffCommits_info_137_v0Wen = RTL_PATH.io_diffCommits_info_137_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_137_vlWen = RTL_PATH.io_diffCommits_info_137_vlWen; \
        force U_IF_NAME.io_diffCommits_info_138_ldest = RTL_PATH.io_diffCommits_info_138_ldest; \
        force U_IF_NAME.io_diffCommits_info_138_pdest = RTL_PATH.io_diffCommits_info_138_pdest; \
        force U_IF_NAME.io_diffCommits_info_138_rfWen = RTL_PATH.io_diffCommits_info_138_rfWen; \
        force U_IF_NAME.io_diffCommits_info_138_fpWen = RTL_PATH.io_diffCommits_info_138_fpWen; \
        force U_IF_NAME.io_diffCommits_info_138_vecWen = RTL_PATH.io_diffCommits_info_138_vecWen; \
        force U_IF_NAME.io_diffCommits_info_138_v0Wen = RTL_PATH.io_diffCommits_info_138_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_138_vlWen = RTL_PATH.io_diffCommits_info_138_vlWen; \
        force U_IF_NAME.io_diffCommits_info_139_ldest = RTL_PATH.io_diffCommits_info_139_ldest; \
        force U_IF_NAME.io_diffCommits_info_139_pdest = RTL_PATH.io_diffCommits_info_139_pdest; \
        force U_IF_NAME.io_diffCommits_info_139_rfWen = RTL_PATH.io_diffCommits_info_139_rfWen; \
        force U_IF_NAME.io_diffCommits_info_139_fpWen = RTL_PATH.io_diffCommits_info_139_fpWen; \
        force U_IF_NAME.io_diffCommits_info_139_vecWen = RTL_PATH.io_diffCommits_info_139_vecWen; \
        force U_IF_NAME.io_diffCommits_info_139_v0Wen = RTL_PATH.io_diffCommits_info_139_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_139_vlWen = RTL_PATH.io_diffCommits_info_139_vlWen; \
        force U_IF_NAME.io_diffCommits_info_140_ldest = RTL_PATH.io_diffCommits_info_140_ldest; \
        force U_IF_NAME.io_diffCommits_info_140_pdest = RTL_PATH.io_diffCommits_info_140_pdest; \
        force U_IF_NAME.io_diffCommits_info_140_rfWen = RTL_PATH.io_diffCommits_info_140_rfWen; \
        force U_IF_NAME.io_diffCommits_info_140_fpWen = RTL_PATH.io_diffCommits_info_140_fpWen; \
        force U_IF_NAME.io_diffCommits_info_140_vecWen = RTL_PATH.io_diffCommits_info_140_vecWen; \
        force U_IF_NAME.io_diffCommits_info_140_v0Wen = RTL_PATH.io_diffCommits_info_140_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_140_vlWen = RTL_PATH.io_diffCommits_info_140_vlWen; \
        force U_IF_NAME.io_diffCommits_info_141_ldest = RTL_PATH.io_diffCommits_info_141_ldest; \
        force U_IF_NAME.io_diffCommits_info_141_pdest = RTL_PATH.io_diffCommits_info_141_pdest; \
        force U_IF_NAME.io_diffCommits_info_141_rfWen = RTL_PATH.io_diffCommits_info_141_rfWen; \
        force U_IF_NAME.io_diffCommits_info_141_fpWen = RTL_PATH.io_diffCommits_info_141_fpWen; \
        force U_IF_NAME.io_diffCommits_info_141_vecWen = RTL_PATH.io_diffCommits_info_141_vecWen; \
        force U_IF_NAME.io_diffCommits_info_141_v0Wen = RTL_PATH.io_diffCommits_info_141_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_141_vlWen = RTL_PATH.io_diffCommits_info_141_vlWen; \
        force U_IF_NAME.io_diffCommits_info_142_ldest = RTL_PATH.io_diffCommits_info_142_ldest; \
        force U_IF_NAME.io_diffCommits_info_142_pdest = RTL_PATH.io_diffCommits_info_142_pdest; \
        force U_IF_NAME.io_diffCommits_info_142_rfWen = RTL_PATH.io_diffCommits_info_142_rfWen; \
        force U_IF_NAME.io_diffCommits_info_142_fpWen = RTL_PATH.io_diffCommits_info_142_fpWen; \
        force U_IF_NAME.io_diffCommits_info_142_vecWen = RTL_PATH.io_diffCommits_info_142_vecWen; \
        force U_IF_NAME.io_diffCommits_info_142_v0Wen = RTL_PATH.io_diffCommits_info_142_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_142_vlWen = RTL_PATH.io_diffCommits_info_142_vlWen; \
        force U_IF_NAME.io_diffCommits_info_143_ldest = RTL_PATH.io_diffCommits_info_143_ldest; \
        force U_IF_NAME.io_diffCommits_info_143_pdest = RTL_PATH.io_diffCommits_info_143_pdest; \
        force U_IF_NAME.io_diffCommits_info_143_rfWen = RTL_PATH.io_diffCommits_info_143_rfWen; \
        force U_IF_NAME.io_diffCommits_info_143_fpWen = RTL_PATH.io_diffCommits_info_143_fpWen; \
        force U_IF_NAME.io_diffCommits_info_143_vecWen = RTL_PATH.io_diffCommits_info_143_vecWen; \
        force U_IF_NAME.io_diffCommits_info_143_v0Wen = RTL_PATH.io_diffCommits_info_143_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_143_vlWen = RTL_PATH.io_diffCommits_info_143_vlWen; \
        force U_IF_NAME.io_diffCommits_info_144_ldest = RTL_PATH.io_diffCommits_info_144_ldest; \
        force U_IF_NAME.io_diffCommits_info_144_pdest = RTL_PATH.io_diffCommits_info_144_pdest; \
        force U_IF_NAME.io_diffCommits_info_144_rfWen = RTL_PATH.io_diffCommits_info_144_rfWen; \
        force U_IF_NAME.io_diffCommits_info_144_fpWen = RTL_PATH.io_diffCommits_info_144_fpWen; \
        force U_IF_NAME.io_diffCommits_info_144_vecWen = RTL_PATH.io_diffCommits_info_144_vecWen; \
        force U_IF_NAME.io_diffCommits_info_144_v0Wen = RTL_PATH.io_diffCommits_info_144_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_144_vlWen = RTL_PATH.io_diffCommits_info_144_vlWen; \
        force U_IF_NAME.io_diffCommits_info_145_ldest = RTL_PATH.io_diffCommits_info_145_ldest; \
        force U_IF_NAME.io_diffCommits_info_145_pdest = RTL_PATH.io_diffCommits_info_145_pdest; \
        force U_IF_NAME.io_diffCommits_info_145_rfWen = RTL_PATH.io_diffCommits_info_145_rfWen; \
        force U_IF_NAME.io_diffCommits_info_145_fpWen = RTL_PATH.io_diffCommits_info_145_fpWen; \
        force U_IF_NAME.io_diffCommits_info_145_vecWen = RTL_PATH.io_diffCommits_info_145_vecWen; \
        force U_IF_NAME.io_diffCommits_info_145_v0Wen = RTL_PATH.io_diffCommits_info_145_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_145_vlWen = RTL_PATH.io_diffCommits_info_145_vlWen; \
        force U_IF_NAME.io_diffCommits_info_146_ldest = RTL_PATH.io_diffCommits_info_146_ldest; \
        force U_IF_NAME.io_diffCommits_info_146_pdest = RTL_PATH.io_diffCommits_info_146_pdest; \
        force U_IF_NAME.io_diffCommits_info_146_rfWen = RTL_PATH.io_diffCommits_info_146_rfWen; \
        force U_IF_NAME.io_diffCommits_info_146_fpWen = RTL_PATH.io_diffCommits_info_146_fpWen; \
        force U_IF_NAME.io_diffCommits_info_146_vecWen = RTL_PATH.io_diffCommits_info_146_vecWen; \
        force U_IF_NAME.io_diffCommits_info_146_v0Wen = RTL_PATH.io_diffCommits_info_146_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_146_vlWen = RTL_PATH.io_diffCommits_info_146_vlWen; \
        force U_IF_NAME.io_diffCommits_info_147_ldest = RTL_PATH.io_diffCommits_info_147_ldest; \
        force U_IF_NAME.io_diffCommits_info_147_pdest = RTL_PATH.io_diffCommits_info_147_pdest; \
        force U_IF_NAME.io_diffCommits_info_147_rfWen = RTL_PATH.io_diffCommits_info_147_rfWen; \
        force U_IF_NAME.io_diffCommits_info_147_fpWen = RTL_PATH.io_diffCommits_info_147_fpWen; \
        force U_IF_NAME.io_diffCommits_info_147_vecWen = RTL_PATH.io_diffCommits_info_147_vecWen; \
        force U_IF_NAME.io_diffCommits_info_147_v0Wen = RTL_PATH.io_diffCommits_info_147_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_147_vlWen = RTL_PATH.io_diffCommits_info_147_vlWen; \
        force U_IF_NAME.io_diffCommits_info_148_ldest = RTL_PATH.io_diffCommits_info_148_ldest; \
        force U_IF_NAME.io_diffCommits_info_148_pdest = RTL_PATH.io_diffCommits_info_148_pdest; \
        force U_IF_NAME.io_diffCommits_info_148_rfWen = RTL_PATH.io_diffCommits_info_148_rfWen; \
        force U_IF_NAME.io_diffCommits_info_148_fpWen = RTL_PATH.io_diffCommits_info_148_fpWen; \
        force U_IF_NAME.io_diffCommits_info_148_vecWen = RTL_PATH.io_diffCommits_info_148_vecWen; \
        force U_IF_NAME.io_diffCommits_info_148_v0Wen = RTL_PATH.io_diffCommits_info_148_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_148_vlWen = RTL_PATH.io_diffCommits_info_148_vlWen; \
        force U_IF_NAME.io_diffCommits_info_149_ldest = RTL_PATH.io_diffCommits_info_149_ldest; \
        force U_IF_NAME.io_diffCommits_info_149_pdest = RTL_PATH.io_diffCommits_info_149_pdest; \
        force U_IF_NAME.io_diffCommits_info_149_rfWen = RTL_PATH.io_diffCommits_info_149_rfWen; \
        force U_IF_NAME.io_diffCommits_info_149_fpWen = RTL_PATH.io_diffCommits_info_149_fpWen; \
        force U_IF_NAME.io_diffCommits_info_149_vecWen = RTL_PATH.io_diffCommits_info_149_vecWen; \
        force U_IF_NAME.io_diffCommits_info_149_v0Wen = RTL_PATH.io_diffCommits_info_149_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_149_vlWen = RTL_PATH.io_diffCommits_info_149_vlWen; \
        force U_IF_NAME.io_diffCommits_info_150_ldest = RTL_PATH.io_diffCommits_info_150_ldest; \
        force U_IF_NAME.io_diffCommits_info_150_pdest = RTL_PATH.io_diffCommits_info_150_pdest; \
        force U_IF_NAME.io_diffCommits_info_150_rfWen = RTL_PATH.io_diffCommits_info_150_rfWen; \
        force U_IF_NAME.io_diffCommits_info_150_fpWen = RTL_PATH.io_diffCommits_info_150_fpWen; \
        force U_IF_NAME.io_diffCommits_info_150_vecWen = RTL_PATH.io_diffCommits_info_150_vecWen; \
        force U_IF_NAME.io_diffCommits_info_150_v0Wen = RTL_PATH.io_diffCommits_info_150_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_150_vlWen = RTL_PATH.io_diffCommits_info_150_vlWen; \
        force U_IF_NAME.io_diffCommits_info_151_ldest = RTL_PATH.io_diffCommits_info_151_ldest; \
        force U_IF_NAME.io_diffCommits_info_151_pdest = RTL_PATH.io_diffCommits_info_151_pdest; \
        force U_IF_NAME.io_diffCommits_info_151_rfWen = RTL_PATH.io_diffCommits_info_151_rfWen; \
        force U_IF_NAME.io_diffCommits_info_151_fpWen = RTL_PATH.io_diffCommits_info_151_fpWen; \
        force U_IF_NAME.io_diffCommits_info_151_vecWen = RTL_PATH.io_diffCommits_info_151_vecWen; \
        force U_IF_NAME.io_diffCommits_info_151_v0Wen = RTL_PATH.io_diffCommits_info_151_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_151_vlWen = RTL_PATH.io_diffCommits_info_151_vlWen; \
        force U_IF_NAME.io_diffCommits_info_152_ldest = RTL_PATH.io_diffCommits_info_152_ldest; \
        force U_IF_NAME.io_diffCommits_info_152_pdest = RTL_PATH.io_diffCommits_info_152_pdest; \
        force U_IF_NAME.io_diffCommits_info_152_rfWen = RTL_PATH.io_diffCommits_info_152_rfWen; \
        force U_IF_NAME.io_diffCommits_info_152_fpWen = RTL_PATH.io_diffCommits_info_152_fpWen; \
        force U_IF_NAME.io_diffCommits_info_152_vecWen = RTL_PATH.io_diffCommits_info_152_vecWen; \
        force U_IF_NAME.io_diffCommits_info_152_v0Wen = RTL_PATH.io_diffCommits_info_152_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_152_vlWen = RTL_PATH.io_diffCommits_info_152_vlWen; \
        force U_IF_NAME.io_diffCommits_info_153_ldest = RTL_PATH.io_diffCommits_info_153_ldest; \
        force U_IF_NAME.io_diffCommits_info_153_pdest = RTL_PATH.io_diffCommits_info_153_pdest; \
        force U_IF_NAME.io_diffCommits_info_153_rfWen = RTL_PATH.io_diffCommits_info_153_rfWen; \
        force U_IF_NAME.io_diffCommits_info_153_fpWen = RTL_PATH.io_diffCommits_info_153_fpWen; \
        force U_IF_NAME.io_diffCommits_info_153_vecWen = RTL_PATH.io_diffCommits_info_153_vecWen; \
        force U_IF_NAME.io_diffCommits_info_153_v0Wen = RTL_PATH.io_diffCommits_info_153_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_153_vlWen = RTL_PATH.io_diffCommits_info_153_vlWen; \
        force U_IF_NAME.io_diffCommits_info_154_ldest = RTL_PATH.io_diffCommits_info_154_ldest; \
        force U_IF_NAME.io_diffCommits_info_154_pdest = RTL_PATH.io_diffCommits_info_154_pdest; \
        force U_IF_NAME.io_diffCommits_info_154_rfWen = RTL_PATH.io_diffCommits_info_154_rfWen; \
        force U_IF_NAME.io_diffCommits_info_154_fpWen = RTL_PATH.io_diffCommits_info_154_fpWen; \
        force U_IF_NAME.io_diffCommits_info_154_vecWen = RTL_PATH.io_diffCommits_info_154_vecWen; \
        force U_IF_NAME.io_diffCommits_info_154_v0Wen = RTL_PATH.io_diffCommits_info_154_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_154_vlWen = RTL_PATH.io_diffCommits_info_154_vlWen; \
        force U_IF_NAME.io_diffCommits_info_155_ldest = RTL_PATH.io_diffCommits_info_155_ldest; \
        force U_IF_NAME.io_diffCommits_info_155_pdest = RTL_PATH.io_diffCommits_info_155_pdest; \
        force U_IF_NAME.io_diffCommits_info_155_rfWen = RTL_PATH.io_diffCommits_info_155_rfWen; \
        force U_IF_NAME.io_diffCommits_info_155_fpWen = RTL_PATH.io_diffCommits_info_155_fpWen; \
        force U_IF_NAME.io_diffCommits_info_155_vecWen = RTL_PATH.io_diffCommits_info_155_vecWen; \
        force U_IF_NAME.io_diffCommits_info_155_v0Wen = RTL_PATH.io_diffCommits_info_155_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_155_vlWen = RTL_PATH.io_diffCommits_info_155_vlWen; \
        force U_IF_NAME.io_diffCommits_info_156_ldest = RTL_PATH.io_diffCommits_info_156_ldest; \
        force U_IF_NAME.io_diffCommits_info_156_pdest = RTL_PATH.io_diffCommits_info_156_pdest; \
        force U_IF_NAME.io_diffCommits_info_156_rfWen = RTL_PATH.io_diffCommits_info_156_rfWen; \
        force U_IF_NAME.io_diffCommits_info_156_fpWen = RTL_PATH.io_diffCommits_info_156_fpWen; \
        force U_IF_NAME.io_diffCommits_info_156_vecWen = RTL_PATH.io_diffCommits_info_156_vecWen; \
        force U_IF_NAME.io_diffCommits_info_156_v0Wen = RTL_PATH.io_diffCommits_info_156_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_156_vlWen = RTL_PATH.io_diffCommits_info_156_vlWen; \
        force U_IF_NAME.io_diffCommits_info_157_ldest = RTL_PATH.io_diffCommits_info_157_ldest; \
        force U_IF_NAME.io_diffCommits_info_157_pdest = RTL_PATH.io_diffCommits_info_157_pdest; \
        force U_IF_NAME.io_diffCommits_info_157_rfWen = RTL_PATH.io_diffCommits_info_157_rfWen; \
        force U_IF_NAME.io_diffCommits_info_157_fpWen = RTL_PATH.io_diffCommits_info_157_fpWen; \
        force U_IF_NAME.io_diffCommits_info_157_vecWen = RTL_PATH.io_diffCommits_info_157_vecWen; \
        force U_IF_NAME.io_diffCommits_info_157_v0Wen = RTL_PATH.io_diffCommits_info_157_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_157_vlWen = RTL_PATH.io_diffCommits_info_157_vlWen; \
        force U_IF_NAME.io_diffCommits_info_158_ldest = RTL_PATH.io_diffCommits_info_158_ldest; \
        force U_IF_NAME.io_diffCommits_info_158_pdest = RTL_PATH.io_diffCommits_info_158_pdest; \
        force U_IF_NAME.io_diffCommits_info_158_rfWen = RTL_PATH.io_diffCommits_info_158_rfWen; \
        force U_IF_NAME.io_diffCommits_info_158_fpWen = RTL_PATH.io_diffCommits_info_158_fpWen; \
        force U_IF_NAME.io_diffCommits_info_158_vecWen = RTL_PATH.io_diffCommits_info_158_vecWen; \
        force U_IF_NAME.io_diffCommits_info_158_v0Wen = RTL_PATH.io_diffCommits_info_158_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_158_vlWen = RTL_PATH.io_diffCommits_info_158_vlWen; \
        force U_IF_NAME.io_diffCommits_info_159_ldest = RTL_PATH.io_diffCommits_info_159_ldest; \
        force U_IF_NAME.io_diffCommits_info_159_pdest = RTL_PATH.io_diffCommits_info_159_pdest; \
        force U_IF_NAME.io_diffCommits_info_159_rfWen = RTL_PATH.io_diffCommits_info_159_rfWen; \
        force U_IF_NAME.io_diffCommits_info_159_fpWen = RTL_PATH.io_diffCommits_info_159_fpWen; \
        force U_IF_NAME.io_diffCommits_info_159_vecWen = RTL_PATH.io_diffCommits_info_159_vecWen; \
        force U_IF_NAME.io_diffCommits_info_159_v0Wen = RTL_PATH.io_diffCommits_info_159_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_159_vlWen = RTL_PATH.io_diffCommits_info_159_vlWen; \
        force U_IF_NAME.io_diffCommits_info_160_ldest = RTL_PATH.io_diffCommits_info_160_ldest; \
        force U_IF_NAME.io_diffCommits_info_160_pdest = RTL_PATH.io_diffCommits_info_160_pdest; \
        force U_IF_NAME.io_diffCommits_info_160_rfWen = RTL_PATH.io_diffCommits_info_160_rfWen; \
        force U_IF_NAME.io_diffCommits_info_160_fpWen = RTL_PATH.io_diffCommits_info_160_fpWen; \
        force U_IF_NAME.io_diffCommits_info_160_vecWen = RTL_PATH.io_diffCommits_info_160_vecWen; \
        force U_IF_NAME.io_diffCommits_info_160_v0Wen = RTL_PATH.io_diffCommits_info_160_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_160_vlWen = RTL_PATH.io_diffCommits_info_160_vlWen; \
        force U_IF_NAME.io_diffCommits_info_161_ldest = RTL_PATH.io_diffCommits_info_161_ldest; \
        force U_IF_NAME.io_diffCommits_info_161_pdest = RTL_PATH.io_diffCommits_info_161_pdest; \
        force U_IF_NAME.io_diffCommits_info_161_rfWen = RTL_PATH.io_diffCommits_info_161_rfWen; \
        force U_IF_NAME.io_diffCommits_info_161_fpWen = RTL_PATH.io_diffCommits_info_161_fpWen; \
        force U_IF_NAME.io_diffCommits_info_161_vecWen = RTL_PATH.io_diffCommits_info_161_vecWen; \
        force U_IF_NAME.io_diffCommits_info_161_v0Wen = RTL_PATH.io_diffCommits_info_161_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_161_vlWen = RTL_PATH.io_diffCommits_info_161_vlWen; \
        force U_IF_NAME.io_diffCommits_info_162_ldest = RTL_PATH.io_diffCommits_info_162_ldest; \
        force U_IF_NAME.io_diffCommits_info_162_pdest = RTL_PATH.io_diffCommits_info_162_pdest; \
        force U_IF_NAME.io_diffCommits_info_162_rfWen = RTL_PATH.io_diffCommits_info_162_rfWen; \
        force U_IF_NAME.io_diffCommits_info_162_fpWen = RTL_PATH.io_diffCommits_info_162_fpWen; \
        force U_IF_NAME.io_diffCommits_info_162_vecWen = RTL_PATH.io_diffCommits_info_162_vecWen; \
        force U_IF_NAME.io_diffCommits_info_162_v0Wen = RTL_PATH.io_diffCommits_info_162_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_162_vlWen = RTL_PATH.io_diffCommits_info_162_vlWen; \
        force U_IF_NAME.io_diffCommits_info_163_ldest = RTL_PATH.io_diffCommits_info_163_ldest; \
        force U_IF_NAME.io_diffCommits_info_163_pdest = RTL_PATH.io_diffCommits_info_163_pdest; \
        force U_IF_NAME.io_diffCommits_info_163_rfWen = RTL_PATH.io_diffCommits_info_163_rfWen; \
        force U_IF_NAME.io_diffCommits_info_163_fpWen = RTL_PATH.io_diffCommits_info_163_fpWen; \
        force U_IF_NAME.io_diffCommits_info_163_vecWen = RTL_PATH.io_diffCommits_info_163_vecWen; \
        force U_IF_NAME.io_diffCommits_info_163_v0Wen = RTL_PATH.io_diffCommits_info_163_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_163_vlWen = RTL_PATH.io_diffCommits_info_163_vlWen; \
        force U_IF_NAME.io_diffCommits_info_164_ldest = RTL_PATH.io_diffCommits_info_164_ldest; \
        force U_IF_NAME.io_diffCommits_info_164_pdest = RTL_PATH.io_diffCommits_info_164_pdest; \
        force U_IF_NAME.io_diffCommits_info_164_rfWen = RTL_PATH.io_diffCommits_info_164_rfWen; \
        force U_IF_NAME.io_diffCommits_info_164_fpWen = RTL_PATH.io_diffCommits_info_164_fpWen; \
        force U_IF_NAME.io_diffCommits_info_164_vecWen = RTL_PATH.io_diffCommits_info_164_vecWen; \
        force U_IF_NAME.io_diffCommits_info_164_v0Wen = RTL_PATH.io_diffCommits_info_164_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_164_vlWen = RTL_PATH.io_diffCommits_info_164_vlWen; \
        force U_IF_NAME.io_diffCommits_info_165_ldest = RTL_PATH.io_diffCommits_info_165_ldest; \
        force U_IF_NAME.io_diffCommits_info_165_pdest = RTL_PATH.io_diffCommits_info_165_pdest; \
        force U_IF_NAME.io_diffCommits_info_165_rfWen = RTL_PATH.io_diffCommits_info_165_rfWen; \
        force U_IF_NAME.io_diffCommits_info_165_fpWen = RTL_PATH.io_diffCommits_info_165_fpWen; \
        force U_IF_NAME.io_diffCommits_info_165_vecWen = RTL_PATH.io_diffCommits_info_165_vecWen; \
        force U_IF_NAME.io_diffCommits_info_165_v0Wen = RTL_PATH.io_diffCommits_info_165_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_165_vlWen = RTL_PATH.io_diffCommits_info_165_vlWen; \
        force U_IF_NAME.io_diffCommits_info_166_ldest = RTL_PATH.io_diffCommits_info_166_ldest; \
        force U_IF_NAME.io_diffCommits_info_166_pdest = RTL_PATH.io_diffCommits_info_166_pdest; \
        force U_IF_NAME.io_diffCommits_info_166_rfWen = RTL_PATH.io_diffCommits_info_166_rfWen; \
        force U_IF_NAME.io_diffCommits_info_166_fpWen = RTL_PATH.io_diffCommits_info_166_fpWen; \
        force U_IF_NAME.io_diffCommits_info_166_vecWen = RTL_PATH.io_diffCommits_info_166_vecWen; \
        force U_IF_NAME.io_diffCommits_info_166_v0Wen = RTL_PATH.io_diffCommits_info_166_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_166_vlWen = RTL_PATH.io_diffCommits_info_166_vlWen; \
        force U_IF_NAME.io_diffCommits_info_167_ldest = RTL_PATH.io_diffCommits_info_167_ldest; \
        force U_IF_NAME.io_diffCommits_info_167_pdest = RTL_PATH.io_diffCommits_info_167_pdest; \
        force U_IF_NAME.io_diffCommits_info_167_rfWen = RTL_PATH.io_diffCommits_info_167_rfWen; \
        force U_IF_NAME.io_diffCommits_info_167_fpWen = RTL_PATH.io_diffCommits_info_167_fpWen; \
        force U_IF_NAME.io_diffCommits_info_167_vecWen = RTL_PATH.io_diffCommits_info_167_vecWen; \
        force U_IF_NAME.io_diffCommits_info_167_v0Wen = RTL_PATH.io_diffCommits_info_167_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_167_vlWen = RTL_PATH.io_diffCommits_info_167_vlWen; \
        force U_IF_NAME.io_diffCommits_info_168_ldest = RTL_PATH.io_diffCommits_info_168_ldest; \
        force U_IF_NAME.io_diffCommits_info_168_pdest = RTL_PATH.io_diffCommits_info_168_pdest; \
        force U_IF_NAME.io_diffCommits_info_168_rfWen = RTL_PATH.io_diffCommits_info_168_rfWen; \
        force U_IF_NAME.io_diffCommits_info_168_fpWen = RTL_PATH.io_diffCommits_info_168_fpWen; \
        force U_IF_NAME.io_diffCommits_info_168_vecWen = RTL_PATH.io_diffCommits_info_168_vecWen; \
        force U_IF_NAME.io_diffCommits_info_168_v0Wen = RTL_PATH.io_diffCommits_info_168_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_168_vlWen = RTL_PATH.io_diffCommits_info_168_vlWen; \
        force U_IF_NAME.io_diffCommits_info_169_ldest = RTL_PATH.io_diffCommits_info_169_ldest; \
        force U_IF_NAME.io_diffCommits_info_169_pdest = RTL_PATH.io_diffCommits_info_169_pdest; \
        force U_IF_NAME.io_diffCommits_info_169_rfWen = RTL_PATH.io_diffCommits_info_169_rfWen; \
        force U_IF_NAME.io_diffCommits_info_169_fpWen = RTL_PATH.io_diffCommits_info_169_fpWen; \
        force U_IF_NAME.io_diffCommits_info_169_vecWen = RTL_PATH.io_diffCommits_info_169_vecWen; \
        force U_IF_NAME.io_diffCommits_info_169_v0Wen = RTL_PATH.io_diffCommits_info_169_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_169_vlWen = RTL_PATH.io_diffCommits_info_169_vlWen; \
        force U_IF_NAME.io_diffCommits_info_170_ldest = RTL_PATH.io_diffCommits_info_170_ldest; \
        force U_IF_NAME.io_diffCommits_info_170_pdest = RTL_PATH.io_diffCommits_info_170_pdest; \
        force U_IF_NAME.io_diffCommits_info_170_rfWen = RTL_PATH.io_diffCommits_info_170_rfWen; \
        force U_IF_NAME.io_diffCommits_info_170_fpWen = RTL_PATH.io_diffCommits_info_170_fpWen; \
        force U_IF_NAME.io_diffCommits_info_170_vecWen = RTL_PATH.io_diffCommits_info_170_vecWen; \
        force U_IF_NAME.io_diffCommits_info_170_v0Wen = RTL_PATH.io_diffCommits_info_170_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_170_vlWen = RTL_PATH.io_diffCommits_info_170_vlWen; \
        force U_IF_NAME.io_diffCommits_info_171_ldest = RTL_PATH.io_diffCommits_info_171_ldest; \
        force U_IF_NAME.io_diffCommits_info_171_pdest = RTL_PATH.io_diffCommits_info_171_pdest; \
        force U_IF_NAME.io_diffCommits_info_171_rfWen = RTL_PATH.io_diffCommits_info_171_rfWen; \
        force U_IF_NAME.io_diffCommits_info_171_fpWen = RTL_PATH.io_diffCommits_info_171_fpWen; \
        force U_IF_NAME.io_diffCommits_info_171_vecWen = RTL_PATH.io_diffCommits_info_171_vecWen; \
        force U_IF_NAME.io_diffCommits_info_171_v0Wen = RTL_PATH.io_diffCommits_info_171_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_171_vlWen = RTL_PATH.io_diffCommits_info_171_vlWen; \
        force U_IF_NAME.io_diffCommits_info_172_ldest = RTL_PATH.io_diffCommits_info_172_ldest; \
        force U_IF_NAME.io_diffCommits_info_172_pdest = RTL_PATH.io_diffCommits_info_172_pdest; \
        force U_IF_NAME.io_diffCommits_info_172_rfWen = RTL_PATH.io_diffCommits_info_172_rfWen; \
        force U_IF_NAME.io_diffCommits_info_172_fpWen = RTL_PATH.io_diffCommits_info_172_fpWen; \
        force U_IF_NAME.io_diffCommits_info_172_vecWen = RTL_PATH.io_diffCommits_info_172_vecWen; \
        force U_IF_NAME.io_diffCommits_info_172_v0Wen = RTL_PATH.io_diffCommits_info_172_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_172_vlWen = RTL_PATH.io_diffCommits_info_172_vlWen; \
        force U_IF_NAME.io_diffCommits_info_173_ldest = RTL_PATH.io_diffCommits_info_173_ldest; \
        force U_IF_NAME.io_diffCommits_info_173_pdest = RTL_PATH.io_diffCommits_info_173_pdest; \
        force U_IF_NAME.io_diffCommits_info_173_rfWen = RTL_PATH.io_diffCommits_info_173_rfWen; \
        force U_IF_NAME.io_diffCommits_info_173_fpWen = RTL_PATH.io_diffCommits_info_173_fpWen; \
        force U_IF_NAME.io_diffCommits_info_173_vecWen = RTL_PATH.io_diffCommits_info_173_vecWen; \
        force U_IF_NAME.io_diffCommits_info_173_v0Wen = RTL_PATH.io_diffCommits_info_173_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_173_vlWen = RTL_PATH.io_diffCommits_info_173_vlWen; \
        force U_IF_NAME.io_diffCommits_info_174_ldest = RTL_PATH.io_diffCommits_info_174_ldest; \
        force U_IF_NAME.io_diffCommits_info_174_pdest = RTL_PATH.io_diffCommits_info_174_pdest; \
        force U_IF_NAME.io_diffCommits_info_174_rfWen = RTL_PATH.io_diffCommits_info_174_rfWen; \
        force U_IF_NAME.io_diffCommits_info_174_fpWen = RTL_PATH.io_diffCommits_info_174_fpWen; \
        force U_IF_NAME.io_diffCommits_info_174_vecWen = RTL_PATH.io_diffCommits_info_174_vecWen; \
        force U_IF_NAME.io_diffCommits_info_174_v0Wen = RTL_PATH.io_diffCommits_info_174_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_174_vlWen = RTL_PATH.io_diffCommits_info_174_vlWen; \
        force U_IF_NAME.io_diffCommits_info_175_ldest = RTL_PATH.io_diffCommits_info_175_ldest; \
        force U_IF_NAME.io_diffCommits_info_175_pdest = RTL_PATH.io_diffCommits_info_175_pdest; \
        force U_IF_NAME.io_diffCommits_info_175_rfWen = RTL_PATH.io_diffCommits_info_175_rfWen; \
        force U_IF_NAME.io_diffCommits_info_175_fpWen = RTL_PATH.io_diffCommits_info_175_fpWen; \
        force U_IF_NAME.io_diffCommits_info_175_vecWen = RTL_PATH.io_diffCommits_info_175_vecWen; \
        force U_IF_NAME.io_diffCommits_info_175_v0Wen = RTL_PATH.io_diffCommits_info_175_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_175_vlWen = RTL_PATH.io_diffCommits_info_175_vlWen; \
        force U_IF_NAME.io_diffCommits_info_176_ldest = RTL_PATH.io_diffCommits_info_176_ldest; \
        force U_IF_NAME.io_diffCommits_info_176_pdest = RTL_PATH.io_diffCommits_info_176_pdest; \
        force U_IF_NAME.io_diffCommits_info_176_rfWen = RTL_PATH.io_diffCommits_info_176_rfWen; \
        force U_IF_NAME.io_diffCommits_info_176_fpWen = RTL_PATH.io_diffCommits_info_176_fpWen; \
        force U_IF_NAME.io_diffCommits_info_176_vecWen = RTL_PATH.io_diffCommits_info_176_vecWen; \
        force U_IF_NAME.io_diffCommits_info_176_v0Wen = RTL_PATH.io_diffCommits_info_176_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_176_vlWen = RTL_PATH.io_diffCommits_info_176_vlWen; \
        force U_IF_NAME.io_diffCommits_info_177_ldest = RTL_PATH.io_diffCommits_info_177_ldest; \
        force U_IF_NAME.io_diffCommits_info_177_pdest = RTL_PATH.io_diffCommits_info_177_pdest; \
        force U_IF_NAME.io_diffCommits_info_177_rfWen = RTL_PATH.io_diffCommits_info_177_rfWen; \
        force U_IF_NAME.io_diffCommits_info_177_fpWen = RTL_PATH.io_diffCommits_info_177_fpWen; \
        force U_IF_NAME.io_diffCommits_info_177_vecWen = RTL_PATH.io_diffCommits_info_177_vecWen; \
        force U_IF_NAME.io_diffCommits_info_177_v0Wen = RTL_PATH.io_diffCommits_info_177_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_177_vlWen = RTL_PATH.io_diffCommits_info_177_vlWen; \
        force U_IF_NAME.io_diffCommits_info_178_ldest = RTL_PATH.io_diffCommits_info_178_ldest; \
        force U_IF_NAME.io_diffCommits_info_178_pdest = RTL_PATH.io_diffCommits_info_178_pdest; \
        force U_IF_NAME.io_diffCommits_info_178_rfWen = RTL_PATH.io_diffCommits_info_178_rfWen; \
        force U_IF_NAME.io_diffCommits_info_178_fpWen = RTL_PATH.io_diffCommits_info_178_fpWen; \
        force U_IF_NAME.io_diffCommits_info_178_vecWen = RTL_PATH.io_diffCommits_info_178_vecWen; \
        force U_IF_NAME.io_diffCommits_info_178_v0Wen = RTL_PATH.io_diffCommits_info_178_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_178_vlWen = RTL_PATH.io_diffCommits_info_178_vlWen; \
        force U_IF_NAME.io_diffCommits_info_179_ldest = RTL_PATH.io_diffCommits_info_179_ldest; \
        force U_IF_NAME.io_diffCommits_info_179_pdest = RTL_PATH.io_diffCommits_info_179_pdest; \
        force U_IF_NAME.io_diffCommits_info_179_rfWen = RTL_PATH.io_diffCommits_info_179_rfWen; \
        force U_IF_NAME.io_diffCommits_info_179_fpWen = RTL_PATH.io_diffCommits_info_179_fpWen; \
        force U_IF_NAME.io_diffCommits_info_179_vecWen = RTL_PATH.io_diffCommits_info_179_vecWen; \
        force U_IF_NAME.io_diffCommits_info_179_v0Wen = RTL_PATH.io_diffCommits_info_179_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_179_vlWen = RTL_PATH.io_diffCommits_info_179_vlWen; \
        force U_IF_NAME.io_diffCommits_info_180_ldest = RTL_PATH.io_diffCommits_info_180_ldest; \
        force U_IF_NAME.io_diffCommits_info_180_pdest = RTL_PATH.io_diffCommits_info_180_pdest; \
        force U_IF_NAME.io_diffCommits_info_180_rfWen = RTL_PATH.io_diffCommits_info_180_rfWen; \
        force U_IF_NAME.io_diffCommits_info_180_fpWen = RTL_PATH.io_diffCommits_info_180_fpWen; \
        force U_IF_NAME.io_diffCommits_info_180_vecWen = RTL_PATH.io_diffCommits_info_180_vecWen; \
        force U_IF_NAME.io_diffCommits_info_180_v0Wen = RTL_PATH.io_diffCommits_info_180_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_180_vlWen = RTL_PATH.io_diffCommits_info_180_vlWen; \
        force U_IF_NAME.io_diffCommits_info_181_ldest = RTL_PATH.io_diffCommits_info_181_ldest; \
        force U_IF_NAME.io_diffCommits_info_181_pdest = RTL_PATH.io_diffCommits_info_181_pdest; \
        force U_IF_NAME.io_diffCommits_info_181_rfWen = RTL_PATH.io_diffCommits_info_181_rfWen; \
        force U_IF_NAME.io_diffCommits_info_181_fpWen = RTL_PATH.io_diffCommits_info_181_fpWen; \
        force U_IF_NAME.io_diffCommits_info_181_vecWen = RTL_PATH.io_diffCommits_info_181_vecWen; \
        force U_IF_NAME.io_diffCommits_info_181_v0Wen = RTL_PATH.io_diffCommits_info_181_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_181_vlWen = RTL_PATH.io_diffCommits_info_181_vlWen; \
        force U_IF_NAME.io_diffCommits_info_182_ldest = RTL_PATH.io_diffCommits_info_182_ldest; \
        force U_IF_NAME.io_diffCommits_info_182_pdest = RTL_PATH.io_diffCommits_info_182_pdest; \
        force U_IF_NAME.io_diffCommits_info_182_rfWen = RTL_PATH.io_diffCommits_info_182_rfWen; \
        force U_IF_NAME.io_diffCommits_info_182_fpWen = RTL_PATH.io_diffCommits_info_182_fpWen; \
        force U_IF_NAME.io_diffCommits_info_182_vecWen = RTL_PATH.io_diffCommits_info_182_vecWen; \
        force U_IF_NAME.io_diffCommits_info_182_v0Wen = RTL_PATH.io_diffCommits_info_182_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_182_vlWen = RTL_PATH.io_diffCommits_info_182_vlWen; \
        force U_IF_NAME.io_diffCommits_info_183_ldest = RTL_PATH.io_diffCommits_info_183_ldest; \
        force U_IF_NAME.io_diffCommits_info_183_pdest = RTL_PATH.io_diffCommits_info_183_pdest; \
        force U_IF_NAME.io_diffCommits_info_183_rfWen = RTL_PATH.io_diffCommits_info_183_rfWen; \
        force U_IF_NAME.io_diffCommits_info_183_fpWen = RTL_PATH.io_diffCommits_info_183_fpWen; \
        force U_IF_NAME.io_diffCommits_info_183_vecWen = RTL_PATH.io_diffCommits_info_183_vecWen; \
        force U_IF_NAME.io_diffCommits_info_183_v0Wen = RTL_PATH.io_diffCommits_info_183_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_183_vlWen = RTL_PATH.io_diffCommits_info_183_vlWen; \
        force U_IF_NAME.io_diffCommits_info_184_ldest = RTL_PATH.io_diffCommits_info_184_ldest; \
        force U_IF_NAME.io_diffCommits_info_184_pdest = RTL_PATH.io_diffCommits_info_184_pdest; \
        force U_IF_NAME.io_diffCommits_info_184_rfWen = RTL_PATH.io_diffCommits_info_184_rfWen; \
        force U_IF_NAME.io_diffCommits_info_184_fpWen = RTL_PATH.io_diffCommits_info_184_fpWen; \
        force U_IF_NAME.io_diffCommits_info_184_vecWen = RTL_PATH.io_diffCommits_info_184_vecWen; \
        force U_IF_NAME.io_diffCommits_info_184_v0Wen = RTL_PATH.io_diffCommits_info_184_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_184_vlWen = RTL_PATH.io_diffCommits_info_184_vlWen; \
        force U_IF_NAME.io_diffCommits_info_185_ldest = RTL_PATH.io_diffCommits_info_185_ldest; \
        force U_IF_NAME.io_diffCommits_info_185_pdest = RTL_PATH.io_diffCommits_info_185_pdest; \
        force U_IF_NAME.io_diffCommits_info_185_rfWen = RTL_PATH.io_diffCommits_info_185_rfWen; \
        force U_IF_NAME.io_diffCommits_info_185_fpWen = RTL_PATH.io_diffCommits_info_185_fpWen; \
        force U_IF_NAME.io_diffCommits_info_185_vecWen = RTL_PATH.io_diffCommits_info_185_vecWen; \
        force U_IF_NAME.io_diffCommits_info_185_v0Wen = RTL_PATH.io_diffCommits_info_185_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_185_vlWen = RTL_PATH.io_diffCommits_info_185_vlWen; \
        force U_IF_NAME.io_diffCommits_info_186_ldest = RTL_PATH.io_diffCommits_info_186_ldest; \
        force U_IF_NAME.io_diffCommits_info_186_pdest = RTL_PATH.io_diffCommits_info_186_pdest; \
        force U_IF_NAME.io_diffCommits_info_186_rfWen = RTL_PATH.io_diffCommits_info_186_rfWen; \
        force U_IF_NAME.io_diffCommits_info_186_fpWen = RTL_PATH.io_diffCommits_info_186_fpWen; \
        force U_IF_NAME.io_diffCommits_info_186_vecWen = RTL_PATH.io_diffCommits_info_186_vecWen; \
        force U_IF_NAME.io_diffCommits_info_186_v0Wen = RTL_PATH.io_diffCommits_info_186_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_186_vlWen = RTL_PATH.io_diffCommits_info_186_vlWen; \
        force U_IF_NAME.io_diffCommits_info_187_ldest = RTL_PATH.io_diffCommits_info_187_ldest; \
        force U_IF_NAME.io_diffCommits_info_187_pdest = RTL_PATH.io_diffCommits_info_187_pdest; \
        force U_IF_NAME.io_diffCommits_info_187_rfWen = RTL_PATH.io_diffCommits_info_187_rfWen; \
        force U_IF_NAME.io_diffCommits_info_187_fpWen = RTL_PATH.io_diffCommits_info_187_fpWen; \
        force U_IF_NAME.io_diffCommits_info_187_vecWen = RTL_PATH.io_diffCommits_info_187_vecWen; \
        force U_IF_NAME.io_diffCommits_info_187_v0Wen = RTL_PATH.io_diffCommits_info_187_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_187_vlWen = RTL_PATH.io_diffCommits_info_187_vlWen; \
        force U_IF_NAME.io_diffCommits_info_188_ldest = RTL_PATH.io_diffCommits_info_188_ldest; \
        force U_IF_NAME.io_diffCommits_info_188_pdest = RTL_PATH.io_diffCommits_info_188_pdest; \
        force U_IF_NAME.io_diffCommits_info_188_rfWen = RTL_PATH.io_diffCommits_info_188_rfWen; \
        force U_IF_NAME.io_diffCommits_info_188_fpWen = RTL_PATH.io_diffCommits_info_188_fpWen; \
        force U_IF_NAME.io_diffCommits_info_188_vecWen = RTL_PATH.io_diffCommits_info_188_vecWen; \
        force U_IF_NAME.io_diffCommits_info_188_v0Wen = RTL_PATH.io_diffCommits_info_188_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_188_vlWen = RTL_PATH.io_diffCommits_info_188_vlWen; \
        force U_IF_NAME.io_diffCommits_info_189_ldest = RTL_PATH.io_diffCommits_info_189_ldest; \
        force U_IF_NAME.io_diffCommits_info_189_pdest = RTL_PATH.io_diffCommits_info_189_pdest; \
        force U_IF_NAME.io_diffCommits_info_189_rfWen = RTL_PATH.io_diffCommits_info_189_rfWen; \
        force U_IF_NAME.io_diffCommits_info_189_fpWen = RTL_PATH.io_diffCommits_info_189_fpWen; \
        force U_IF_NAME.io_diffCommits_info_189_vecWen = RTL_PATH.io_diffCommits_info_189_vecWen; \
        force U_IF_NAME.io_diffCommits_info_189_v0Wen = RTL_PATH.io_diffCommits_info_189_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_189_vlWen = RTL_PATH.io_diffCommits_info_189_vlWen; \
        force U_IF_NAME.io_diffCommits_info_190_ldest = RTL_PATH.io_diffCommits_info_190_ldest; \
        force U_IF_NAME.io_diffCommits_info_190_pdest = RTL_PATH.io_diffCommits_info_190_pdest; \
        force U_IF_NAME.io_diffCommits_info_190_rfWen = RTL_PATH.io_diffCommits_info_190_rfWen; \
        force U_IF_NAME.io_diffCommits_info_190_fpWen = RTL_PATH.io_diffCommits_info_190_fpWen; \
        force U_IF_NAME.io_diffCommits_info_190_vecWen = RTL_PATH.io_diffCommits_info_190_vecWen; \
        force U_IF_NAME.io_diffCommits_info_190_v0Wen = RTL_PATH.io_diffCommits_info_190_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_190_vlWen = RTL_PATH.io_diffCommits_info_190_vlWen; \
        force U_IF_NAME.io_diffCommits_info_191_ldest = RTL_PATH.io_diffCommits_info_191_ldest; \
        force U_IF_NAME.io_diffCommits_info_191_pdest = RTL_PATH.io_diffCommits_info_191_pdest; \
        force U_IF_NAME.io_diffCommits_info_191_rfWen = RTL_PATH.io_diffCommits_info_191_rfWen; \
        force U_IF_NAME.io_diffCommits_info_191_fpWen = RTL_PATH.io_diffCommits_info_191_fpWen; \
        force U_IF_NAME.io_diffCommits_info_191_vecWen = RTL_PATH.io_diffCommits_info_191_vecWen; \
        force U_IF_NAME.io_diffCommits_info_191_v0Wen = RTL_PATH.io_diffCommits_info_191_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_191_vlWen = RTL_PATH.io_diffCommits_info_191_vlWen; \
        force U_IF_NAME.io_diffCommits_info_192_ldest = RTL_PATH.io_diffCommits_info_192_ldest; \
        force U_IF_NAME.io_diffCommits_info_192_pdest = RTL_PATH.io_diffCommits_info_192_pdest; \
        force U_IF_NAME.io_diffCommits_info_192_rfWen = RTL_PATH.io_diffCommits_info_192_rfWen; \
        force U_IF_NAME.io_diffCommits_info_192_fpWen = RTL_PATH.io_diffCommits_info_192_fpWen; \
        force U_IF_NAME.io_diffCommits_info_192_vecWen = RTL_PATH.io_diffCommits_info_192_vecWen; \
        force U_IF_NAME.io_diffCommits_info_192_v0Wen = RTL_PATH.io_diffCommits_info_192_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_192_vlWen = RTL_PATH.io_diffCommits_info_192_vlWen; \
        force U_IF_NAME.io_diffCommits_info_193_ldest = RTL_PATH.io_diffCommits_info_193_ldest; \
        force U_IF_NAME.io_diffCommits_info_193_pdest = RTL_PATH.io_diffCommits_info_193_pdest; \
        force U_IF_NAME.io_diffCommits_info_193_rfWen = RTL_PATH.io_diffCommits_info_193_rfWen; \
        force U_IF_NAME.io_diffCommits_info_193_fpWen = RTL_PATH.io_diffCommits_info_193_fpWen; \
        force U_IF_NAME.io_diffCommits_info_193_vecWen = RTL_PATH.io_diffCommits_info_193_vecWen; \
        force U_IF_NAME.io_diffCommits_info_193_v0Wen = RTL_PATH.io_diffCommits_info_193_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_193_vlWen = RTL_PATH.io_diffCommits_info_193_vlWen; \
        force U_IF_NAME.io_diffCommits_info_194_ldest = RTL_PATH.io_diffCommits_info_194_ldest; \
        force U_IF_NAME.io_diffCommits_info_194_pdest = RTL_PATH.io_diffCommits_info_194_pdest; \
        force U_IF_NAME.io_diffCommits_info_194_rfWen = RTL_PATH.io_diffCommits_info_194_rfWen; \
        force U_IF_NAME.io_diffCommits_info_194_fpWen = RTL_PATH.io_diffCommits_info_194_fpWen; \
        force U_IF_NAME.io_diffCommits_info_194_vecWen = RTL_PATH.io_diffCommits_info_194_vecWen; \
        force U_IF_NAME.io_diffCommits_info_194_v0Wen = RTL_PATH.io_diffCommits_info_194_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_194_vlWen = RTL_PATH.io_diffCommits_info_194_vlWen; \
        force U_IF_NAME.io_diffCommits_info_195_ldest = RTL_PATH.io_diffCommits_info_195_ldest; \
        force U_IF_NAME.io_diffCommits_info_195_pdest = RTL_PATH.io_diffCommits_info_195_pdest; \
        force U_IF_NAME.io_diffCommits_info_195_rfWen = RTL_PATH.io_diffCommits_info_195_rfWen; \
        force U_IF_NAME.io_diffCommits_info_195_fpWen = RTL_PATH.io_diffCommits_info_195_fpWen; \
        force U_IF_NAME.io_diffCommits_info_195_vecWen = RTL_PATH.io_diffCommits_info_195_vecWen; \
        force U_IF_NAME.io_diffCommits_info_195_v0Wen = RTL_PATH.io_diffCommits_info_195_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_195_vlWen = RTL_PATH.io_diffCommits_info_195_vlWen; \
        force U_IF_NAME.io_diffCommits_info_196_ldest = RTL_PATH.io_diffCommits_info_196_ldest; \
        force U_IF_NAME.io_diffCommits_info_196_pdest = RTL_PATH.io_diffCommits_info_196_pdest; \
        force U_IF_NAME.io_diffCommits_info_196_rfWen = RTL_PATH.io_diffCommits_info_196_rfWen; \
        force U_IF_NAME.io_diffCommits_info_196_fpWen = RTL_PATH.io_diffCommits_info_196_fpWen; \
        force U_IF_NAME.io_diffCommits_info_196_vecWen = RTL_PATH.io_diffCommits_info_196_vecWen; \
        force U_IF_NAME.io_diffCommits_info_196_v0Wen = RTL_PATH.io_diffCommits_info_196_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_196_vlWen = RTL_PATH.io_diffCommits_info_196_vlWen; \
        force U_IF_NAME.io_diffCommits_info_197_ldest = RTL_PATH.io_diffCommits_info_197_ldest; \
        force U_IF_NAME.io_diffCommits_info_197_pdest = RTL_PATH.io_diffCommits_info_197_pdest; \
        force U_IF_NAME.io_diffCommits_info_197_rfWen = RTL_PATH.io_diffCommits_info_197_rfWen; \
        force U_IF_NAME.io_diffCommits_info_197_fpWen = RTL_PATH.io_diffCommits_info_197_fpWen; \
        force U_IF_NAME.io_diffCommits_info_197_vecWen = RTL_PATH.io_diffCommits_info_197_vecWen; \
        force U_IF_NAME.io_diffCommits_info_197_v0Wen = RTL_PATH.io_diffCommits_info_197_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_197_vlWen = RTL_PATH.io_diffCommits_info_197_vlWen; \
        force U_IF_NAME.io_diffCommits_info_198_ldest = RTL_PATH.io_diffCommits_info_198_ldest; \
        force U_IF_NAME.io_diffCommits_info_198_pdest = RTL_PATH.io_diffCommits_info_198_pdest; \
        force U_IF_NAME.io_diffCommits_info_198_rfWen = RTL_PATH.io_diffCommits_info_198_rfWen; \
        force U_IF_NAME.io_diffCommits_info_198_fpWen = RTL_PATH.io_diffCommits_info_198_fpWen; \
        force U_IF_NAME.io_diffCommits_info_198_vecWen = RTL_PATH.io_diffCommits_info_198_vecWen; \
        force U_IF_NAME.io_diffCommits_info_198_v0Wen = RTL_PATH.io_diffCommits_info_198_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_198_vlWen = RTL_PATH.io_diffCommits_info_198_vlWen; \
        force U_IF_NAME.io_diffCommits_info_199_ldest = RTL_PATH.io_diffCommits_info_199_ldest; \
        force U_IF_NAME.io_diffCommits_info_199_pdest = RTL_PATH.io_diffCommits_info_199_pdest; \
        force U_IF_NAME.io_diffCommits_info_199_rfWen = RTL_PATH.io_diffCommits_info_199_rfWen; \
        force U_IF_NAME.io_diffCommits_info_199_fpWen = RTL_PATH.io_diffCommits_info_199_fpWen; \
        force U_IF_NAME.io_diffCommits_info_199_vecWen = RTL_PATH.io_diffCommits_info_199_vecWen; \
        force U_IF_NAME.io_diffCommits_info_199_v0Wen = RTL_PATH.io_diffCommits_info_199_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_199_vlWen = RTL_PATH.io_diffCommits_info_199_vlWen; \
        force U_IF_NAME.io_diffCommits_info_200_ldest = RTL_PATH.io_diffCommits_info_200_ldest; \
        force U_IF_NAME.io_diffCommits_info_200_pdest = RTL_PATH.io_diffCommits_info_200_pdest; \
        force U_IF_NAME.io_diffCommits_info_200_rfWen = RTL_PATH.io_diffCommits_info_200_rfWen; \
        force U_IF_NAME.io_diffCommits_info_200_fpWen = RTL_PATH.io_diffCommits_info_200_fpWen; \
        force U_IF_NAME.io_diffCommits_info_200_vecWen = RTL_PATH.io_diffCommits_info_200_vecWen; \
        force U_IF_NAME.io_diffCommits_info_200_v0Wen = RTL_PATH.io_diffCommits_info_200_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_200_vlWen = RTL_PATH.io_diffCommits_info_200_vlWen; \
        force U_IF_NAME.io_diffCommits_info_201_ldest = RTL_PATH.io_diffCommits_info_201_ldest; \
        force U_IF_NAME.io_diffCommits_info_201_pdest = RTL_PATH.io_diffCommits_info_201_pdest; \
        force U_IF_NAME.io_diffCommits_info_201_rfWen = RTL_PATH.io_diffCommits_info_201_rfWen; \
        force U_IF_NAME.io_diffCommits_info_201_fpWen = RTL_PATH.io_diffCommits_info_201_fpWen; \
        force U_IF_NAME.io_diffCommits_info_201_vecWen = RTL_PATH.io_diffCommits_info_201_vecWen; \
        force U_IF_NAME.io_diffCommits_info_201_v0Wen = RTL_PATH.io_diffCommits_info_201_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_201_vlWen = RTL_PATH.io_diffCommits_info_201_vlWen; \
        force U_IF_NAME.io_diffCommits_info_202_ldest = RTL_PATH.io_diffCommits_info_202_ldest; \
        force U_IF_NAME.io_diffCommits_info_202_pdest = RTL_PATH.io_diffCommits_info_202_pdest; \
        force U_IF_NAME.io_diffCommits_info_202_rfWen = RTL_PATH.io_diffCommits_info_202_rfWen; \
        force U_IF_NAME.io_diffCommits_info_202_fpWen = RTL_PATH.io_diffCommits_info_202_fpWen; \
        force U_IF_NAME.io_diffCommits_info_202_vecWen = RTL_PATH.io_diffCommits_info_202_vecWen; \
        force U_IF_NAME.io_diffCommits_info_202_v0Wen = RTL_PATH.io_diffCommits_info_202_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_202_vlWen = RTL_PATH.io_diffCommits_info_202_vlWen; \
        force U_IF_NAME.io_diffCommits_info_203_ldest = RTL_PATH.io_diffCommits_info_203_ldest; \
        force U_IF_NAME.io_diffCommits_info_203_pdest = RTL_PATH.io_diffCommits_info_203_pdest; \
        force U_IF_NAME.io_diffCommits_info_203_rfWen = RTL_PATH.io_diffCommits_info_203_rfWen; \
        force U_IF_NAME.io_diffCommits_info_203_fpWen = RTL_PATH.io_diffCommits_info_203_fpWen; \
        force U_IF_NAME.io_diffCommits_info_203_vecWen = RTL_PATH.io_diffCommits_info_203_vecWen; \
        force U_IF_NAME.io_diffCommits_info_203_v0Wen = RTL_PATH.io_diffCommits_info_203_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_203_vlWen = RTL_PATH.io_diffCommits_info_203_vlWen; \
        force U_IF_NAME.io_diffCommits_info_204_ldest = RTL_PATH.io_diffCommits_info_204_ldest; \
        force U_IF_NAME.io_diffCommits_info_204_pdest = RTL_PATH.io_diffCommits_info_204_pdest; \
        force U_IF_NAME.io_diffCommits_info_204_rfWen = RTL_PATH.io_diffCommits_info_204_rfWen; \
        force U_IF_NAME.io_diffCommits_info_204_fpWen = RTL_PATH.io_diffCommits_info_204_fpWen; \
        force U_IF_NAME.io_diffCommits_info_204_vecWen = RTL_PATH.io_diffCommits_info_204_vecWen; \
        force U_IF_NAME.io_diffCommits_info_204_v0Wen = RTL_PATH.io_diffCommits_info_204_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_204_vlWen = RTL_PATH.io_diffCommits_info_204_vlWen; \
        force U_IF_NAME.io_diffCommits_info_205_ldest = RTL_PATH.io_diffCommits_info_205_ldest; \
        force U_IF_NAME.io_diffCommits_info_205_pdest = RTL_PATH.io_diffCommits_info_205_pdest; \
        force U_IF_NAME.io_diffCommits_info_205_rfWen = RTL_PATH.io_diffCommits_info_205_rfWen; \
        force U_IF_NAME.io_diffCommits_info_205_fpWen = RTL_PATH.io_diffCommits_info_205_fpWen; \
        force U_IF_NAME.io_diffCommits_info_205_vecWen = RTL_PATH.io_diffCommits_info_205_vecWen; \
        force U_IF_NAME.io_diffCommits_info_205_v0Wen = RTL_PATH.io_diffCommits_info_205_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_205_vlWen = RTL_PATH.io_diffCommits_info_205_vlWen; \
        force U_IF_NAME.io_diffCommits_info_206_ldest = RTL_PATH.io_diffCommits_info_206_ldest; \
        force U_IF_NAME.io_diffCommits_info_206_pdest = RTL_PATH.io_diffCommits_info_206_pdest; \
        force U_IF_NAME.io_diffCommits_info_206_rfWen = RTL_PATH.io_diffCommits_info_206_rfWen; \
        force U_IF_NAME.io_diffCommits_info_206_fpWen = RTL_PATH.io_diffCommits_info_206_fpWen; \
        force U_IF_NAME.io_diffCommits_info_206_vecWen = RTL_PATH.io_diffCommits_info_206_vecWen; \
        force U_IF_NAME.io_diffCommits_info_206_v0Wen = RTL_PATH.io_diffCommits_info_206_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_206_vlWen = RTL_PATH.io_diffCommits_info_206_vlWen; \
        force U_IF_NAME.io_diffCommits_info_207_ldest = RTL_PATH.io_diffCommits_info_207_ldest; \
        force U_IF_NAME.io_diffCommits_info_207_pdest = RTL_PATH.io_diffCommits_info_207_pdest; \
        force U_IF_NAME.io_diffCommits_info_207_rfWen = RTL_PATH.io_diffCommits_info_207_rfWen; \
        force U_IF_NAME.io_diffCommits_info_207_fpWen = RTL_PATH.io_diffCommits_info_207_fpWen; \
        force U_IF_NAME.io_diffCommits_info_207_vecWen = RTL_PATH.io_diffCommits_info_207_vecWen; \
        force U_IF_NAME.io_diffCommits_info_207_v0Wen = RTL_PATH.io_diffCommits_info_207_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_207_vlWen = RTL_PATH.io_diffCommits_info_207_vlWen; \
        force U_IF_NAME.io_diffCommits_info_208_ldest = RTL_PATH.io_diffCommits_info_208_ldest; \
        force U_IF_NAME.io_diffCommits_info_208_pdest = RTL_PATH.io_diffCommits_info_208_pdest; \
        force U_IF_NAME.io_diffCommits_info_208_rfWen = RTL_PATH.io_diffCommits_info_208_rfWen; \
        force U_IF_NAME.io_diffCommits_info_208_fpWen = RTL_PATH.io_diffCommits_info_208_fpWen; \
        force U_IF_NAME.io_diffCommits_info_208_vecWen = RTL_PATH.io_diffCommits_info_208_vecWen; \
        force U_IF_NAME.io_diffCommits_info_208_v0Wen = RTL_PATH.io_diffCommits_info_208_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_208_vlWen = RTL_PATH.io_diffCommits_info_208_vlWen; \
        force U_IF_NAME.io_diffCommits_info_209_ldest = RTL_PATH.io_diffCommits_info_209_ldest; \
        force U_IF_NAME.io_diffCommits_info_209_pdest = RTL_PATH.io_diffCommits_info_209_pdest; \
        force U_IF_NAME.io_diffCommits_info_209_rfWen = RTL_PATH.io_diffCommits_info_209_rfWen; \
        force U_IF_NAME.io_diffCommits_info_209_fpWen = RTL_PATH.io_diffCommits_info_209_fpWen; \
        force U_IF_NAME.io_diffCommits_info_209_vecWen = RTL_PATH.io_diffCommits_info_209_vecWen; \
        force U_IF_NAME.io_diffCommits_info_209_v0Wen = RTL_PATH.io_diffCommits_info_209_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_209_vlWen = RTL_PATH.io_diffCommits_info_209_vlWen; \
        force U_IF_NAME.io_diffCommits_info_210_ldest = RTL_PATH.io_diffCommits_info_210_ldest; \
        force U_IF_NAME.io_diffCommits_info_210_pdest = RTL_PATH.io_diffCommits_info_210_pdest; \
        force U_IF_NAME.io_diffCommits_info_210_rfWen = RTL_PATH.io_diffCommits_info_210_rfWen; \
        force U_IF_NAME.io_diffCommits_info_210_fpWen = RTL_PATH.io_diffCommits_info_210_fpWen; \
        force U_IF_NAME.io_diffCommits_info_210_vecWen = RTL_PATH.io_diffCommits_info_210_vecWen; \
        force U_IF_NAME.io_diffCommits_info_210_v0Wen = RTL_PATH.io_diffCommits_info_210_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_210_vlWen = RTL_PATH.io_diffCommits_info_210_vlWen; \
        force U_IF_NAME.io_diffCommits_info_211_ldest = RTL_PATH.io_diffCommits_info_211_ldest; \
        force U_IF_NAME.io_diffCommits_info_211_pdest = RTL_PATH.io_diffCommits_info_211_pdest; \
        force U_IF_NAME.io_diffCommits_info_211_rfWen = RTL_PATH.io_diffCommits_info_211_rfWen; \
        force U_IF_NAME.io_diffCommits_info_211_fpWen = RTL_PATH.io_diffCommits_info_211_fpWen; \
        force U_IF_NAME.io_diffCommits_info_211_vecWen = RTL_PATH.io_diffCommits_info_211_vecWen; \
        force U_IF_NAME.io_diffCommits_info_211_v0Wen = RTL_PATH.io_diffCommits_info_211_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_211_vlWen = RTL_PATH.io_diffCommits_info_211_vlWen; \
        force U_IF_NAME.io_diffCommits_info_212_ldest = RTL_PATH.io_diffCommits_info_212_ldest; \
        force U_IF_NAME.io_diffCommits_info_212_pdest = RTL_PATH.io_diffCommits_info_212_pdest; \
        force U_IF_NAME.io_diffCommits_info_212_rfWen = RTL_PATH.io_diffCommits_info_212_rfWen; \
        force U_IF_NAME.io_diffCommits_info_212_fpWen = RTL_PATH.io_diffCommits_info_212_fpWen; \
        force U_IF_NAME.io_diffCommits_info_212_vecWen = RTL_PATH.io_diffCommits_info_212_vecWen; \
        force U_IF_NAME.io_diffCommits_info_212_v0Wen = RTL_PATH.io_diffCommits_info_212_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_212_vlWen = RTL_PATH.io_diffCommits_info_212_vlWen; \
        force U_IF_NAME.io_diffCommits_info_213_ldest = RTL_PATH.io_diffCommits_info_213_ldest; \
        force U_IF_NAME.io_diffCommits_info_213_pdest = RTL_PATH.io_diffCommits_info_213_pdest; \
        force U_IF_NAME.io_diffCommits_info_213_rfWen = RTL_PATH.io_diffCommits_info_213_rfWen; \
        force U_IF_NAME.io_diffCommits_info_213_fpWen = RTL_PATH.io_diffCommits_info_213_fpWen; \
        force U_IF_NAME.io_diffCommits_info_213_vecWen = RTL_PATH.io_diffCommits_info_213_vecWen; \
        force U_IF_NAME.io_diffCommits_info_213_v0Wen = RTL_PATH.io_diffCommits_info_213_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_213_vlWen = RTL_PATH.io_diffCommits_info_213_vlWen; \
        force U_IF_NAME.io_diffCommits_info_214_ldest = RTL_PATH.io_diffCommits_info_214_ldest; \
        force U_IF_NAME.io_diffCommits_info_214_pdest = RTL_PATH.io_diffCommits_info_214_pdest; \
        force U_IF_NAME.io_diffCommits_info_214_rfWen = RTL_PATH.io_diffCommits_info_214_rfWen; \
        force U_IF_NAME.io_diffCommits_info_214_fpWen = RTL_PATH.io_diffCommits_info_214_fpWen; \
        force U_IF_NAME.io_diffCommits_info_214_vecWen = RTL_PATH.io_diffCommits_info_214_vecWen; \
        force U_IF_NAME.io_diffCommits_info_214_v0Wen = RTL_PATH.io_diffCommits_info_214_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_214_vlWen = RTL_PATH.io_diffCommits_info_214_vlWen; \
        force U_IF_NAME.io_diffCommits_info_215_ldest = RTL_PATH.io_diffCommits_info_215_ldest; \
        force U_IF_NAME.io_diffCommits_info_215_pdest = RTL_PATH.io_diffCommits_info_215_pdest; \
        force U_IF_NAME.io_diffCommits_info_215_rfWen = RTL_PATH.io_diffCommits_info_215_rfWen; \
        force U_IF_NAME.io_diffCommits_info_215_fpWen = RTL_PATH.io_diffCommits_info_215_fpWen; \
        force U_IF_NAME.io_diffCommits_info_215_vecWen = RTL_PATH.io_diffCommits_info_215_vecWen; \
        force U_IF_NAME.io_diffCommits_info_215_v0Wen = RTL_PATH.io_diffCommits_info_215_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_215_vlWen = RTL_PATH.io_diffCommits_info_215_vlWen; \
        force U_IF_NAME.io_diffCommits_info_216_ldest = RTL_PATH.io_diffCommits_info_216_ldest; \
        force U_IF_NAME.io_diffCommits_info_216_pdest = RTL_PATH.io_diffCommits_info_216_pdest; \
        force U_IF_NAME.io_diffCommits_info_216_rfWen = RTL_PATH.io_diffCommits_info_216_rfWen; \
        force U_IF_NAME.io_diffCommits_info_216_fpWen = RTL_PATH.io_diffCommits_info_216_fpWen; \
        force U_IF_NAME.io_diffCommits_info_216_vecWen = RTL_PATH.io_diffCommits_info_216_vecWen; \
        force U_IF_NAME.io_diffCommits_info_216_v0Wen = RTL_PATH.io_diffCommits_info_216_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_216_vlWen = RTL_PATH.io_diffCommits_info_216_vlWen; \
        force U_IF_NAME.io_diffCommits_info_217_ldest = RTL_PATH.io_diffCommits_info_217_ldest; \
        force U_IF_NAME.io_diffCommits_info_217_pdest = RTL_PATH.io_diffCommits_info_217_pdest; \
        force U_IF_NAME.io_diffCommits_info_217_rfWen = RTL_PATH.io_diffCommits_info_217_rfWen; \
        force U_IF_NAME.io_diffCommits_info_217_fpWen = RTL_PATH.io_diffCommits_info_217_fpWen; \
        force U_IF_NAME.io_diffCommits_info_217_vecWen = RTL_PATH.io_diffCommits_info_217_vecWen; \
        force U_IF_NAME.io_diffCommits_info_217_v0Wen = RTL_PATH.io_diffCommits_info_217_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_217_vlWen = RTL_PATH.io_diffCommits_info_217_vlWen; \
        force U_IF_NAME.io_diffCommits_info_218_ldest = RTL_PATH.io_diffCommits_info_218_ldest; \
        force U_IF_NAME.io_diffCommits_info_218_pdest = RTL_PATH.io_diffCommits_info_218_pdest; \
        force U_IF_NAME.io_diffCommits_info_218_rfWen = RTL_PATH.io_diffCommits_info_218_rfWen; \
        force U_IF_NAME.io_diffCommits_info_218_fpWen = RTL_PATH.io_diffCommits_info_218_fpWen; \
        force U_IF_NAME.io_diffCommits_info_218_vecWen = RTL_PATH.io_diffCommits_info_218_vecWen; \
        force U_IF_NAME.io_diffCommits_info_218_v0Wen = RTL_PATH.io_diffCommits_info_218_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_218_vlWen = RTL_PATH.io_diffCommits_info_218_vlWen; \
        force U_IF_NAME.io_diffCommits_info_219_ldest = RTL_PATH.io_diffCommits_info_219_ldest; \
        force U_IF_NAME.io_diffCommits_info_219_pdest = RTL_PATH.io_diffCommits_info_219_pdest; \
        force U_IF_NAME.io_diffCommits_info_219_rfWen = RTL_PATH.io_diffCommits_info_219_rfWen; \
        force U_IF_NAME.io_diffCommits_info_219_fpWen = RTL_PATH.io_diffCommits_info_219_fpWen; \
        force U_IF_NAME.io_diffCommits_info_219_vecWen = RTL_PATH.io_diffCommits_info_219_vecWen; \
        force U_IF_NAME.io_diffCommits_info_219_v0Wen = RTL_PATH.io_diffCommits_info_219_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_219_vlWen = RTL_PATH.io_diffCommits_info_219_vlWen; \
        force U_IF_NAME.io_diffCommits_info_220_ldest = RTL_PATH.io_diffCommits_info_220_ldest; \
        force U_IF_NAME.io_diffCommits_info_220_pdest = RTL_PATH.io_diffCommits_info_220_pdest; \
        force U_IF_NAME.io_diffCommits_info_220_rfWen = RTL_PATH.io_diffCommits_info_220_rfWen; \
        force U_IF_NAME.io_diffCommits_info_220_fpWen = RTL_PATH.io_diffCommits_info_220_fpWen; \
        force U_IF_NAME.io_diffCommits_info_220_vecWen = RTL_PATH.io_diffCommits_info_220_vecWen; \
        force U_IF_NAME.io_diffCommits_info_220_v0Wen = RTL_PATH.io_diffCommits_info_220_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_220_vlWen = RTL_PATH.io_diffCommits_info_220_vlWen; \
        force U_IF_NAME.io_diffCommits_info_221_ldest = RTL_PATH.io_diffCommits_info_221_ldest; \
        force U_IF_NAME.io_diffCommits_info_221_pdest = RTL_PATH.io_diffCommits_info_221_pdest; \
        force U_IF_NAME.io_diffCommits_info_221_rfWen = RTL_PATH.io_diffCommits_info_221_rfWen; \
        force U_IF_NAME.io_diffCommits_info_221_fpWen = RTL_PATH.io_diffCommits_info_221_fpWen; \
        force U_IF_NAME.io_diffCommits_info_221_vecWen = RTL_PATH.io_diffCommits_info_221_vecWen; \
        force U_IF_NAME.io_diffCommits_info_221_v0Wen = RTL_PATH.io_diffCommits_info_221_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_221_vlWen = RTL_PATH.io_diffCommits_info_221_vlWen; \
        force U_IF_NAME.io_diffCommits_info_222_ldest = RTL_PATH.io_diffCommits_info_222_ldest; \
        force U_IF_NAME.io_diffCommits_info_222_pdest = RTL_PATH.io_diffCommits_info_222_pdest; \
        force U_IF_NAME.io_diffCommits_info_222_rfWen = RTL_PATH.io_diffCommits_info_222_rfWen; \
        force U_IF_NAME.io_diffCommits_info_222_fpWen = RTL_PATH.io_diffCommits_info_222_fpWen; \
        force U_IF_NAME.io_diffCommits_info_222_vecWen = RTL_PATH.io_diffCommits_info_222_vecWen; \
        force U_IF_NAME.io_diffCommits_info_222_v0Wen = RTL_PATH.io_diffCommits_info_222_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_222_vlWen = RTL_PATH.io_diffCommits_info_222_vlWen; \
        force U_IF_NAME.io_diffCommits_info_223_ldest = RTL_PATH.io_diffCommits_info_223_ldest; \
        force U_IF_NAME.io_diffCommits_info_223_pdest = RTL_PATH.io_diffCommits_info_223_pdest; \
        force U_IF_NAME.io_diffCommits_info_223_rfWen = RTL_PATH.io_diffCommits_info_223_rfWen; \
        force U_IF_NAME.io_diffCommits_info_223_fpWen = RTL_PATH.io_diffCommits_info_223_fpWen; \
        force U_IF_NAME.io_diffCommits_info_223_vecWen = RTL_PATH.io_diffCommits_info_223_vecWen; \
        force U_IF_NAME.io_diffCommits_info_223_v0Wen = RTL_PATH.io_diffCommits_info_223_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_223_vlWen = RTL_PATH.io_diffCommits_info_223_vlWen; \
        force U_IF_NAME.io_diffCommits_info_224_ldest = RTL_PATH.io_diffCommits_info_224_ldest; \
        force U_IF_NAME.io_diffCommits_info_224_pdest = RTL_PATH.io_diffCommits_info_224_pdest; \
        force U_IF_NAME.io_diffCommits_info_224_rfWen = RTL_PATH.io_diffCommits_info_224_rfWen; \
        force U_IF_NAME.io_diffCommits_info_224_fpWen = RTL_PATH.io_diffCommits_info_224_fpWen; \
        force U_IF_NAME.io_diffCommits_info_224_vecWen = RTL_PATH.io_diffCommits_info_224_vecWen; \
        force U_IF_NAME.io_diffCommits_info_224_v0Wen = RTL_PATH.io_diffCommits_info_224_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_224_vlWen = RTL_PATH.io_diffCommits_info_224_vlWen; \
        force U_IF_NAME.io_diffCommits_info_225_ldest = RTL_PATH.io_diffCommits_info_225_ldest; \
        force U_IF_NAME.io_diffCommits_info_225_pdest = RTL_PATH.io_diffCommits_info_225_pdest; \
        force U_IF_NAME.io_diffCommits_info_225_rfWen = RTL_PATH.io_diffCommits_info_225_rfWen; \
        force U_IF_NAME.io_diffCommits_info_225_fpWen = RTL_PATH.io_diffCommits_info_225_fpWen; \
        force U_IF_NAME.io_diffCommits_info_225_vecWen = RTL_PATH.io_diffCommits_info_225_vecWen; \
        force U_IF_NAME.io_diffCommits_info_225_v0Wen = RTL_PATH.io_diffCommits_info_225_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_225_vlWen = RTL_PATH.io_diffCommits_info_225_vlWen; \
        force U_IF_NAME.io_diffCommits_info_226_ldest = RTL_PATH.io_diffCommits_info_226_ldest; \
        force U_IF_NAME.io_diffCommits_info_226_pdest = RTL_PATH.io_diffCommits_info_226_pdest; \
        force U_IF_NAME.io_diffCommits_info_226_rfWen = RTL_PATH.io_diffCommits_info_226_rfWen; \
        force U_IF_NAME.io_diffCommits_info_226_fpWen = RTL_PATH.io_diffCommits_info_226_fpWen; \
        force U_IF_NAME.io_diffCommits_info_226_vecWen = RTL_PATH.io_diffCommits_info_226_vecWen; \
        force U_IF_NAME.io_diffCommits_info_226_v0Wen = RTL_PATH.io_diffCommits_info_226_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_226_vlWen = RTL_PATH.io_diffCommits_info_226_vlWen; \
        force U_IF_NAME.io_diffCommits_info_227_ldest = RTL_PATH.io_diffCommits_info_227_ldest; \
        force U_IF_NAME.io_diffCommits_info_227_pdest = RTL_PATH.io_diffCommits_info_227_pdest; \
        force U_IF_NAME.io_diffCommits_info_227_rfWen = RTL_PATH.io_diffCommits_info_227_rfWen; \
        force U_IF_NAME.io_diffCommits_info_227_fpWen = RTL_PATH.io_diffCommits_info_227_fpWen; \
        force U_IF_NAME.io_diffCommits_info_227_vecWen = RTL_PATH.io_diffCommits_info_227_vecWen; \
        force U_IF_NAME.io_diffCommits_info_227_v0Wen = RTL_PATH.io_diffCommits_info_227_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_227_vlWen = RTL_PATH.io_diffCommits_info_227_vlWen; \
        force U_IF_NAME.io_diffCommits_info_228_ldest = RTL_PATH.io_diffCommits_info_228_ldest; \
        force U_IF_NAME.io_diffCommits_info_228_pdest = RTL_PATH.io_diffCommits_info_228_pdest; \
        force U_IF_NAME.io_diffCommits_info_228_rfWen = RTL_PATH.io_diffCommits_info_228_rfWen; \
        force U_IF_NAME.io_diffCommits_info_228_fpWen = RTL_PATH.io_diffCommits_info_228_fpWen; \
        force U_IF_NAME.io_diffCommits_info_228_vecWen = RTL_PATH.io_diffCommits_info_228_vecWen; \
        force U_IF_NAME.io_diffCommits_info_228_v0Wen = RTL_PATH.io_diffCommits_info_228_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_228_vlWen = RTL_PATH.io_diffCommits_info_228_vlWen; \
        force U_IF_NAME.io_diffCommits_info_229_ldest = RTL_PATH.io_diffCommits_info_229_ldest; \
        force U_IF_NAME.io_diffCommits_info_229_pdest = RTL_PATH.io_diffCommits_info_229_pdest; \
        force U_IF_NAME.io_diffCommits_info_229_rfWen = RTL_PATH.io_diffCommits_info_229_rfWen; \
        force U_IF_NAME.io_diffCommits_info_229_fpWen = RTL_PATH.io_diffCommits_info_229_fpWen; \
        force U_IF_NAME.io_diffCommits_info_229_vecWen = RTL_PATH.io_diffCommits_info_229_vecWen; \
        force U_IF_NAME.io_diffCommits_info_229_v0Wen = RTL_PATH.io_diffCommits_info_229_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_229_vlWen = RTL_PATH.io_diffCommits_info_229_vlWen; \
        force U_IF_NAME.io_diffCommits_info_230_ldest = RTL_PATH.io_diffCommits_info_230_ldest; \
        force U_IF_NAME.io_diffCommits_info_230_pdest = RTL_PATH.io_diffCommits_info_230_pdest; \
        force U_IF_NAME.io_diffCommits_info_230_rfWen = RTL_PATH.io_diffCommits_info_230_rfWen; \
        force U_IF_NAME.io_diffCommits_info_230_fpWen = RTL_PATH.io_diffCommits_info_230_fpWen; \
        force U_IF_NAME.io_diffCommits_info_230_vecWen = RTL_PATH.io_diffCommits_info_230_vecWen; \
        force U_IF_NAME.io_diffCommits_info_230_v0Wen = RTL_PATH.io_diffCommits_info_230_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_230_vlWen = RTL_PATH.io_diffCommits_info_230_vlWen; \
        force U_IF_NAME.io_diffCommits_info_231_ldest = RTL_PATH.io_diffCommits_info_231_ldest; \
        force U_IF_NAME.io_diffCommits_info_231_pdest = RTL_PATH.io_diffCommits_info_231_pdest; \
        force U_IF_NAME.io_diffCommits_info_231_rfWen = RTL_PATH.io_diffCommits_info_231_rfWen; \
        force U_IF_NAME.io_diffCommits_info_231_fpWen = RTL_PATH.io_diffCommits_info_231_fpWen; \
        force U_IF_NAME.io_diffCommits_info_231_vecWen = RTL_PATH.io_diffCommits_info_231_vecWen; \
        force U_IF_NAME.io_diffCommits_info_231_v0Wen = RTL_PATH.io_diffCommits_info_231_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_231_vlWen = RTL_PATH.io_diffCommits_info_231_vlWen; \
        force U_IF_NAME.io_diffCommits_info_232_ldest = RTL_PATH.io_diffCommits_info_232_ldest; \
        force U_IF_NAME.io_diffCommits_info_232_pdest = RTL_PATH.io_diffCommits_info_232_pdest; \
        force U_IF_NAME.io_diffCommits_info_232_rfWen = RTL_PATH.io_diffCommits_info_232_rfWen; \
        force U_IF_NAME.io_diffCommits_info_232_fpWen = RTL_PATH.io_diffCommits_info_232_fpWen; \
        force U_IF_NAME.io_diffCommits_info_232_vecWen = RTL_PATH.io_diffCommits_info_232_vecWen; \
        force U_IF_NAME.io_diffCommits_info_232_v0Wen = RTL_PATH.io_diffCommits_info_232_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_232_vlWen = RTL_PATH.io_diffCommits_info_232_vlWen; \
        force U_IF_NAME.io_diffCommits_info_233_ldest = RTL_PATH.io_diffCommits_info_233_ldest; \
        force U_IF_NAME.io_diffCommits_info_233_pdest = RTL_PATH.io_diffCommits_info_233_pdest; \
        force U_IF_NAME.io_diffCommits_info_233_rfWen = RTL_PATH.io_diffCommits_info_233_rfWen; \
        force U_IF_NAME.io_diffCommits_info_233_fpWen = RTL_PATH.io_diffCommits_info_233_fpWen; \
        force U_IF_NAME.io_diffCommits_info_233_vecWen = RTL_PATH.io_diffCommits_info_233_vecWen; \
        force U_IF_NAME.io_diffCommits_info_233_v0Wen = RTL_PATH.io_diffCommits_info_233_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_233_vlWen = RTL_PATH.io_diffCommits_info_233_vlWen; \
        force U_IF_NAME.io_diffCommits_info_234_ldest = RTL_PATH.io_diffCommits_info_234_ldest; \
        force U_IF_NAME.io_diffCommits_info_234_pdest = RTL_PATH.io_diffCommits_info_234_pdest; \
        force U_IF_NAME.io_diffCommits_info_234_rfWen = RTL_PATH.io_diffCommits_info_234_rfWen; \
        force U_IF_NAME.io_diffCommits_info_234_fpWen = RTL_PATH.io_diffCommits_info_234_fpWen; \
        force U_IF_NAME.io_diffCommits_info_234_vecWen = RTL_PATH.io_diffCommits_info_234_vecWen; \
        force U_IF_NAME.io_diffCommits_info_234_v0Wen = RTL_PATH.io_diffCommits_info_234_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_234_vlWen = RTL_PATH.io_diffCommits_info_234_vlWen; \
        force U_IF_NAME.io_diffCommits_info_235_ldest = RTL_PATH.io_diffCommits_info_235_ldest; \
        force U_IF_NAME.io_diffCommits_info_235_pdest = RTL_PATH.io_diffCommits_info_235_pdest; \
        force U_IF_NAME.io_diffCommits_info_235_rfWen = RTL_PATH.io_diffCommits_info_235_rfWen; \
        force U_IF_NAME.io_diffCommits_info_235_fpWen = RTL_PATH.io_diffCommits_info_235_fpWen; \
        force U_IF_NAME.io_diffCommits_info_235_vecWen = RTL_PATH.io_diffCommits_info_235_vecWen; \
        force U_IF_NAME.io_diffCommits_info_235_v0Wen = RTL_PATH.io_diffCommits_info_235_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_235_vlWen = RTL_PATH.io_diffCommits_info_235_vlWen; \
        force U_IF_NAME.io_diffCommits_info_236_ldest = RTL_PATH.io_diffCommits_info_236_ldest; \
        force U_IF_NAME.io_diffCommits_info_236_pdest = RTL_PATH.io_diffCommits_info_236_pdest; \
        force U_IF_NAME.io_diffCommits_info_236_rfWen = RTL_PATH.io_diffCommits_info_236_rfWen; \
        force U_IF_NAME.io_diffCommits_info_236_fpWen = RTL_PATH.io_diffCommits_info_236_fpWen; \
        force U_IF_NAME.io_diffCommits_info_236_vecWen = RTL_PATH.io_diffCommits_info_236_vecWen; \
        force U_IF_NAME.io_diffCommits_info_236_v0Wen = RTL_PATH.io_diffCommits_info_236_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_236_vlWen = RTL_PATH.io_diffCommits_info_236_vlWen; \
        force U_IF_NAME.io_diffCommits_info_237_ldest = RTL_PATH.io_diffCommits_info_237_ldest; \
        force U_IF_NAME.io_diffCommits_info_237_pdest = RTL_PATH.io_diffCommits_info_237_pdest; \
        force U_IF_NAME.io_diffCommits_info_237_rfWen = RTL_PATH.io_diffCommits_info_237_rfWen; \
        force U_IF_NAME.io_diffCommits_info_237_fpWen = RTL_PATH.io_diffCommits_info_237_fpWen; \
        force U_IF_NAME.io_diffCommits_info_237_vecWen = RTL_PATH.io_diffCommits_info_237_vecWen; \
        force U_IF_NAME.io_diffCommits_info_237_v0Wen = RTL_PATH.io_diffCommits_info_237_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_237_vlWen = RTL_PATH.io_diffCommits_info_237_vlWen; \
        force U_IF_NAME.io_diffCommits_info_238_ldest = RTL_PATH.io_diffCommits_info_238_ldest; \
        force U_IF_NAME.io_diffCommits_info_238_pdest = RTL_PATH.io_diffCommits_info_238_pdest; \
        force U_IF_NAME.io_diffCommits_info_238_rfWen = RTL_PATH.io_diffCommits_info_238_rfWen; \
        force U_IF_NAME.io_diffCommits_info_238_fpWen = RTL_PATH.io_diffCommits_info_238_fpWen; \
        force U_IF_NAME.io_diffCommits_info_238_vecWen = RTL_PATH.io_diffCommits_info_238_vecWen; \
        force U_IF_NAME.io_diffCommits_info_238_v0Wen = RTL_PATH.io_diffCommits_info_238_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_238_vlWen = RTL_PATH.io_diffCommits_info_238_vlWen; \
        force U_IF_NAME.io_diffCommits_info_239_ldest = RTL_PATH.io_diffCommits_info_239_ldest; \
        force U_IF_NAME.io_diffCommits_info_239_pdest = RTL_PATH.io_diffCommits_info_239_pdest; \
        force U_IF_NAME.io_diffCommits_info_239_rfWen = RTL_PATH.io_diffCommits_info_239_rfWen; \
        force U_IF_NAME.io_diffCommits_info_239_fpWen = RTL_PATH.io_diffCommits_info_239_fpWen; \
        force U_IF_NAME.io_diffCommits_info_239_vecWen = RTL_PATH.io_diffCommits_info_239_vecWen; \
        force U_IF_NAME.io_diffCommits_info_239_v0Wen = RTL_PATH.io_diffCommits_info_239_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_239_vlWen = RTL_PATH.io_diffCommits_info_239_vlWen; \
        force U_IF_NAME.io_diffCommits_info_240_ldest = RTL_PATH.io_diffCommits_info_240_ldest; \
        force U_IF_NAME.io_diffCommits_info_240_pdest = RTL_PATH.io_diffCommits_info_240_pdest; \
        force U_IF_NAME.io_diffCommits_info_240_rfWen = RTL_PATH.io_diffCommits_info_240_rfWen; \
        force U_IF_NAME.io_diffCommits_info_240_fpWen = RTL_PATH.io_diffCommits_info_240_fpWen; \
        force U_IF_NAME.io_diffCommits_info_240_vecWen = RTL_PATH.io_diffCommits_info_240_vecWen; \
        force U_IF_NAME.io_diffCommits_info_240_v0Wen = RTL_PATH.io_diffCommits_info_240_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_240_vlWen = RTL_PATH.io_diffCommits_info_240_vlWen; \
        force U_IF_NAME.io_diffCommits_info_241_ldest = RTL_PATH.io_diffCommits_info_241_ldest; \
        force U_IF_NAME.io_diffCommits_info_241_pdest = RTL_PATH.io_diffCommits_info_241_pdest; \
        force U_IF_NAME.io_diffCommits_info_241_rfWen = RTL_PATH.io_diffCommits_info_241_rfWen; \
        force U_IF_NAME.io_diffCommits_info_241_fpWen = RTL_PATH.io_diffCommits_info_241_fpWen; \
        force U_IF_NAME.io_diffCommits_info_241_vecWen = RTL_PATH.io_diffCommits_info_241_vecWen; \
        force U_IF_NAME.io_diffCommits_info_241_v0Wen = RTL_PATH.io_diffCommits_info_241_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_241_vlWen = RTL_PATH.io_diffCommits_info_241_vlWen; \
        force U_IF_NAME.io_diffCommits_info_242_ldest = RTL_PATH.io_diffCommits_info_242_ldest; \
        force U_IF_NAME.io_diffCommits_info_242_pdest = RTL_PATH.io_diffCommits_info_242_pdest; \
        force U_IF_NAME.io_diffCommits_info_242_rfWen = RTL_PATH.io_diffCommits_info_242_rfWen; \
        force U_IF_NAME.io_diffCommits_info_242_fpWen = RTL_PATH.io_diffCommits_info_242_fpWen; \
        force U_IF_NAME.io_diffCommits_info_242_vecWen = RTL_PATH.io_diffCommits_info_242_vecWen; \
        force U_IF_NAME.io_diffCommits_info_242_v0Wen = RTL_PATH.io_diffCommits_info_242_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_242_vlWen = RTL_PATH.io_diffCommits_info_242_vlWen; \
        force U_IF_NAME.io_diffCommits_info_243_ldest = RTL_PATH.io_diffCommits_info_243_ldest; \
        force U_IF_NAME.io_diffCommits_info_243_pdest = RTL_PATH.io_diffCommits_info_243_pdest; \
        force U_IF_NAME.io_diffCommits_info_243_rfWen = RTL_PATH.io_diffCommits_info_243_rfWen; \
        force U_IF_NAME.io_diffCommits_info_243_fpWen = RTL_PATH.io_diffCommits_info_243_fpWen; \
        force U_IF_NAME.io_diffCommits_info_243_vecWen = RTL_PATH.io_diffCommits_info_243_vecWen; \
        force U_IF_NAME.io_diffCommits_info_243_v0Wen = RTL_PATH.io_diffCommits_info_243_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_243_vlWen = RTL_PATH.io_diffCommits_info_243_vlWen; \
        force U_IF_NAME.io_diffCommits_info_244_ldest = RTL_PATH.io_diffCommits_info_244_ldest; \
        force U_IF_NAME.io_diffCommits_info_244_pdest = RTL_PATH.io_diffCommits_info_244_pdest; \
        force U_IF_NAME.io_diffCommits_info_244_rfWen = RTL_PATH.io_diffCommits_info_244_rfWen; \
        force U_IF_NAME.io_diffCommits_info_244_fpWen = RTL_PATH.io_diffCommits_info_244_fpWen; \
        force U_IF_NAME.io_diffCommits_info_244_vecWen = RTL_PATH.io_diffCommits_info_244_vecWen; \
        force U_IF_NAME.io_diffCommits_info_244_v0Wen = RTL_PATH.io_diffCommits_info_244_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_244_vlWen = RTL_PATH.io_diffCommits_info_244_vlWen; \
        force U_IF_NAME.io_diffCommits_info_245_ldest = RTL_PATH.io_diffCommits_info_245_ldest; \
        force U_IF_NAME.io_diffCommits_info_245_pdest = RTL_PATH.io_diffCommits_info_245_pdest; \
        force U_IF_NAME.io_diffCommits_info_245_rfWen = RTL_PATH.io_diffCommits_info_245_rfWen; \
        force U_IF_NAME.io_diffCommits_info_245_fpWen = RTL_PATH.io_diffCommits_info_245_fpWen; \
        force U_IF_NAME.io_diffCommits_info_245_vecWen = RTL_PATH.io_diffCommits_info_245_vecWen; \
        force U_IF_NAME.io_diffCommits_info_245_v0Wen = RTL_PATH.io_diffCommits_info_245_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_245_vlWen = RTL_PATH.io_diffCommits_info_245_vlWen; \
        force U_IF_NAME.io_diffCommits_info_246_ldest = RTL_PATH.io_diffCommits_info_246_ldest; \
        force U_IF_NAME.io_diffCommits_info_246_pdest = RTL_PATH.io_diffCommits_info_246_pdest; \
        force U_IF_NAME.io_diffCommits_info_246_rfWen = RTL_PATH.io_diffCommits_info_246_rfWen; \
        force U_IF_NAME.io_diffCommits_info_246_fpWen = RTL_PATH.io_diffCommits_info_246_fpWen; \
        force U_IF_NAME.io_diffCommits_info_246_vecWen = RTL_PATH.io_diffCommits_info_246_vecWen; \
        force U_IF_NAME.io_diffCommits_info_246_v0Wen = RTL_PATH.io_diffCommits_info_246_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_246_vlWen = RTL_PATH.io_diffCommits_info_246_vlWen; \
        force U_IF_NAME.io_diffCommits_info_247_ldest = RTL_PATH.io_diffCommits_info_247_ldest; \
        force U_IF_NAME.io_diffCommits_info_247_pdest = RTL_PATH.io_diffCommits_info_247_pdest; \
        force U_IF_NAME.io_diffCommits_info_247_rfWen = RTL_PATH.io_diffCommits_info_247_rfWen; \
        force U_IF_NAME.io_diffCommits_info_247_fpWen = RTL_PATH.io_diffCommits_info_247_fpWen; \
        force U_IF_NAME.io_diffCommits_info_247_vecWen = RTL_PATH.io_diffCommits_info_247_vecWen; \
        force U_IF_NAME.io_diffCommits_info_247_v0Wen = RTL_PATH.io_diffCommits_info_247_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_247_vlWen = RTL_PATH.io_diffCommits_info_247_vlWen; \
        force U_IF_NAME.io_diffCommits_info_248_ldest = RTL_PATH.io_diffCommits_info_248_ldest; \
        force U_IF_NAME.io_diffCommits_info_248_pdest = RTL_PATH.io_diffCommits_info_248_pdest; \
        force U_IF_NAME.io_diffCommits_info_248_rfWen = RTL_PATH.io_diffCommits_info_248_rfWen; \
        force U_IF_NAME.io_diffCommits_info_248_fpWen = RTL_PATH.io_diffCommits_info_248_fpWen; \
        force U_IF_NAME.io_diffCommits_info_248_vecWen = RTL_PATH.io_diffCommits_info_248_vecWen; \
        force U_IF_NAME.io_diffCommits_info_248_v0Wen = RTL_PATH.io_diffCommits_info_248_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_248_vlWen = RTL_PATH.io_diffCommits_info_248_vlWen; \
        force U_IF_NAME.io_diffCommits_info_249_ldest = RTL_PATH.io_diffCommits_info_249_ldest; \
        force U_IF_NAME.io_diffCommits_info_249_pdest = RTL_PATH.io_diffCommits_info_249_pdest; \
        force U_IF_NAME.io_diffCommits_info_249_rfWen = RTL_PATH.io_diffCommits_info_249_rfWen; \
        force U_IF_NAME.io_diffCommits_info_249_fpWen = RTL_PATH.io_diffCommits_info_249_fpWen; \
        force U_IF_NAME.io_diffCommits_info_249_vecWen = RTL_PATH.io_diffCommits_info_249_vecWen; \
        force U_IF_NAME.io_diffCommits_info_249_v0Wen = RTL_PATH.io_diffCommits_info_249_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_249_vlWen = RTL_PATH.io_diffCommits_info_249_vlWen; \
        force U_IF_NAME.io_diffCommits_info_250_ldest = RTL_PATH.io_diffCommits_info_250_ldest; \
        force U_IF_NAME.io_diffCommits_info_250_pdest = RTL_PATH.io_diffCommits_info_250_pdest; \
        force U_IF_NAME.io_diffCommits_info_250_rfWen = RTL_PATH.io_diffCommits_info_250_rfWen; \
        force U_IF_NAME.io_diffCommits_info_250_fpWen = RTL_PATH.io_diffCommits_info_250_fpWen; \
        force U_IF_NAME.io_diffCommits_info_250_vecWen = RTL_PATH.io_diffCommits_info_250_vecWen; \
        force U_IF_NAME.io_diffCommits_info_250_v0Wen = RTL_PATH.io_diffCommits_info_250_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_250_vlWen = RTL_PATH.io_diffCommits_info_250_vlWen; \
        force U_IF_NAME.io_diffCommits_info_251_ldest = RTL_PATH.io_diffCommits_info_251_ldest; \
        force U_IF_NAME.io_diffCommits_info_251_pdest = RTL_PATH.io_diffCommits_info_251_pdest; \
        force U_IF_NAME.io_diffCommits_info_251_rfWen = RTL_PATH.io_diffCommits_info_251_rfWen; \
        force U_IF_NAME.io_diffCommits_info_251_fpWen = RTL_PATH.io_diffCommits_info_251_fpWen; \
        force U_IF_NAME.io_diffCommits_info_251_vecWen = RTL_PATH.io_diffCommits_info_251_vecWen; \
        force U_IF_NAME.io_diffCommits_info_251_v0Wen = RTL_PATH.io_diffCommits_info_251_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_251_vlWen = RTL_PATH.io_diffCommits_info_251_vlWen; \
        force U_IF_NAME.io_diffCommits_info_252_ldest = RTL_PATH.io_diffCommits_info_252_ldest; \
        force U_IF_NAME.io_diffCommits_info_252_pdest = RTL_PATH.io_diffCommits_info_252_pdest; \
        force U_IF_NAME.io_diffCommits_info_252_rfWen = RTL_PATH.io_diffCommits_info_252_rfWen; \
        force U_IF_NAME.io_diffCommits_info_252_fpWen = RTL_PATH.io_diffCommits_info_252_fpWen; \
        force U_IF_NAME.io_diffCommits_info_252_vecWen = RTL_PATH.io_diffCommits_info_252_vecWen; \
        force U_IF_NAME.io_diffCommits_info_252_v0Wen = RTL_PATH.io_diffCommits_info_252_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_252_vlWen = RTL_PATH.io_diffCommits_info_252_vlWen; \
        force U_IF_NAME.io_diffCommits_info_253_ldest = RTL_PATH.io_diffCommits_info_253_ldest; \
        force U_IF_NAME.io_diffCommits_info_253_pdest = RTL_PATH.io_diffCommits_info_253_pdest; \
        force U_IF_NAME.io_diffCommits_info_253_rfWen = RTL_PATH.io_diffCommits_info_253_rfWen; \
        force U_IF_NAME.io_diffCommits_info_253_fpWen = RTL_PATH.io_diffCommits_info_253_fpWen; \
        force U_IF_NAME.io_diffCommits_info_253_vecWen = RTL_PATH.io_diffCommits_info_253_vecWen; \
        force U_IF_NAME.io_diffCommits_info_253_v0Wen = RTL_PATH.io_diffCommits_info_253_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_253_vlWen = RTL_PATH.io_diffCommits_info_253_vlWen; \
        force U_IF_NAME.io_diffCommits_info_254_ldest = RTL_PATH.io_diffCommits_info_254_ldest; \
        force U_IF_NAME.io_diffCommits_info_254_pdest = RTL_PATH.io_diffCommits_info_254_pdest; \
        force U_IF_NAME.io_diffCommits_info_254_rfWen = RTL_PATH.io_diffCommits_info_254_rfWen; \
        force U_IF_NAME.io_diffCommits_info_254_fpWen = RTL_PATH.io_diffCommits_info_254_fpWen; \
        force U_IF_NAME.io_diffCommits_info_254_vecWen = RTL_PATH.io_diffCommits_info_254_vecWen; \
        force U_IF_NAME.io_diffCommits_info_254_v0Wen = RTL_PATH.io_diffCommits_info_254_v0Wen; \
        force U_IF_NAME.io_diffCommits_info_254_vlWen = RTL_PATH.io_diffCommits_info_254_vlWen; \
        force U_IF_NAME.io_diffCommits_info_255_ldest = RTL_PATH.io_diffCommits_info_255_ldest; \
        force U_IF_NAME.io_diffCommits_info_255_pdest = RTL_PATH.io_diffCommits_info_255_pdest; \
        force U_IF_NAME.io_diffCommits_info_256_ldest = RTL_PATH.io_diffCommits_info_256_ldest; \
        force U_IF_NAME.io_diffCommits_info_256_pdest = RTL_PATH.io_diffCommits_info_256_pdest; \
        force U_IF_NAME.io_diffCommits_info_257_ldest = RTL_PATH.io_diffCommits_info_257_ldest; \
        force U_IF_NAME.io_diffCommits_info_257_pdest = RTL_PATH.io_diffCommits_info_257_pdest; \
        force U_IF_NAME.io_diffCommits_info_258_ldest = RTL_PATH.io_diffCommits_info_258_ldest; \
        force U_IF_NAME.io_diffCommits_info_258_pdest = RTL_PATH.io_diffCommits_info_258_pdest; \
        force U_IF_NAME.io_diffCommits_info_259_ldest = RTL_PATH.io_diffCommits_info_259_ldest; \
        force U_IF_NAME.io_diffCommits_info_259_pdest = RTL_PATH.io_diffCommits_info_259_pdest; \
        force U_IF_NAME.io_diffCommits_info_260_ldest = RTL_PATH.io_diffCommits_info_260_ldest; \
        force U_IF_NAME.io_diffCommits_info_260_pdest = RTL_PATH.io_diffCommits_info_260_pdest; \
        force U_IF_NAME.io_diffCommits_info_261_ldest = RTL_PATH.io_diffCommits_info_261_ldest; \
        force U_IF_NAME.io_diffCommits_info_261_pdest = RTL_PATH.io_diffCommits_info_261_pdest; \
        force U_IF_NAME.io_diffCommits_info_262_ldest = RTL_PATH.io_diffCommits_info_262_ldest; \
        force U_IF_NAME.io_diffCommits_info_262_pdest = RTL_PATH.io_diffCommits_info_262_pdest; \
        force U_IF_NAME.io_diffCommits_info_263_ldest = RTL_PATH.io_diffCommits_info_263_ldest; \
        force U_IF_NAME.io_diffCommits_info_263_pdest = RTL_PATH.io_diffCommits_info_263_pdest; \
        force U_IF_NAME.io_diffCommits_info_264_ldest = RTL_PATH.io_diffCommits_info_264_ldest; \
        force U_IF_NAME.io_diffCommits_info_264_pdest = RTL_PATH.io_diffCommits_info_264_pdest; \
        force U_IF_NAME.io_diffCommits_info_265_ldest = RTL_PATH.io_diffCommits_info_265_ldest; \
        force U_IF_NAME.io_diffCommits_info_265_pdest = RTL_PATH.io_diffCommits_info_265_pdest; \
        force U_IF_NAME.io_diffCommits_info_266_ldest = RTL_PATH.io_diffCommits_info_266_ldest; \
        force U_IF_NAME.io_diffCommits_info_266_pdest = RTL_PATH.io_diffCommits_info_266_pdest; \
        force U_IF_NAME.io_diffCommits_info_267_ldest = RTL_PATH.io_diffCommits_info_267_ldest; \
        force U_IF_NAME.io_diffCommits_info_267_pdest = RTL_PATH.io_diffCommits_info_267_pdest; \
        force U_IF_NAME.io_diffCommits_info_268_ldest = RTL_PATH.io_diffCommits_info_268_ldest; \
        force U_IF_NAME.io_diffCommits_info_268_pdest = RTL_PATH.io_diffCommits_info_268_pdest; \
        force U_IF_NAME.io_diffCommits_info_269_ldest = RTL_PATH.io_diffCommits_info_269_ldest; \
        force U_IF_NAME.io_diffCommits_info_269_pdest = RTL_PATH.io_diffCommits_info_269_pdest; \
        force U_IF_NAME.io_diffCommits_info_270_ldest = RTL_PATH.io_diffCommits_info_270_ldest; \
        force U_IF_NAME.io_diffCommits_info_270_pdest = RTL_PATH.io_diffCommits_info_270_pdest; \
        force U_IF_NAME.io_diffCommits_info_271_ldest = RTL_PATH.io_diffCommits_info_271_ldest; \
        force U_IF_NAME.io_diffCommits_info_271_pdest = RTL_PATH.io_diffCommits_info_271_pdest; \
        force U_IF_NAME.io_diffCommits_info_272_ldest = RTL_PATH.io_diffCommits_info_272_ldest; \
        force U_IF_NAME.io_diffCommits_info_272_pdest = RTL_PATH.io_diffCommits_info_272_pdest; \
        force U_IF_NAME.io_diffCommits_info_273_ldest = RTL_PATH.io_diffCommits_info_273_ldest; \
        force U_IF_NAME.io_diffCommits_info_273_pdest = RTL_PATH.io_diffCommits_info_273_pdest; \
        force U_IF_NAME.io_diffCommits_info_274_ldest = RTL_PATH.io_diffCommits_info_274_ldest; \
        force U_IF_NAME.io_diffCommits_info_274_pdest = RTL_PATH.io_diffCommits_info_274_pdest; \
        force U_IF_NAME.io_diffCommits_info_275_ldest = RTL_PATH.io_diffCommits_info_275_ldest; \
        force U_IF_NAME.io_diffCommits_info_275_pdest = RTL_PATH.io_diffCommits_info_275_pdest; \
        force U_IF_NAME.io_diffCommits_info_276_ldest = RTL_PATH.io_diffCommits_info_276_ldest; \
        force U_IF_NAME.io_diffCommits_info_276_pdest = RTL_PATH.io_diffCommits_info_276_pdest; \
        force U_IF_NAME.io_diffCommits_info_277_ldest = RTL_PATH.io_diffCommits_info_277_ldest; \
        force U_IF_NAME.io_diffCommits_info_277_pdest = RTL_PATH.io_diffCommits_info_277_pdest; \
        force U_IF_NAME.io_diffCommits_info_278_ldest = RTL_PATH.io_diffCommits_info_278_ldest; \
        force U_IF_NAME.io_diffCommits_info_278_pdest = RTL_PATH.io_diffCommits_info_278_pdest; \
        force U_IF_NAME.io_diffCommits_info_279_ldest = RTL_PATH.io_diffCommits_info_279_ldest; \
        force U_IF_NAME.io_diffCommits_info_279_pdest = RTL_PATH.io_diffCommits_info_279_pdest; \
        force U_IF_NAME.io_diffCommits_info_280_ldest = RTL_PATH.io_diffCommits_info_280_ldest; \
        force U_IF_NAME.io_diffCommits_info_280_pdest = RTL_PATH.io_diffCommits_info_280_pdest; \
        force U_IF_NAME.io_diffCommits_info_281_ldest = RTL_PATH.io_diffCommits_info_281_ldest; \
        force U_IF_NAME.io_diffCommits_info_281_pdest = RTL_PATH.io_diffCommits_info_281_pdest; \
        force U_IF_NAME.io_diffCommits_info_282_ldest = RTL_PATH.io_diffCommits_info_282_ldest; \
        force U_IF_NAME.io_diffCommits_info_282_pdest = RTL_PATH.io_diffCommits_info_282_pdest; \
        force U_IF_NAME.io_diffCommits_info_283_ldest = RTL_PATH.io_diffCommits_info_283_ldest; \
        force U_IF_NAME.io_diffCommits_info_283_pdest = RTL_PATH.io_diffCommits_info_283_pdest; \
        force U_IF_NAME.io_diffCommits_info_284_ldest = RTL_PATH.io_diffCommits_info_284_ldest; \
        force U_IF_NAME.io_diffCommits_info_284_pdest = RTL_PATH.io_diffCommits_info_284_pdest; \
        force U_IF_NAME.io_diffCommits_info_285_ldest = RTL_PATH.io_diffCommits_info_285_ldest; \
        force U_IF_NAME.io_diffCommits_info_285_pdest = RTL_PATH.io_diffCommits_info_285_pdest; \
        force U_IF_NAME.io_diffCommits_info_286_ldest = RTL_PATH.io_diffCommits_info_286_ldest; \
        force U_IF_NAME.io_diffCommits_info_286_pdest = RTL_PATH.io_diffCommits_info_286_pdest; \
        force U_IF_NAME.io_diffCommits_info_287_ldest = RTL_PATH.io_diffCommits_info_287_ldest; \
        force U_IF_NAME.io_diffCommits_info_287_pdest = RTL_PATH.io_diffCommits_info_287_pdest; \
        force U_IF_NAME.io_diffCommits_info_288_ldest = RTL_PATH.io_diffCommits_info_288_ldest; \
        force U_IF_NAME.io_diffCommits_info_288_pdest = RTL_PATH.io_diffCommits_info_288_pdest; \
        force U_IF_NAME.io_diffCommits_info_289_ldest = RTL_PATH.io_diffCommits_info_289_ldest; \
        force U_IF_NAME.io_diffCommits_info_289_pdest = RTL_PATH.io_diffCommits_info_289_pdest; \
        force U_IF_NAME.io_diffCommits_info_290_ldest = RTL_PATH.io_diffCommits_info_290_ldest; \
        force U_IF_NAME.io_diffCommits_info_290_pdest = RTL_PATH.io_diffCommits_info_290_pdest; \
        force U_IF_NAME.io_diffCommits_info_291_ldest = RTL_PATH.io_diffCommits_info_291_ldest; \
        force U_IF_NAME.io_diffCommits_info_291_pdest = RTL_PATH.io_diffCommits_info_291_pdest; \
        force U_IF_NAME.io_diffCommits_info_292_ldest = RTL_PATH.io_diffCommits_info_292_ldest; \
        force U_IF_NAME.io_diffCommits_info_292_pdest = RTL_PATH.io_diffCommits_info_292_pdest; \
        force U_IF_NAME.io_diffCommits_info_293_ldest = RTL_PATH.io_diffCommits_info_293_ldest; \
        force U_IF_NAME.io_diffCommits_info_293_pdest = RTL_PATH.io_diffCommits_info_293_pdest; \
        force U_IF_NAME.io_diffCommits_info_294_ldest = RTL_PATH.io_diffCommits_info_294_ldest; \
        force U_IF_NAME.io_diffCommits_info_294_pdest = RTL_PATH.io_diffCommits_info_294_pdest; \
        force U_IF_NAME.io_diffCommits_info_295_ldest = RTL_PATH.io_diffCommits_info_295_ldest; \
        force U_IF_NAME.io_diffCommits_info_295_pdest = RTL_PATH.io_diffCommits_info_295_pdest; \
        force U_IF_NAME.io_diffCommits_info_296_ldest = RTL_PATH.io_diffCommits_info_296_ldest; \
        force U_IF_NAME.io_diffCommits_info_296_pdest = RTL_PATH.io_diffCommits_info_296_pdest; \
        force U_IF_NAME.io_diffCommits_info_297_ldest = RTL_PATH.io_diffCommits_info_297_ldest; \
        force U_IF_NAME.io_diffCommits_info_297_pdest = RTL_PATH.io_diffCommits_info_297_pdest; \
        force U_IF_NAME.io_diffCommits_info_298_ldest = RTL_PATH.io_diffCommits_info_298_ldest; \
        force U_IF_NAME.io_diffCommits_info_298_pdest = RTL_PATH.io_diffCommits_info_298_pdest; \
        force U_IF_NAME.io_diffCommits_info_299_ldest = RTL_PATH.io_diffCommits_info_299_ldest; \
        force U_IF_NAME.io_diffCommits_info_299_pdest = RTL_PATH.io_diffCommits_info_299_pdest; \
        force U_IF_NAME.io_diffCommits_info_300_ldest = RTL_PATH.io_diffCommits_info_300_ldest; \
        force U_IF_NAME.io_diffCommits_info_300_pdest = RTL_PATH.io_diffCommits_info_300_pdest; \
        force U_IF_NAME.io_diffCommits_info_301_ldest = RTL_PATH.io_diffCommits_info_301_ldest; \
        force U_IF_NAME.io_diffCommits_info_301_pdest = RTL_PATH.io_diffCommits_info_301_pdest; \
        force U_IF_NAME.io_diffCommits_info_302_ldest = RTL_PATH.io_diffCommits_info_302_ldest; \
        force U_IF_NAME.io_diffCommits_info_302_pdest = RTL_PATH.io_diffCommits_info_302_pdest; \
        force U_IF_NAME.io_diffCommits_info_303_ldest = RTL_PATH.io_diffCommits_info_303_ldest; \
        force U_IF_NAME.io_diffCommits_info_303_pdest = RTL_PATH.io_diffCommits_info_303_pdest; \
        force U_IF_NAME.io_diffCommits_info_304_ldest = RTL_PATH.io_diffCommits_info_304_ldest; \
        force U_IF_NAME.io_diffCommits_info_304_pdest = RTL_PATH.io_diffCommits_info_304_pdest; \
        force U_IF_NAME.io_diffCommits_info_305_ldest = RTL_PATH.io_diffCommits_info_305_ldest; \
        force U_IF_NAME.io_diffCommits_info_305_pdest = RTL_PATH.io_diffCommits_info_305_pdest; \
        force U_IF_NAME.io_diffCommits_info_306_ldest = RTL_PATH.io_diffCommits_info_306_ldest; \
        force U_IF_NAME.io_diffCommits_info_306_pdest = RTL_PATH.io_diffCommits_info_306_pdest; \
        force U_IF_NAME.io_diffCommits_info_307_ldest = RTL_PATH.io_diffCommits_info_307_ldest; \
        force U_IF_NAME.io_diffCommits_info_307_pdest = RTL_PATH.io_diffCommits_info_307_pdest; \
        force U_IF_NAME.io_diffCommits_info_308_ldest = RTL_PATH.io_diffCommits_info_308_ldest; \
        force U_IF_NAME.io_diffCommits_info_308_pdest = RTL_PATH.io_diffCommits_info_308_pdest; \
        force U_IF_NAME.io_diffCommits_info_309_ldest = RTL_PATH.io_diffCommits_info_309_ldest; \
        force U_IF_NAME.io_diffCommits_info_309_pdest = RTL_PATH.io_diffCommits_info_309_pdest; \
        force U_IF_NAME.io_diffCommits_info_310_ldest = RTL_PATH.io_diffCommits_info_310_ldest; \
        force U_IF_NAME.io_diffCommits_info_310_pdest = RTL_PATH.io_diffCommits_info_310_pdest; \
        force U_IF_NAME.io_diffCommits_info_311_ldest = RTL_PATH.io_diffCommits_info_311_ldest; \
        force U_IF_NAME.io_diffCommits_info_311_pdest = RTL_PATH.io_diffCommits_info_311_pdest; \
        force U_IF_NAME.io_diffCommits_info_312_ldest = RTL_PATH.io_diffCommits_info_312_ldest; \
        force U_IF_NAME.io_diffCommits_info_312_pdest = RTL_PATH.io_diffCommits_info_312_pdest; \
        force U_IF_NAME.io_diffCommits_info_313_ldest = RTL_PATH.io_diffCommits_info_313_ldest; \
        force U_IF_NAME.io_diffCommits_info_313_pdest = RTL_PATH.io_diffCommits_info_313_pdest; \
        force U_IF_NAME.io_diffCommits_info_314_ldest = RTL_PATH.io_diffCommits_info_314_ldest; \
        force U_IF_NAME.io_diffCommits_info_314_pdest = RTL_PATH.io_diffCommits_info_314_pdest; \
        force U_IF_NAME.io_diffCommits_info_315_ldest = RTL_PATH.io_diffCommits_info_315_ldest; \
        force U_IF_NAME.io_diffCommits_info_315_pdest = RTL_PATH.io_diffCommits_info_315_pdest; \
        force U_IF_NAME.io_diffCommits_info_316_ldest = RTL_PATH.io_diffCommits_info_316_ldest; \
        force U_IF_NAME.io_diffCommits_info_316_pdest = RTL_PATH.io_diffCommits_info_316_pdest; \
        force U_IF_NAME.io_diffCommits_info_317_ldest = RTL_PATH.io_diffCommits_info_317_ldest; \
        force U_IF_NAME.io_diffCommits_info_317_pdest = RTL_PATH.io_diffCommits_info_317_pdest; \
        force U_IF_NAME.io_diffCommits_info_318_ldest = RTL_PATH.io_diffCommits_info_318_ldest; \
        force U_IF_NAME.io_diffCommits_info_318_pdest = RTL_PATH.io_diffCommits_info_318_pdest; \
        force U_IF_NAME.io_diffCommits_info_319_ldest = RTL_PATH.io_diffCommits_info_319_ldest; \
        force U_IF_NAME.io_diffCommits_info_319_pdest = RTL_PATH.io_diffCommits_info_319_pdest; \
        force U_IF_NAME.io_diffCommits_info_320_ldest = RTL_PATH.io_diffCommits_info_320_ldest; \
        force U_IF_NAME.io_diffCommits_info_320_pdest = RTL_PATH.io_diffCommits_info_320_pdest; \
        force U_IF_NAME.io_diffCommits_info_321_ldest = RTL_PATH.io_diffCommits_info_321_ldest; \
        force U_IF_NAME.io_diffCommits_info_321_pdest = RTL_PATH.io_diffCommits_info_321_pdest; \
        force U_IF_NAME.io_diffCommits_info_322_ldest = RTL_PATH.io_diffCommits_info_322_ldest; \
        force U_IF_NAME.io_diffCommits_info_322_pdest = RTL_PATH.io_diffCommits_info_322_pdest; \
        force U_IF_NAME.io_diffCommits_info_323_ldest = RTL_PATH.io_diffCommits_info_323_ldest; \
        force U_IF_NAME.io_diffCommits_info_323_pdest = RTL_PATH.io_diffCommits_info_323_pdest; \
        force U_IF_NAME.io_diffCommits_info_324_ldest = RTL_PATH.io_diffCommits_info_324_ldest; \
        force U_IF_NAME.io_diffCommits_info_324_pdest = RTL_PATH.io_diffCommits_info_324_pdest; \
        force U_IF_NAME.io_diffCommits_info_325_ldest = RTL_PATH.io_diffCommits_info_325_ldest; \
        force U_IF_NAME.io_diffCommits_info_325_pdest = RTL_PATH.io_diffCommits_info_325_pdest; \
        force U_IF_NAME.io_diffCommits_info_326_ldest = RTL_PATH.io_diffCommits_info_326_ldest; \
        force U_IF_NAME.io_diffCommits_info_326_pdest = RTL_PATH.io_diffCommits_info_326_pdest; \
        force U_IF_NAME.io_diffCommits_info_327_ldest = RTL_PATH.io_diffCommits_info_327_ldest; \
        force U_IF_NAME.io_diffCommits_info_327_pdest = RTL_PATH.io_diffCommits_info_327_pdest; \
        force U_IF_NAME.io_diffCommits_info_328_ldest = RTL_PATH.io_diffCommits_info_328_ldest; \
        force U_IF_NAME.io_diffCommits_info_328_pdest = RTL_PATH.io_diffCommits_info_328_pdest; \
        force U_IF_NAME.io_diffCommits_info_329_ldest = RTL_PATH.io_diffCommits_info_329_ldest; \
        force U_IF_NAME.io_diffCommits_info_329_pdest = RTL_PATH.io_diffCommits_info_329_pdest; \
        force U_IF_NAME.io_diffCommits_info_330_ldest = RTL_PATH.io_diffCommits_info_330_ldest; \
        force U_IF_NAME.io_diffCommits_info_330_pdest = RTL_PATH.io_diffCommits_info_330_pdest; \
        force U_IF_NAME.io_diffCommits_info_331_ldest = RTL_PATH.io_diffCommits_info_331_ldest; \
        force U_IF_NAME.io_diffCommits_info_331_pdest = RTL_PATH.io_diffCommits_info_331_pdest; \
        force U_IF_NAME.io_diffCommits_info_332_ldest = RTL_PATH.io_diffCommits_info_332_ldest; \
        force U_IF_NAME.io_diffCommits_info_332_pdest = RTL_PATH.io_diffCommits_info_332_pdest; \
        force U_IF_NAME.io_diffCommits_info_333_ldest = RTL_PATH.io_diffCommits_info_333_ldest; \
        force U_IF_NAME.io_diffCommits_info_333_pdest = RTL_PATH.io_diffCommits_info_333_pdest; \
        force U_IF_NAME.io_diffCommits_info_334_ldest = RTL_PATH.io_diffCommits_info_334_ldest; \
        force U_IF_NAME.io_diffCommits_info_334_pdest = RTL_PATH.io_diffCommits_info_334_pdest; \
        force U_IF_NAME.io_diffCommits_info_335_ldest = RTL_PATH.io_diffCommits_info_335_ldest; \
        force U_IF_NAME.io_diffCommits_info_335_pdest = RTL_PATH.io_diffCommits_info_335_pdest; \
        force U_IF_NAME.io_diffCommits_info_336_ldest = RTL_PATH.io_diffCommits_info_336_ldest; \
        force U_IF_NAME.io_diffCommits_info_336_pdest = RTL_PATH.io_diffCommits_info_336_pdest; \
        force U_IF_NAME.io_diffCommits_info_337_ldest = RTL_PATH.io_diffCommits_info_337_ldest; \
        force U_IF_NAME.io_diffCommits_info_337_pdest = RTL_PATH.io_diffCommits_info_337_pdest; \
        force U_IF_NAME.io_diffCommits_info_338_ldest = RTL_PATH.io_diffCommits_info_338_ldest; \
        force U_IF_NAME.io_diffCommits_info_338_pdest = RTL_PATH.io_diffCommits_info_338_pdest; \
        force U_IF_NAME.io_diffCommits_info_339_ldest = RTL_PATH.io_diffCommits_info_339_ldest; \
        force U_IF_NAME.io_diffCommits_info_339_pdest = RTL_PATH.io_diffCommits_info_339_pdest; \
        force U_IF_NAME.io_diffCommits_info_340_ldest = RTL_PATH.io_diffCommits_info_340_ldest; \
        force U_IF_NAME.io_diffCommits_info_340_pdest = RTL_PATH.io_diffCommits_info_340_pdest; \
        force U_IF_NAME.io_diffCommits_info_341_ldest = RTL_PATH.io_diffCommits_info_341_ldest; \
        force U_IF_NAME.io_diffCommits_info_341_pdest = RTL_PATH.io_diffCommits_info_341_pdest; \
        force U_IF_NAME.io_diffCommits_info_342_ldest = RTL_PATH.io_diffCommits_info_342_ldest; \
        force U_IF_NAME.io_diffCommits_info_342_pdest = RTL_PATH.io_diffCommits_info_342_pdest; \
        force U_IF_NAME.io_diffCommits_info_343_ldest = RTL_PATH.io_diffCommits_info_343_ldest; \
        force U_IF_NAME.io_diffCommits_info_343_pdest = RTL_PATH.io_diffCommits_info_343_pdest; \
        force U_IF_NAME.io_diffCommits_info_344_ldest = RTL_PATH.io_diffCommits_info_344_ldest; \
        force U_IF_NAME.io_diffCommits_info_344_pdest = RTL_PATH.io_diffCommits_info_344_pdest; \
        force U_IF_NAME.io_diffCommits_info_345_ldest = RTL_PATH.io_diffCommits_info_345_ldest; \
        force U_IF_NAME.io_diffCommits_info_345_pdest = RTL_PATH.io_diffCommits_info_345_pdest; \
        force U_IF_NAME.io_diffCommits_info_346_ldest = RTL_PATH.io_diffCommits_info_346_ldest; \
        force U_IF_NAME.io_diffCommits_info_346_pdest = RTL_PATH.io_diffCommits_info_346_pdest; \
        force U_IF_NAME.io_diffCommits_info_347_ldest = RTL_PATH.io_diffCommits_info_347_ldest; \
        force U_IF_NAME.io_diffCommits_info_347_pdest = RTL_PATH.io_diffCommits_info_347_pdest; \
        force U_IF_NAME.io_diffCommits_info_348_ldest = RTL_PATH.io_diffCommits_info_348_ldest; \
        force U_IF_NAME.io_diffCommits_info_348_pdest = RTL_PATH.io_diffCommits_info_348_pdest; \
        force U_IF_NAME.io_diffCommits_info_349_ldest = RTL_PATH.io_diffCommits_info_349_ldest; \
        force U_IF_NAME.io_diffCommits_info_349_pdest = RTL_PATH.io_diffCommits_info_349_pdest; \
        force U_IF_NAME.io_diffCommits_info_350_ldest = RTL_PATH.io_diffCommits_info_350_ldest; \
        force U_IF_NAME.io_diffCommits_info_350_pdest = RTL_PATH.io_diffCommits_info_350_pdest; \
        force U_IF_NAME.io_diffCommits_info_351_ldest = RTL_PATH.io_diffCommits_info_351_ldest; \
        force U_IF_NAME.io_diffCommits_info_351_pdest = RTL_PATH.io_diffCommits_info_351_pdest; \
        force U_IF_NAME.io_diffCommits_info_352_ldest = RTL_PATH.io_diffCommits_info_352_ldest; \
        force U_IF_NAME.io_diffCommits_info_352_pdest = RTL_PATH.io_diffCommits_info_352_pdest; \
        force U_IF_NAME.io_diffCommits_info_353_ldest = RTL_PATH.io_diffCommits_info_353_ldest; \
        force U_IF_NAME.io_diffCommits_info_353_pdest = RTL_PATH.io_diffCommits_info_353_pdest; \
        force U_IF_NAME.io_diffCommits_info_354_ldest = RTL_PATH.io_diffCommits_info_354_ldest; \
        force U_IF_NAME.io_diffCommits_info_354_pdest = RTL_PATH.io_diffCommits_info_354_pdest; \
        force U_IF_NAME.io_diffCommits_info_355_ldest = RTL_PATH.io_diffCommits_info_355_ldest; \
        force U_IF_NAME.io_diffCommits_info_355_pdest = RTL_PATH.io_diffCommits_info_355_pdest; \
        force U_IF_NAME.io_diffCommits_info_356_ldest = RTL_PATH.io_diffCommits_info_356_ldest; \
        force U_IF_NAME.io_diffCommits_info_356_pdest = RTL_PATH.io_diffCommits_info_356_pdest; \
        force U_IF_NAME.io_diffCommits_info_357_ldest = RTL_PATH.io_diffCommits_info_357_ldest; \
        force U_IF_NAME.io_diffCommits_info_357_pdest = RTL_PATH.io_diffCommits_info_357_pdest; \
        force U_IF_NAME.io_diffCommits_info_358_ldest = RTL_PATH.io_diffCommits_info_358_ldest; \
        force U_IF_NAME.io_diffCommits_info_358_pdest = RTL_PATH.io_diffCommits_info_358_pdest; \
        force U_IF_NAME.io_diffCommits_info_359_ldest = RTL_PATH.io_diffCommits_info_359_ldest; \
        force U_IF_NAME.io_diffCommits_info_359_pdest = RTL_PATH.io_diffCommits_info_359_pdest; \
        force U_IF_NAME.io_diffCommits_info_360_ldest = RTL_PATH.io_diffCommits_info_360_ldest; \
        force U_IF_NAME.io_diffCommits_info_360_pdest = RTL_PATH.io_diffCommits_info_360_pdest; \
        force U_IF_NAME.io_diffCommits_info_361_ldest = RTL_PATH.io_diffCommits_info_361_ldest; \
        force U_IF_NAME.io_diffCommits_info_361_pdest = RTL_PATH.io_diffCommits_info_361_pdest; \
        force U_IF_NAME.io_diffCommits_info_362_ldest = RTL_PATH.io_diffCommits_info_362_ldest; \
        force U_IF_NAME.io_diffCommits_info_362_pdest = RTL_PATH.io_diffCommits_info_362_pdest; \
        force U_IF_NAME.io_diffCommits_info_363_ldest = RTL_PATH.io_diffCommits_info_363_ldest; \
        force U_IF_NAME.io_diffCommits_info_363_pdest = RTL_PATH.io_diffCommits_info_363_pdest; \
        force U_IF_NAME.io_diffCommits_info_364_ldest = RTL_PATH.io_diffCommits_info_364_ldest; \
        force U_IF_NAME.io_diffCommits_info_364_pdest = RTL_PATH.io_diffCommits_info_364_pdest; \
        force U_IF_NAME.io_diffCommits_info_365_ldest = RTL_PATH.io_diffCommits_info_365_ldest; \
        force U_IF_NAME.io_diffCommits_info_365_pdest = RTL_PATH.io_diffCommits_info_365_pdest; \
        force U_IF_NAME.io_diffCommits_info_366_ldest = RTL_PATH.io_diffCommits_info_366_ldest; \
        force U_IF_NAME.io_diffCommits_info_366_pdest = RTL_PATH.io_diffCommits_info_366_pdest; \
        force U_IF_NAME.io_diffCommits_info_367_ldest = RTL_PATH.io_diffCommits_info_367_ldest; \
        force U_IF_NAME.io_diffCommits_info_367_pdest = RTL_PATH.io_diffCommits_info_367_pdest; \
        force U_IF_NAME.io_diffCommits_info_368_ldest = RTL_PATH.io_diffCommits_info_368_ldest; \
        force U_IF_NAME.io_diffCommits_info_368_pdest = RTL_PATH.io_diffCommits_info_368_pdest; \
        force U_IF_NAME.io_diffCommits_info_369_ldest = RTL_PATH.io_diffCommits_info_369_ldest; \
        force U_IF_NAME.io_diffCommits_info_369_pdest = RTL_PATH.io_diffCommits_info_369_pdest; \
        force U_IF_NAME.io_diffCommits_info_370_ldest = RTL_PATH.io_diffCommits_info_370_ldest; \
        force U_IF_NAME.io_diffCommits_info_370_pdest = RTL_PATH.io_diffCommits_info_370_pdest; \
        force U_IF_NAME.io_diffCommits_info_371_ldest = RTL_PATH.io_diffCommits_info_371_ldest; \
        force U_IF_NAME.io_diffCommits_info_371_pdest = RTL_PATH.io_diffCommits_info_371_pdest; \
        force U_IF_NAME.io_diffCommits_info_372_ldest = RTL_PATH.io_diffCommits_info_372_ldest; \
        force U_IF_NAME.io_diffCommits_info_372_pdest = RTL_PATH.io_diffCommits_info_372_pdest; \
        force U_IF_NAME.io_diffCommits_info_373_ldest = RTL_PATH.io_diffCommits_info_373_ldest; \
        force U_IF_NAME.io_diffCommits_info_373_pdest = RTL_PATH.io_diffCommits_info_373_pdest; \
        force U_IF_NAME.io_diffCommits_info_374_ldest = RTL_PATH.io_diffCommits_info_374_ldest; \
        force U_IF_NAME.io_diffCommits_info_374_pdest = RTL_PATH.io_diffCommits_info_374_pdest; \
        force U_IF_NAME.io_diffCommits_info_375_ldest = RTL_PATH.io_diffCommits_info_375_ldest; \
        force U_IF_NAME.io_diffCommits_info_375_pdest = RTL_PATH.io_diffCommits_info_375_pdest; \
        force U_IF_NAME.io_diffCommits_info_376_ldest = RTL_PATH.io_diffCommits_info_376_ldest; \
        force U_IF_NAME.io_diffCommits_info_376_pdest = RTL_PATH.io_diffCommits_info_376_pdest; \
        force U_IF_NAME.io_diffCommits_info_377_ldest = RTL_PATH.io_diffCommits_info_377_ldest; \
        force U_IF_NAME.io_diffCommits_info_377_pdest = RTL_PATH.io_diffCommits_info_377_pdest; \
        force U_IF_NAME.io_diffCommits_info_378_ldest = RTL_PATH.io_diffCommits_info_378_ldest; \
        force U_IF_NAME.io_diffCommits_info_378_pdest = RTL_PATH.io_diffCommits_info_378_pdest; \
        force U_IF_NAME.io_diffCommits_info_379_ldest = RTL_PATH.io_diffCommits_info_379_ldest; \
        force U_IF_NAME.io_diffCommits_info_379_pdest = RTL_PATH.io_diffCommits_info_379_pdest; \
        force U_IF_NAME.io_diffCommits_info_380_ldest = RTL_PATH.io_diffCommits_info_380_ldest; \
        force U_IF_NAME.io_diffCommits_info_380_pdest = RTL_PATH.io_diffCommits_info_380_pdest; \
        force U_IF_NAME.io_diffCommits_info_381_ldest = RTL_PATH.io_diffCommits_info_381_ldest; \
        force U_IF_NAME.io_diffCommits_info_381_pdest = RTL_PATH.io_diffCommits_info_381_pdest; \
        force U_IF_NAME.io_diffCommits_info_382_ldest = RTL_PATH.io_diffCommits_info_382_ldest; \
        force U_IF_NAME.io_diffCommits_info_382_pdest = RTL_PATH.io_diffCommits_info_382_pdest; \
        force U_IF_NAME.io_diffCommits_info_383_ldest = RTL_PATH.io_diffCommits_info_383_ldest; \
        force U_IF_NAME.io_diffCommits_info_383_pdest = RTL_PATH.io_diffCommits_info_383_pdest; \
        force U_IF_NAME.io_diffCommits_info_384_ldest = RTL_PATH.io_diffCommits_info_384_ldest; \
        force U_IF_NAME.io_diffCommits_info_384_pdest = RTL_PATH.io_diffCommits_info_384_pdest; \
        force U_IF_NAME.io_diffCommits_info_385_ldest = RTL_PATH.io_diffCommits_info_385_ldest; \
        force U_IF_NAME.io_diffCommits_info_385_pdest = RTL_PATH.io_diffCommits_info_385_pdest; \
        force U_IF_NAME.io_diffCommits_info_386_ldest = RTL_PATH.io_diffCommits_info_386_ldest; \
        force U_IF_NAME.io_diffCommits_info_386_pdest = RTL_PATH.io_diffCommits_info_386_pdest; \
        force U_IF_NAME.io_diffCommits_info_387_ldest = RTL_PATH.io_diffCommits_info_387_ldest; \
        force U_IF_NAME.io_diffCommits_info_387_pdest = RTL_PATH.io_diffCommits_info_387_pdest; \
        force U_IF_NAME.io_diffCommits_info_388_ldest = RTL_PATH.io_diffCommits_info_388_ldest; \
        force U_IF_NAME.io_diffCommits_info_388_pdest = RTL_PATH.io_diffCommits_info_388_pdest; \
        force U_IF_NAME.io_diffCommits_info_389_ldest = RTL_PATH.io_diffCommits_info_389_ldest; \
        force U_IF_NAME.io_diffCommits_info_389_pdest = RTL_PATH.io_diffCommits_info_389_pdest; \
        force U_IF_NAME.io_lsq_scommit = RTL_PATH.io_lsq_scommit; \
        force U_IF_NAME.io_lsq_pendingMMIOld = RTL_PATH.io_lsq_pendingMMIOld; \
        force U_IF_NAME.io_lsq_pendingst = RTL_PATH.io_lsq_pendingst; \
        force U_IF_NAME.io_lsq_pendingPtr_flag = RTL_PATH.io_lsq_pendingPtr_flag; \
        force U_IF_NAME.io_lsq_pendingPtr_value = RTL_PATH.io_lsq_pendingPtr_value; \
        force U_IF_NAME.io_robDeqPtr_flag = RTL_PATH.io_robDeqPtr_flag; \
        force U_IF_NAME.io_robDeqPtr_value = RTL_PATH.io_robDeqPtr_value; \
        force U_IF_NAME.io_csr_fflags_valid = RTL_PATH.io_csr_fflags_valid; \
        force U_IF_NAME.io_csr_fflags_bits = RTL_PATH.io_csr_fflags_bits; \
        force U_IF_NAME.io_csr_vxsat_valid = RTL_PATH.io_csr_vxsat_valid; \
        force U_IF_NAME.io_csr_vxsat_bits = RTL_PATH.io_csr_vxsat_bits; \
        force U_IF_NAME.io_csr_vstart_valid = RTL_PATH.io_csr_vstart_valid; \
        force U_IF_NAME.io_csr_vstart_bits = RTL_PATH.io_csr_vstart_bits; \
        force U_IF_NAME.io_csr_dirty_fs = RTL_PATH.io_csr_dirty_fs; \
        force U_IF_NAME.io_csr_dirty_vs = RTL_PATH.io_csr_dirty_vs; \
        force U_IF_NAME.io_csr_perfinfo_retiredInstr = RTL_PATH.io_csr_perfinfo_retiredInstr; \
        force U_IF_NAME.io_cpu_halt = RTL_PATH.io_cpu_halt; \
        force U_IF_NAME.io_wfi_wfiReq = RTL_PATH.io_wfi_wfiReq; \
        force U_IF_NAME.io_toDecode_isResumeVType = RTL_PATH.io_toDecode_isResumeVType; \
        force U_IF_NAME.io_toDecode_walkToArchVType = RTL_PATH.io_toDecode_walkToArchVType; \
        force U_IF_NAME.io_toDecode_walkVType_valid = RTL_PATH.io_toDecode_walkVType_valid; \
        force U_IF_NAME.io_toDecode_walkVType_bits_illegal = RTL_PATH.io_toDecode_walkVType_bits_illegal; \
        force U_IF_NAME.io_toDecode_walkVType_bits_vma = RTL_PATH.io_toDecode_walkVType_bits_vma; \
        force U_IF_NAME.io_toDecode_walkVType_bits_vta = RTL_PATH.io_toDecode_walkVType_bits_vta; \
        force U_IF_NAME.io_toDecode_walkVType_bits_vsew = RTL_PATH.io_toDecode_walkVType_bits_vsew; \
        force U_IF_NAME.io_toDecode_walkVType_bits_vlmul = RTL_PATH.io_toDecode_walkVType_bits_vlmul; \
        force U_IF_NAME.io_toDecode_commitVType_vtype_valid = RTL_PATH.io_toDecode_commitVType_vtype_valid; \
        force U_IF_NAME.io_toDecode_commitVType_vtype_bits_illegal = RTL_PATH.io_toDecode_commitVType_vtype_bits_illegal; \
        force U_IF_NAME.io_toDecode_commitVType_vtype_bits_vma = RTL_PATH.io_toDecode_commitVType_vtype_bits_vma; \
        force U_IF_NAME.io_toDecode_commitVType_vtype_bits_vta = RTL_PATH.io_toDecode_commitVType_vtype_bits_vta; \
        force U_IF_NAME.io_toDecode_commitVType_vtype_bits_vsew = RTL_PATH.io_toDecode_commitVType_vtype_bits_vsew; \
        force U_IF_NAME.io_toDecode_commitVType_vtype_bits_vlmul = RTL_PATH.io_toDecode_commitVType_vtype_bits_vlmul; \
        force U_IF_NAME.io_toDecode_commitVType_hasVsetvl = RTL_PATH.io_toDecode_commitVType_hasVsetvl; \
        force U_IF_NAME.io_readGPAMemAddr_valid = RTL_PATH.io_readGPAMemAddr_valid; \
        force U_IF_NAME.io_readGPAMemAddr_bits_ftqPtr_value = RTL_PATH.io_readGPAMemAddr_bits_ftqPtr_value; \
        force U_IF_NAME.io_readGPAMemAddr_bits_ftqOffset = RTL_PATH.io_readGPAMemAddr_bits_ftqOffset; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_0_valid = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_0_valid; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_0_bits_lreg = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_0_bits_lreg; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_0_bits_preg = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_0_bits_preg; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_1_valid = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_1_valid; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_1_bits_lreg = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_1_bits_lreg; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_1_bits_preg = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_1_bits_preg; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_2_valid = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_2_valid; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_2_bits_lreg = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_2_bits_lreg; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_2_bits_preg = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_2_bits_preg; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_3_valid = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_3_valid; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_3_bits_lreg = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_3_bits_lreg; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_3_bits_preg = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_3_bits_preg; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_4_valid = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_4_valid; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_4_bits_lreg = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_4_bits_lreg; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_4_bits_preg = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_4_bits_preg; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_5_valid = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_5_valid; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_5_bits_lreg = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_5_bits_lreg; \
        force U_IF_NAME.io_toVecExcpMod_logicPhyRegMap_5_bits_preg = RTL_PATH.io_toVecExcpMod_logicPhyRegMap_5_bits_preg; \
        force U_IF_NAME.io_toVecExcpMod_excpInfo_valid = RTL_PATH.io_toVecExcpMod_excpInfo_valid; \
        force U_IF_NAME.io_toVecExcpMod_excpInfo_bits_vstart = RTL_PATH.io_toVecExcpMod_excpInfo_bits_vstart; \
        force U_IF_NAME.io_toVecExcpMod_excpInfo_bits_vsew = RTL_PATH.io_toVecExcpMod_excpInfo_bits_vsew; \
        force U_IF_NAME.io_toVecExcpMod_excpInfo_bits_veew = RTL_PATH.io_toVecExcpMod_excpInfo_bits_veew; \
        force U_IF_NAME.io_toVecExcpMod_excpInfo_bits_vlmul = RTL_PATH.io_toVecExcpMod_excpInfo_bits_vlmul; \
        force U_IF_NAME.io_toVecExcpMod_excpInfo_bits_nf = RTL_PATH.io_toVecExcpMod_excpInfo_bits_nf; \
        force U_IF_NAME.io_toVecExcpMod_excpInfo_bits_isStride = RTL_PATH.io_toVecExcpMod_excpInfo_bits_isStride; \
        force U_IF_NAME.io_toVecExcpMod_excpInfo_bits_isIndexed = RTL_PATH.io_toVecExcpMod_excpInfo_bits_isIndexed; \
        force U_IF_NAME.io_toVecExcpMod_excpInfo_bits_isWhole = RTL_PATH.io_toVecExcpMod_excpInfo_bits_isWhole; \
        force U_IF_NAME.io_toVecExcpMod_excpInfo_bits_isVlm = RTL_PATH.io_toVecExcpMod_excpInfo_bits_isVlm; \
        force U_IF_NAME.io_storeDebugInfo_1_pc = RTL_PATH.io_storeDebugInfo_1_pc; \
        force U_IF_NAME.io_perf_0_value = RTL_PATH.io_perf_0_value; \
        force U_IF_NAME.io_perf_1_value = RTL_PATH.io_perf_1_value; \
        force U_IF_NAME.io_perf_2_value = RTL_PATH.io_perf_2_value; \
        force U_IF_NAME.io_perf_3_value = RTL_PATH.io_perf_3_value; \
        force U_IF_NAME.io_perf_4_value = RTL_PATH.io_perf_4_value; \
        force U_IF_NAME.io_perf_5_value = RTL_PATH.io_perf_5_value; \
        force U_IF_NAME.io_perf_6_value = RTL_PATH.io_perf_6_value; \
        force U_IF_NAME.io_perf_7_value = RTL_PATH.io_perf_7_value; \
        force U_IF_NAME.io_perf_8_value = RTL_PATH.io_perf_8_value; \
        force U_IF_NAME.io_perf_9_value = RTL_PATH.io_perf_9_value; \
        force U_IF_NAME.io_perf_10_value = RTL_PATH.io_perf_10_value; \
        force U_IF_NAME.io_perf_11_value = RTL_PATH.io_perf_11_value; \
        force U_IF_NAME.io_perf_12_value = RTL_PATH.io_perf_12_value; \
        force U_IF_NAME.io_perf_13_value = RTL_PATH.io_perf_13_value; \
        force U_IF_NAME.io_perf_14_value = RTL_PATH.io_perf_14_value; \
        force U_IF_NAME.io_perf_15_value = RTL_PATH.io_perf_15_value; \
        force U_IF_NAME.io_perf_16_value = RTL_PATH.io_perf_16_value; \
        force U_IF_NAME.io_perf_17_value = RTL_PATH.io_perf_17_value; \
        force U_IF_NAME.io_error_0 = RTL_PATH.io_error_0; \
    end \
    `endif

`endif

//=========================================================
//File name    : rename_in_agent_driver.sv
//Author       : nanyunhao
//Module name  : rename_in_agent_driver
//Discribution : rename_in_agent_driver : driver
//Date         : 2026-01-22
//=========================================================
`ifndef RENAME_IN_AGENT_DRIVER__SV
`define RENAME_IN_AGENT_DRIVER__SV

class rename_in_agent_driver  extends tcnt_driver_base#(virtual rename_in_agent_interface,rename_in_agent_cfg,rename_in_agent_xaction);

    `uvm_component_utils(rename_in_agent_driver)

    extern function new(string name, uvm_component parent);
    extern virtual function void build_phase(uvm_phase phase);
    extern virtual task reset_phase(uvm_phase phase);
    extern task main_phase(uvm_phase phase);
    extern task send_pkt(rename_in_agent_xaction tr);
    extern task drive_idle(tcnt_dec_base::drv_mode_e drv_mode);
endclass:rename_in_agent_driver

function rename_in_agent_driver::new(string name, uvm_component parent);
    super.new(name,parent);
endfunction:new

function void rename_in_agent_driver::build_phase(uvm_phase phase);
    super.build_phase(phase);
endfunction:build_phase

task rename_in_agent_driver::reset_phase(uvm_phase phase);

    super.reset_phase(phase);
    phase.raise_objection(this);

    repeat(2) begin
        @this.vif.drv_mp.drv_cb;
        this.drive_idle(this.cfg.drv_mode);
    end
    wait(vif.rst_n == 1'b1);
    repeat(20) begin
        @this.vif.drv_mp.drv_cb;
        this.drive_idle(this.cfg.drv_mode);
    end

    phase.drop_objection(this);
endtask:reset_phase

task rename_in_agent_driver::main_phase(uvm_phase phase);
    super.main_phase(phase);
    //while(1) begin
    if(this.cfg.sqr_sw==tcnt_dec_base::ON && this.cfg.drv_sw==tcnt_dec_base::ON) begin
        while(1) begin
            seq_item_port.try_next_item(req);
            if(req!=null) begin
                repeat(req.pre_pkt_gap) begin
                    @this.vif.drv_mp.drv_cb;
                    this.drive_idle(this.cfg.drv_mode);
                end
                @this.vif.drv_mp.drv_cb;
                this.send_pkt(req);
                repeat(req.post_pkt_gap) begin
                    @this.vif.drv_mp.drv_cb;
                    this.drive_idle(this.cfg.drv_mode);
                end
                seq_item_port.item_done();
            end
            else begin
                @this.vif.drv_mp.drv_cb;
                this.drive_idle(this.cfg.drv_mode);
            end
        end
    end
    else if (this.cfg.drv_sw==tcnt_dec_base::ON) begin
        while(1) begin
            @this.vif.drv_mp.drv_cb;
            `uvm_fatal(get_type_name(), $sformatf("sqr_sw==OFF & drv_sw==ON, please give a driver send task!"))
            //send task
        end
    end
endtask:main_phase

task rename_in_agent_driver::send_pkt(rename_in_agent_xaction tr);
    vif.drv_mp.drv_cb.clock <= tr.clock; 
    vif.drv_mp.drv_cb.reset <= tr.reset; 
    vif.drv_mp.drv_cb.io_hartId <= tr.io_hartId; 
    vif.drv_mp.drv_cb.io_enq_req_0_valid <= tr.io_enq_req_0_valid; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_instr <= tr.io_enq_req_0_bits_instr; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_pc <= tr.io_enq_req_0_bits_pc; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_0 <= tr.io_enq_req_0_bits_exceptionVec_0; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_1 <= tr.io_enq_req_0_bits_exceptionVec_1; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_2 <= tr.io_enq_req_0_bits_exceptionVec_2; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_3 <= tr.io_enq_req_0_bits_exceptionVec_3; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_12 <= tr.io_enq_req_0_bits_exceptionVec_12; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_20 <= tr.io_enq_req_0_bits_exceptionVec_20; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_22 <= tr.io_enq_req_0_bits_exceptionVec_22; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_isFetchMalAddr <= tr.io_enq_req_0_bits_isFetchMalAddr; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_hasException <= tr.io_enq_req_0_bits_hasException; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_trigger <= tr.io_enq_req_0_bits_trigger; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_preDecodeInfo_isRVC <= tr.io_enq_req_0_bits_preDecodeInfo_isRVC; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_crossPageIPFFix <= tr.io_enq_req_0_bits_crossPageIPFFix; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_ftqPtr_flag <= tr.io_enq_req_0_bits_ftqPtr_flag; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_ftqPtr_value <= tr.io_enq_req_0_bits_ftqPtr_value; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_ftqOffset <= tr.io_enq_req_0_bits_ftqOffset; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_ldest <= tr.io_enq_req_0_bits_ldest; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_fuType <= tr.io_enq_req_0_bits_fuType; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_fuOpType <= tr.io_enq_req_0_bits_fuOpType; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_rfWen <= tr.io_enq_req_0_bits_rfWen; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_fpWen <= tr.io_enq_req_0_bits_fpWen; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_vecWen <= tr.io_enq_req_0_bits_vecWen; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_v0Wen <= tr.io_enq_req_0_bits_v0Wen; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_vlWen <= tr.io_enq_req_0_bits_vlWen; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_isXSTrap <= tr.io_enq_req_0_bits_isXSTrap; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_waitForward <= tr.io_enq_req_0_bits_waitForward; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_blockBackward <= tr.io_enq_req_0_bits_blockBackward; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_flushPipe <= tr.io_enq_req_0_bits_flushPipe; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vill <= tr.io_enq_req_0_bits_vpu_vill; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vma <= tr.io_enq_req_0_bits_vpu_vma; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vta <= tr.io_enq_req_0_bits_vpu_vta; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vsew <= tr.io_enq_req_0_bits_vpu_vsew; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vlmul <= tr.io_enq_req_0_bits_vpu_vlmul; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVill <= tr.io_enq_req_0_bits_vpu_specVill; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVma <= tr.io_enq_req_0_bits_vpu_specVma; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVta <= tr.io_enq_req_0_bits_vpu_specVta; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVsew <= tr.io_enq_req_0_bits_vpu_specVsew; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVlmul <= tr.io_enq_req_0_bits_vpu_specVlmul; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_vlsInstr <= tr.io_enq_req_0_bits_vlsInstr; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_wfflags <= tr.io_enq_req_0_bits_wfflags; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_isMove <= tr.io_enq_req_0_bits_isMove; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_isVset <= tr.io_enq_req_0_bits_isVset; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_firstUop <= tr.io_enq_req_0_bits_firstUop; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_lastUop <= tr.io_enq_req_0_bits_lastUop; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_numWB <= tr.io_enq_req_0_bits_numWB; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_commitType <= tr.io_enq_req_0_bits_commitType; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_pdest <= tr.io_enq_req_0_bits_pdest; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_robIdx_flag <= tr.io_enq_req_0_bits_robIdx_flag; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_robIdx_value <= tr.io_enq_req_0_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_instrSize <= tr.io_enq_req_0_bits_instrSize; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_dirtyFs <= tr.io_enq_req_0_bits_dirtyFs; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_dirtyVs <= tr.io_enq_req_0_bits_dirtyVs; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_traceBlockInPipe_itype <= tr.io_enq_req_0_bits_traceBlockInPipe_itype; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_traceBlockInPipe_iretire <= tr.io_enq_req_0_bits_traceBlockInPipe_iretire; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_traceBlockInPipe_ilastsize <= tr.io_enq_req_0_bits_traceBlockInPipe_ilastsize; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_eliminatedMove <= tr.io_enq_req_0_bits_eliminatedMove; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_snapshot <= tr.io_enq_req_0_bits_snapshot; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_lqIdx_value <= tr.io_enq_req_0_bits_lqIdx_value; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_sqIdx_value <= tr.io_enq_req_0_bits_sqIdx_value; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_singleStep <= tr.io_enq_req_0_bits_singleStep; 
    vif.drv_mp.drv_cb.io_enq_req_0_bits_debug_sim_trig <= tr.io_enq_req_0_bits_debug_sim_trig; 
    vif.drv_mp.drv_cb.io_enq_req_1_valid <= tr.io_enq_req_1_valid; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_instr <= tr.io_enq_req_1_bits_instr; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_pc <= tr.io_enq_req_1_bits_pc; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_0 <= tr.io_enq_req_1_bits_exceptionVec_0; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_1 <= tr.io_enq_req_1_bits_exceptionVec_1; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_2 <= tr.io_enq_req_1_bits_exceptionVec_2; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_3 <= tr.io_enq_req_1_bits_exceptionVec_3; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_12 <= tr.io_enq_req_1_bits_exceptionVec_12; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_20 <= tr.io_enq_req_1_bits_exceptionVec_20; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_22 <= tr.io_enq_req_1_bits_exceptionVec_22; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_isFetchMalAddr <= tr.io_enq_req_1_bits_isFetchMalAddr; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_hasException <= tr.io_enq_req_1_bits_hasException; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_trigger <= tr.io_enq_req_1_bits_trigger; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_preDecodeInfo_isRVC <= tr.io_enq_req_1_bits_preDecodeInfo_isRVC; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_crossPageIPFFix <= tr.io_enq_req_1_bits_crossPageIPFFix; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_ftqPtr_flag <= tr.io_enq_req_1_bits_ftqPtr_flag; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_ftqPtr_value <= tr.io_enq_req_1_bits_ftqPtr_value; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_ftqOffset <= tr.io_enq_req_1_bits_ftqOffset; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_ldest <= tr.io_enq_req_1_bits_ldest; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_fuType <= tr.io_enq_req_1_bits_fuType; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_fuOpType <= tr.io_enq_req_1_bits_fuOpType; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_rfWen <= tr.io_enq_req_1_bits_rfWen; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_fpWen <= tr.io_enq_req_1_bits_fpWen; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_vecWen <= tr.io_enq_req_1_bits_vecWen; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_v0Wen <= tr.io_enq_req_1_bits_v0Wen; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_vlWen <= tr.io_enq_req_1_bits_vlWen; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_isXSTrap <= tr.io_enq_req_1_bits_isXSTrap; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_waitForward <= tr.io_enq_req_1_bits_waitForward; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_blockBackward <= tr.io_enq_req_1_bits_blockBackward; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_flushPipe <= tr.io_enq_req_1_bits_flushPipe; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vill <= tr.io_enq_req_1_bits_vpu_vill; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vma <= tr.io_enq_req_1_bits_vpu_vma; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vta <= tr.io_enq_req_1_bits_vpu_vta; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vsew <= tr.io_enq_req_1_bits_vpu_vsew; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vlmul <= tr.io_enq_req_1_bits_vpu_vlmul; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVill <= tr.io_enq_req_1_bits_vpu_specVill; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVma <= tr.io_enq_req_1_bits_vpu_specVma; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVta <= tr.io_enq_req_1_bits_vpu_specVta; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVsew <= tr.io_enq_req_1_bits_vpu_specVsew; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVlmul <= tr.io_enq_req_1_bits_vpu_specVlmul; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_vlsInstr <= tr.io_enq_req_1_bits_vlsInstr; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_wfflags <= tr.io_enq_req_1_bits_wfflags; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_isMove <= tr.io_enq_req_1_bits_isMove; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_isVset <= tr.io_enq_req_1_bits_isVset; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_firstUop <= tr.io_enq_req_1_bits_firstUop; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_lastUop <= tr.io_enq_req_1_bits_lastUop; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_numWB <= tr.io_enq_req_1_bits_numWB; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_commitType <= tr.io_enq_req_1_bits_commitType; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_pdest <= tr.io_enq_req_1_bits_pdest; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_robIdx_flag <= tr.io_enq_req_1_bits_robIdx_flag; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_robIdx_value <= tr.io_enq_req_1_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_instrSize <= tr.io_enq_req_1_bits_instrSize; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_dirtyFs <= tr.io_enq_req_1_bits_dirtyFs; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_dirtyVs <= tr.io_enq_req_1_bits_dirtyVs; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_traceBlockInPipe_itype <= tr.io_enq_req_1_bits_traceBlockInPipe_itype; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_traceBlockInPipe_iretire <= tr.io_enq_req_1_bits_traceBlockInPipe_iretire; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_traceBlockInPipe_ilastsize <= tr.io_enq_req_1_bits_traceBlockInPipe_ilastsize; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_eliminatedMove <= tr.io_enq_req_1_bits_eliminatedMove; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_snapshot <= tr.io_enq_req_1_bits_snapshot; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_lqIdx_value <= tr.io_enq_req_1_bits_lqIdx_value; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_sqIdx_value <= tr.io_enq_req_1_bits_sqIdx_value; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_singleStep <= tr.io_enq_req_1_bits_singleStep; 
    vif.drv_mp.drv_cb.io_enq_req_1_bits_debug_sim_trig <= tr.io_enq_req_1_bits_debug_sim_trig; 
    vif.drv_mp.drv_cb.io_enq_req_2_valid <= tr.io_enq_req_2_valid; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_instr <= tr.io_enq_req_2_bits_instr; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_pc <= tr.io_enq_req_2_bits_pc; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_0 <= tr.io_enq_req_2_bits_exceptionVec_0; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_1 <= tr.io_enq_req_2_bits_exceptionVec_1; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_2 <= tr.io_enq_req_2_bits_exceptionVec_2; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_3 <= tr.io_enq_req_2_bits_exceptionVec_3; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_12 <= tr.io_enq_req_2_bits_exceptionVec_12; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_20 <= tr.io_enq_req_2_bits_exceptionVec_20; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_22 <= tr.io_enq_req_2_bits_exceptionVec_22; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_isFetchMalAddr <= tr.io_enq_req_2_bits_isFetchMalAddr; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_hasException <= tr.io_enq_req_2_bits_hasException; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_trigger <= tr.io_enq_req_2_bits_trigger; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_preDecodeInfo_isRVC <= tr.io_enq_req_2_bits_preDecodeInfo_isRVC; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_crossPageIPFFix <= tr.io_enq_req_2_bits_crossPageIPFFix; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_ftqPtr_flag <= tr.io_enq_req_2_bits_ftqPtr_flag; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_ftqPtr_value <= tr.io_enq_req_2_bits_ftqPtr_value; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_ftqOffset <= tr.io_enq_req_2_bits_ftqOffset; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_ldest <= tr.io_enq_req_2_bits_ldest; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_fuType <= tr.io_enq_req_2_bits_fuType; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_fuOpType <= tr.io_enq_req_2_bits_fuOpType; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_rfWen <= tr.io_enq_req_2_bits_rfWen; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_fpWen <= tr.io_enq_req_2_bits_fpWen; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_vecWen <= tr.io_enq_req_2_bits_vecWen; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_v0Wen <= tr.io_enq_req_2_bits_v0Wen; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_vlWen <= tr.io_enq_req_2_bits_vlWen; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_isXSTrap <= tr.io_enq_req_2_bits_isXSTrap; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_waitForward <= tr.io_enq_req_2_bits_waitForward; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_blockBackward <= tr.io_enq_req_2_bits_blockBackward; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_flushPipe <= tr.io_enq_req_2_bits_flushPipe; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vill <= tr.io_enq_req_2_bits_vpu_vill; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vma <= tr.io_enq_req_2_bits_vpu_vma; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vta <= tr.io_enq_req_2_bits_vpu_vta; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vsew <= tr.io_enq_req_2_bits_vpu_vsew; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vlmul <= tr.io_enq_req_2_bits_vpu_vlmul; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVill <= tr.io_enq_req_2_bits_vpu_specVill; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVma <= tr.io_enq_req_2_bits_vpu_specVma; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVta <= tr.io_enq_req_2_bits_vpu_specVta; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVsew <= tr.io_enq_req_2_bits_vpu_specVsew; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVlmul <= tr.io_enq_req_2_bits_vpu_specVlmul; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_vlsInstr <= tr.io_enq_req_2_bits_vlsInstr; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_wfflags <= tr.io_enq_req_2_bits_wfflags; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_isMove <= tr.io_enq_req_2_bits_isMove; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_isVset <= tr.io_enq_req_2_bits_isVset; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_firstUop <= tr.io_enq_req_2_bits_firstUop; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_lastUop <= tr.io_enq_req_2_bits_lastUop; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_numWB <= tr.io_enq_req_2_bits_numWB; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_commitType <= tr.io_enq_req_2_bits_commitType; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_pdest <= tr.io_enq_req_2_bits_pdest; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_robIdx_flag <= tr.io_enq_req_2_bits_robIdx_flag; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_robIdx_value <= tr.io_enq_req_2_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_instrSize <= tr.io_enq_req_2_bits_instrSize; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_dirtyFs <= tr.io_enq_req_2_bits_dirtyFs; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_dirtyVs <= tr.io_enq_req_2_bits_dirtyVs; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_traceBlockInPipe_itype <= tr.io_enq_req_2_bits_traceBlockInPipe_itype; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_traceBlockInPipe_iretire <= tr.io_enq_req_2_bits_traceBlockInPipe_iretire; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_traceBlockInPipe_ilastsize <= tr.io_enq_req_2_bits_traceBlockInPipe_ilastsize; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_eliminatedMove <= tr.io_enq_req_2_bits_eliminatedMove; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_snapshot <= tr.io_enq_req_2_bits_snapshot; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_lqIdx_value <= tr.io_enq_req_2_bits_lqIdx_value; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_sqIdx_value <= tr.io_enq_req_2_bits_sqIdx_value; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_singleStep <= tr.io_enq_req_2_bits_singleStep; 
    vif.drv_mp.drv_cb.io_enq_req_2_bits_debug_sim_trig <= tr.io_enq_req_2_bits_debug_sim_trig; 
    vif.drv_mp.drv_cb.io_enq_req_3_valid <= tr.io_enq_req_3_valid; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_instr <= tr.io_enq_req_3_bits_instr; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_pc <= tr.io_enq_req_3_bits_pc; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_0 <= tr.io_enq_req_3_bits_exceptionVec_0; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_1 <= tr.io_enq_req_3_bits_exceptionVec_1; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_2 <= tr.io_enq_req_3_bits_exceptionVec_2; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_3 <= tr.io_enq_req_3_bits_exceptionVec_3; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_12 <= tr.io_enq_req_3_bits_exceptionVec_12; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_20 <= tr.io_enq_req_3_bits_exceptionVec_20; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_22 <= tr.io_enq_req_3_bits_exceptionVec_22; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_isFetchMalAddr <= tr.io_enq_req_3_bits_isFetchMalAddr; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_hasException <= tr.io_enq_req_3_bits_hasException; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_trigger <= tr.io_enq_req_3_bits_trigger; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_preDecodeInfo_isRVC <= tr.io_enq_req_3_bits_preDecodeInfo_isRVC; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_crossPageIPFFix <= tr.io_enq_req_3_bits_crossPageIPFFix; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_ftqPtr_flag <= tr.io_enq_req_3_bits_ftqPtr_flag; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_ftqPtr_value <= tr.io_enq_req_3_bits_ftqPtr_value; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_ftqOffset <= tr.io_enq_req_3_bits_ftqOffset; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_ldest <= tr.io_enq_req_3_bits_ldest; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_fuType <= tr.io_enq_req_3_bits_fuType; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_fuOpType <= tr.io_enq_req_3_bits_fuOpType; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_rfWen <= tr.io_enq_req_3_bits_rfWen; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_fpWen <= tr.io_enq_req_3_bits_fpWen; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_vecWen <= tr.io_enq_req_3_bits_vecWen; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_v0Wen <= tr.io_enq_req_3_bits_v0Wen; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_vlWen <= tr.io_enq_req_3_bits_vlWen; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_isXSTrap <= tr.io_enq_req_3_bits_isXSTrap; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_waitForward <= tr.io_enq_req_3_bits_waitForward; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_blockBackward <= tr.io_enq_req_3_bits_blockBackward; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_flushPipe <= tr.io_enq_req_3_bits_flushPipe; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vill <= tr.io_enq_req_3_bits_vpu_vill; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vma <= tr.io_enq_req_3_bits_vpu_vma; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vta <= tr.io_enq_req_3_bits_vpu_vta; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vsew <= tr.io_enq_req_3_bits_vpu_vsew; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vlmul <= tr.io_enq_req_3_bits_vpu_vlmul; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVill <= tr.io_enq_req_3_bits_vpu_specVill; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVma <= tr.io_enq_req_3_bits_vpu_specVma; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVta <= tr.io_enq_req_3_bits_vpu_specVta; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVsew <= tr.io_enq_req_3_bits_vpu_specVsew; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVlmul <= tr.io_enq_req_3_bits_vpu_specVlmul; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_vlsInstr <= tr.io_enq_req_3_bits_vlsInstr; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_wfflags <= tr.io_enq_req_3_bits_wfflags; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_isMove <= tr.io_enq_req_3_bits_isMove; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_isVset <= tr.io_enq_req_3_bits_isVset; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_firstUop <= tr.io_enq_req_3_bits_firstUop; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_lastUop <= tr.io_enq_req_3_bits_lastUop; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_numWB <= tr.io_enq_req_3_bits_numWB; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_commitType <= tr.io_enq_req_3_bits_commitType; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_pdest <= tr.io_enq_req_3_bits_pdest; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_robIdx_flag <= tr.io_enq_req_3_bits_robIdx_flag; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_robIdx_value <= tr.io_enq_req_3_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_instrSize <= tr.io_enq_req_3_bits_instrSize; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_dirtyFs <= tr.io_enq_req_3_bits_dirtyFs; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_dirtyVs <= tr.io_enq_req_3_bits_dirtyVs; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_traceBlockInPipe_itype <= tr.io_enq_req_3_bits_traceBlockInPipe_itype; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_traceBlockInPipe_iretire <= tr.io_enq_req_3_bits_traceBlockInPipe_iretire; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_traceBlockInPipe_ilastsize <= tr.io_enq_req_3_bits_traceBlockInPipe_ilastsize; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_eliminatedMove <= tr.io_enq_req_3_bits_eliminatedMove; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_snapshot <= tr.io_enq_req_3_bits_snapshot; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_lqIdx_value <= tr.io_enq_req_3_bits_lqIdx_value; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_sqIdx_value <= tr.io_enq_req_3_bits_sqIdx_value; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_singleStep <= tr.io_enq_req_3_bits_singleStep; 
    vif.drv_mp.drv_cb.io_enq_req_3_bits_debug_sim_trig <= tr.io_enq_req_3_bits_debug_sim_trig; 
    vif.drv_mp.drv_cb.io_enq_req_4_valid <= tr.io_enq_req_4_valid; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_instr <= tr.io_enq_req_4_bits_instr; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_pc <= tr.io_enq_req_4_bits_pc; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_0 <= tr.io_enq_req_4_bits_exceptionVec_0; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_1 <= tr.io_enq_req_4_bits_exceptionVec_1; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_2 <= tr.io_enq_req_4_bits_exceptionVec_2; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_3 <= tr.io_enq_req_4_bits_exceptionVec_3; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_12 <= tr.io_enq_req_4_bits_exceptionVec_12; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_20 <= tr.io_enq_req_4_bits_exceptionVec_20; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_22 <= tr.io_enq_req_4_bits_exceptionVec_22; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_isFetchMalAddr <= tr.io_enq_req_4_bits_isFetchMalAddr; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_hasException <= tr.io_enq_req_4_bits_hasException; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_trigger <= tr.io_enq_req_4_bits_trigger; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_preDecodeInfo_isRVC <= tr.io_enq_req_4_bits_preDecodeInfo_isRVC; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_crossPageIPFFix <= tr.io_enq_req_4_bits_crossPageIPFFix; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_ftqPtr_flag <= tr.io_enq_req_4_bits_ftqPtr_flag; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_ftqPtr_value <= tr.io_enq_req_4_bits_ftqPtr_value; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_ftqOffset <= tr.io_enq_req_4_bits_ftqOffset; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_ldest <= tr.io_enq_req_4_bits_ldest; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_fuType <= tr.io_enq_req_4_bits_fuType; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_fuOpType <= tr.io_enq_req_4_bits_fuOpType; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_rfWen <= tr.io_enq_req_4_bits_rfWen; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_fpWen <= tr.io_enq_req_4_bits_fpWen; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_vecWen <= tr.io_enq_req_4_bits_vecWen; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_v0Wen <= tr.io_enq_req_4_bits_v0Wen; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_vlWen <= tr.io_enq_req_4_bits_vlWen; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_isXSTrap <= tr.io_enq_req_4_bits_isXSTrap; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_waitForward <= tr.io_enq_req_4_bits_waitForward; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_blockBackward <= tr.io_enq_req_4_bits_blockBackward; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_flushPipe <= tr.io_enq_req_4_bits_flushPipe; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vill <= tr.io_enq_req_4_bits_vpu_vill; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vma <= tr.io_enq_req_4_bits_vpu_vma; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vta <= tr.io_enq_req_4_bits_vpu_vta; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vsew <= tr.io_enq_req_4_bits_vpu_vsew; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vlmul <= tr.io_enq_req_4_bits_vpu_vlmul; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVill <= tr.io_enq_req_4_bits_vpu_specVill; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVma <= tr.io_enq_req_4_bits_vpu_specVma; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVta <= tr.io_enq_req_4_bits_vpu_specVta; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVsew <= tr.io_enq_req_4_bits_vpu_specVsew; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVlmul <= tr.io_enq_req_4_bits_vpu_specVlmul; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_vlsInstr <= tr.io_enq_req_4_bits_vlsInstr; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_wfflags <= tr.io_enq_req_4_bits_wfflags; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_isMove <= tr.io_enq_req_4_bits_isMove; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_isVset <= tr.io_enq_req_4_bits_isVset; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_firstUop <= tr.io_enq_req_4_bits_firstUop; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_lastUop <= tr.io_enq_req_4_bits_lastUop; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_numWB <= tr.io_enq_req_4_bits_numWB; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_commitType <= tr.io_enq_req_4_bits_commitType; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_pdest <= tr.io_enq_req_4_bits_pdest; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_robIdx_flag <= tr.io_enq_req_4_bits_robIdx_flag; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_robIdx_value <= tr.io_enq_req_4_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_instrSize <= tr.io_enq_req_4_bits_instrSize; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_dirtyFs <= tr.io_enq_req_4_bits_dirtyFs; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_dirtyVs <= tr.io_enq_req_4_bits_dirtyVs; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_traceBlockInPipe_itype <= tr.io_enq_req_4_bits_traceBlockInPipe_itype; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_traceBlockInPipe_iretire <= tr.io_enq_req_4_bits_traceBlockInPipe_iretire; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_traceBlockInPipe_ilastsize <= tr.io_enq_req_4_bits_traceBlockInPipe_ilastsize; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_eliminatedMove <= tr.io_enq_req_4_bits_eliminatedMove; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_snapshot <= tr.io_enq_req_4_bits_snapshot; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_lqIdx_value <= tr.io_enq_req_4_bits_lqIdx_value; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_sqIdx_value <= tr.io_enq_req_4_bits_sqIdx_value; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_singleStep <= tr.io_enq_req_4_bits_singleStep; 
    vif.drv_mp.drv_cb.io_enq_req_4_bits_debug_sim_trig <= tr.io_enq_req_4_bits_debug_sim_trig; 
    vif.drv_mp.drv_cb.io_enq_req_5_valid <= tr.io_enq_req_5_valid; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_instr <= tr.io_enq_req_5_bits_instr; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_pc <= tr.io_enq_req_5_bits_pc; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_0 <= tr.io_enq_req_5_bits_exceptionVec_0; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_1 <= tr.io_enq_req_5_bits_exceptionVec_1; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_2 <= tr.io_enq_req_5_bits_exceptionVec_2; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_3 <= tr.io_enq_req_5_bits_exceptionVec_3; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_12 <= tr.io_enq_req_5_bits_exceptionVec_12; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_20 <= tr.io_enq_req_5_bits_exceptionVec_20; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_22 <= tr.io_enq_req_5_bits_exceptionVec_22; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_isFetchMalAddr <= tr.io_enq_req_5_bits_isFetchMalAddr; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_hasException <= tr.io_enq_req_5_bits_hasException; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_trigger <= tr.io_enq_req_5_bits_trigger; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_preDecodeInfo_isRVC <= tr.io_enq_req_5_bits_preDecodeInfo_isRVC; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_crossPageIPFFix <= tr.io_enq_req_5_bits_crossPageIPFFix; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_ftqPtr_flag <= tr.io_enq_req_5_bits_ftqPtr_flag; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_ftqPtr_value <= tr.io_enq_req_5_bits_ftqPtr_value; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_ftqOffset <= tr.io_enq_req_5_bits_ftqOffset; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_ldest <= tr.io_enq_req_5_bits_ldest; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_fuType <= tr.io_enq_req_5_bits_fuType; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_fuOpType <= tr.io_enq_req_5_bits_fuOpType; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_rfWen <= tr.io_enq_req_5_bits_rfWen; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_fpWen <= tr.io_enq_req_5_bits_fpWen; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_vecWen <= tr.io_enq_req_5_bits_vecWen; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_v0Wen <= tr.io_enq_req_5_bits_v0Wen; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_vlWen <= tr.io_enq_req_5_bits_vlWen; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_isXSTrap <= tr.io_enq_req_5_bits_isXSTrap; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_waitForward <= tr.io_enq_req_5_bits_waitForward; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_blockBackward <= tr.io_enq_req_5_bits_blockBackward; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_flushPipe <= tr.io_enq_req_5_bits_flushPipe; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vill <= tr.io_enq_req_5_bits_vpu_vill; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vma <= tr.io_enq_req_5_bits_vpu_vma; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vta <= tr.io_enq_req_5_bits_vpu_vta; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vsew <= tr.io_enq_req_5_bits_vpu_vsew; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vlmul <= tr.io_enq_req_5_bits_vpu_vlmul; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVill <= tr.io_enq_req_5_bits_vpu_specVill; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVma <= tr.io_enq_req_5_bits_vpu_specVma; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVta <= tr.io_enq_req_5_bits_vpu_specVta; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVsew <= tr.io_enq_req_5_bits_vpu_specVsew; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVlmul <= tr.io_enq_req_5_bits_vpu_specVlmul; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_vlsInstr <= tr.io_enq_req_5_bits_vlsInstr; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_wfflags <= tr.io_enq_req_5_bits_wfflags; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_isMove <= tr.io_enq_req_5_bits_isMove; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_isVset <= tr.io_enq_req_5_bits_isVset; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_firstUop <= tr.io_enq_req_5_bits_firstUop; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_lastUop <= tr.io_enq_req_5_bits_lastUop; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_numWB <= tr.io_enq_req_5_bits_numWB; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_commitType <= tr.io_enq_req_5_bits_commitType; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_pdest <= tr.io_enq_req_5_bits_pdest; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_robIdx_flag <= tr.io_enq_req_5_bits_robIdx_flag; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_robIdx_value <= tr.io_enq_req_5_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_instrSize <= tr.io_enq_req_5_bits_instrSize; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_dirtyFs <= tr.io_enq_req_5_bits_dirtyFs; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_dirtyVs <= tr.io_enq_req_5_bits_dirtyVs; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_traceBlockInPipe_itype <= tr.io_enq_req_5_bits_traceBlockInPipe_itype; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_traceBlockInPipe_iretire <= tr.io_enq_req_5_bits_traceBlockInPipe_iretire; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_traceBlockInPipe_ilastsize <= tr.io_enq_req_5_bits_traceBlockInPipe_ilastsize; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_eliminatedMove <= tr.io_enq_req_5_bits_eliminatedMove; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_snapshot <= tr.io_enq_req_5_bits_snapshot; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_lqIdx_value <= tr.io_enq_req_5_bits_lqIdx_value; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_sqIdx_value <= tr.io_enq_req_5_bits_sqIdx_value; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_singleStep <= tr.io_enq_req_5_bits_singleStep; 
    vif.drv_mp.drv_cb.io_enq_req_5_bits_debug_sim_trig <= tr.io_enq_req_5_bits_debug_sim_trig; 

endtask:send_pkt

task rename_in_agent_driver::drive_idle(tcnt_dec_base::drv_mode_e drv_mode);

    if(drv_mode==tcnt_dec_base::DRV_0) begin
        vif.drv_mp.drv_cb.clock <= '0;
        vif.drv_mp.drv_cb.reset <= '0;
        vif.drv_mp.drv_cb.io_hartId <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_valid <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_instr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_pc <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_0 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_1 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_3 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_12 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_20 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_22 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_isFetchMalAddr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_hasException <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_trigger <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_preDecodeInfo_isRVC <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_crossPageIPFFix <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_ftqPtr_flag <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_ftqPtr_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_ftqOffset <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_ldest <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_fuType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_fuOpType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_rfWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_fpWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vlWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_isXSTrap <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_waitForward <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_blockBackward <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_flushPipe <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vill <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vma <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vta <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vsew <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vlmul <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVill <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVma <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVta <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVsew <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVlmul <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vlsInstr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_wfflags <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_isMove <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_isVset <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_firstUop <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_lastUop <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_numWB <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_commitType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_instrSize <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_dirtyFs <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_dirtyVs <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_traceBlockInPipe_itype <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_traceBlockInPipe_iretire <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_traceBlockInPipe_ilastsize <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_snapshot <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_lqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_sqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_singleStep <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_debug_sim_trig <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_valid <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_instr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_pc <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_0 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_1 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_3 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_12 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_20 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_22 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_isFetchMalAddr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_hasException <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_trigger <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_preDecodeInfo_isRVC <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_crossPageIPFFix <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_ftqPtr_flag <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_ftqPtr_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_ftqOffset <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_ldest <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_fuType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_fuOpType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_rfWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_fpWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vlWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_isXSTrap <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_waitForward <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_blockBackward <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_flushPipe <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vill <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vma <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vta <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vsew <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vlmul <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVill <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVma <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVta <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVsew <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVlmul <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vlsInstr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_wfflags <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_isMove <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_isVset <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_firstUop <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_lastUop <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_numWB <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_commitType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_instrSize <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_dirtyFs <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_dirtyVs <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_traceBlockInPipe_itype <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_traceBlockInPipe_iretire <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_traceBlockInPipe_ilastsize <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_snapshot <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_lqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_sqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_singleStep <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_debug_sim_trig <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_valid <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_instr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_pc <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_0 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_1 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_3 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_12 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_20 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_22 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_isFetchMalAddr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_hasException <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_trigger <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_preDecodeInfo_isRVC <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_crossPageIPFFix <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_ftqPtr_flag <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_ftqPtr_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_ftqOffset <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_ldest <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_fuType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_fuOpType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_rfWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_fpWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vlWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_isXSTrap <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_waitForward <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_blockBackward <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_flushPipe <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vill <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vma <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vta <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vsew <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vlmul <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVill <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVma <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVta <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVsew <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVlmul <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vlsInstr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_wfflags <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_isMove <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_isVset <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_firstUop <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_lastUop <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_numWB <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_commitType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_instrSize <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_dirtyFs <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_dirtyVs <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_traceBlockInPipe_itype <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_traceBlockInPipe_iretire <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_traceBlockInPipe_ilastsize <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_snapshot <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_lqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_sqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_singleStep <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_debug_sim_trig <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_valid <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_instr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_pc <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_0 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_1 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_3 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_12 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_20 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_22 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_isFetchMalAddr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_hasException <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_trigger <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_preDecodeInfo_isRVC <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_crossPageIPFFix <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_ftqPtr_flag <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_ftqPtr_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_ftqOffset <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_ldest <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_fuType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_fuOpType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_rfWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_fpWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vlWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_isXSTrap <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_waitForward <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_blockBackward <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_flushPipe <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vill <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vma <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vta <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vsew <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vlmul <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVill <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVma <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVta <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVsew <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVlmul <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vlsInstr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_wfflags <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_isMove <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_isVset <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_firstUop <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_lastUop <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_numWB <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_commitType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_instrSize <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_dirtyFs <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_dirtyVs <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_traceBlockInPipe_itype <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_traceBlockInPipe_iretire <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_traceBlockInPipe_ilastsize <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_snapshot <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_lqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_sqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_singleStep <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_debug_sim_trig <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_valid <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_instr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_pc <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_0 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_1 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_3 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_12 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_20 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_22 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_isFetchMalAddr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_hasException <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_trigger <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_preDecodeInfo_isRVC <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_crossPageIPFFix <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_ftqPtr_flag <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_ftqPtr_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_ftqOffset <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_ldest <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_fuType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_fuOpType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_rfWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_fpWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vlWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_isXSTrap <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_waitForward <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_blockBackward <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_flushPipe <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vill <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vma <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vta <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vsew <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vlmul <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVill <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVma <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVta <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVsew <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVlmul <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vlsInstr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_wfflags <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_isMove <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_isVset <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_firstUop <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_lastUop <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_numWB <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_commitType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_instrSize <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_dirtyFs <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_dirtyVs <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_traceBlockInPipe_itype <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_traceBlockInPipe_iretire <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_traceBlockInPipe_ilastsize <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_snapshot <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_lqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_sqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_singleStep <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_debug_sim_trig <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_valid <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_instr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_pc <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_0 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_1 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_3 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_12 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_20 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_22 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_isFetchMalAddr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_hasException <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_trigger <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_preDecodeInfo_isRVC <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_crossPageIPFFix <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_ftqPtr_flag <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_ftqPtr_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_ftqOffset <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_ldest <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_fuType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_fuOpType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_rfWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_fpWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vlWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_isXSTrap <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_waitForward <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_blockBackward <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_flushPipe <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vill <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vma <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vta <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vsew <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vlmul <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVill <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVma <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVta <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVsew <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVlmul <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vlsInstr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_wfflags <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_isMove <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_isVset <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_firstUop <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_lastUop <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_numWB <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_commitType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_instrSize <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_dirtyFs <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_dirtyVs <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_traceBlockInPipe_itype <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_traceBlockInPipe_iretire <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_traceBlockInPipe_ilastsize <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_snapshot <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_lqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_sqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_singleStep <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_debug_sim_trig <= '0;

    end
    else if(drv_mode==tcnt_dec_base::DRV_1) begin
        vif.drv_mp.drv_cb.clock <= '1;
        vif.drv_mp.drv_cb.reset <= '1;
        vif.drv_mp.drv_cb.io_hartId <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_valid <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_instr <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_pc <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_0 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_1 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_2 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_3 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_12 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_20 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_22 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_isFetchMalAddr <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_hasException <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_trigger <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_preDecodeInfo_isRVC <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_crossPageIPFFix <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_ftqPtr_flag <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_ftqPtr_value <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_ftqOffset <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_ldest <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_fuType <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_fuOpType <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_rfWen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_fpWen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vecWen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_v0Wen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vlWen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_isXSTrap <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_waitForward <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_blockBackward <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_flushPipe <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vill <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vma <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vta <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vsew <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vlmul <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVill <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVma <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVta <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVsew <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVlmul <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vlsInstr <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_wfflags <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_isMove <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_isVset <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_firstUop <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_lastUop <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_numWB <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_commitType <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_pdest <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_robIdx_flag <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_instrSize <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_dirtyFs <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_dirtyVs <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_traceBlockInPipe_itype <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_traceBlockInPipe_iretire <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_traceBlockInPipe_ilastsize <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_eliminatedMove <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_snapshot <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_lqIdx_value <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_sqIdx_value <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_singleStep <= '1;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_debug_sim_trig <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_valid <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_instr <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_pc <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_0 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_1 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_2 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_3 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_12 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_20 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_22 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_isFetchMalAddr <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_hasException <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_trigger <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_preDecodeInfo_isRVC <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_crossPageIPFFix <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_ftqPtr_flag <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_ftqPtr_value <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_ftqOffset <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_ldest <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_fuType <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_fuOpType <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_rfWen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_fpWen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vecWen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_v0Wen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vlWen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_isXSTrap <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_waitForward <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_blockBackward <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_flushPipe <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vill <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vma <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vta <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vsew <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vlmul <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVill <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVma <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVta <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVsew <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVlmul <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vlsInstr <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_wfflags <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_isMove <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_isVset <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_firstUop <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_lastUop <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_numWB <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_commitType <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_pdest <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_robIdx_flag <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_instrSize <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_dirtyFs <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_dirtyVs <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_traceBlockInPipe_itype <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_traceBlockInPipe_iretire <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_traceBlockInPipe_ilastsize <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_eliminatedMove <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_snapshot <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_lqIdx_value <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_sqIdx_value <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_singleStep <= '1;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_debug_sim_trig <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_valid <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_instr <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_pc <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_0 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_1 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_2 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_3 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_12 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_20 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_22 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_isFetchMalAddr <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_hasException <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_trigger <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_preDecodeInfo_isRVC <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_crossPageIPFFix <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_ftqPtr_flag <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_ftqPtr_value <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_ftqOffset <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_ldest <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_fuType <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_fuOpType <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_rfWen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_fpWen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vecWen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_v0Wen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vlWen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_isXSTrap <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_waitForward <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_blockBackward <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_flushPipe <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vill <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vma <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vta <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vsew <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vlmul <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVill <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVma <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVta <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVsew <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVlmul <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vlsInstr <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_wfflags <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_isMove <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_isVset <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_firstUop <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_lastUop <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_numWB <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_commitType <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_pdest <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_robIdx_flag <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_instrSize <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_dirtyFs <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_dirtyVs <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_traceBlockInPipe_itype <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_traceBlockInPipe_iretire <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_traceBlockInPipe_ilastsize <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_eliminatedMove <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_snapshot <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_lqIdx_value <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_sqIdx_value <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_singleStep <= '1;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_debug_sim_trig <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_valid <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_instr <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_pc <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_0 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_1 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_2 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_3 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_12 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_20 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_22 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_isFetchMalAddr <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_hasException <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_trigger <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_preDecodeInfo_isRVC <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_crossPageIPFFix <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_ftqPtr_flag <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_ftqPtr_value <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_ftqOffset <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_ldest <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_fuType <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_fuOpType <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_rfWen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_fpWen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vecWen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_v0Wen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vlWen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_isXSTrap <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_waitForward <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_blockBackward <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_flushPipe <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vill <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vma <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vta <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vsew <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vlmul <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVill <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVma <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVta <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVsew <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVlmul <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vlsInstr <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_wfflags <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_isMove <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_isVset <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_firstUop <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_lastUop <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_numWB <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_commitType <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_pdest <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_robIdx_flag <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_instrSize <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_dirtyFs <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_dirtyVs <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_traceBlockInPipe_itype <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_traceBlockInPipe_iretire <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_traceBlockInPipe_ilastsize <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_eliminatedMove <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_snapshot <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_lqIdx_value <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_sqIdx_value <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_singleStep <= '1;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_debug_sim_trig <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_valid <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_instr <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_pc <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_0 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_1 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_2 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_3 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_12 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_20 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_22 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_isFetchMalAddr <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_hasException <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_trigger <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_preDecodeInfo_isRVC <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_crossPageIPFFix <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_ftqPtr_flag <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_ftqPtr_value <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_ftqOffset <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_ldest <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_fuType <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_fuOpType <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_rfWen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_fpWen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vecWen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_v0Wen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vlWen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_isXSTrap <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_waitForward <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_blockBackward <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_flushPipe <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vill <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vma <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vta <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vsew <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vlmul <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVill <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVma <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVta <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVsew <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVlmul <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vlsInstr <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_wfflags <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_isMove <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_isVset <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_firstUop <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_lastUop <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_numWB <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_commitType <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_pdest <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_robIdx_flag <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_instrSize <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_dirtyFs <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_dirtyVs <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_traceBlockInPipe_itype <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_traceBlockInPipe_iretire <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_traceBlockInPipe_ilastsize <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_eliminatedMove <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_snapshot <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_lqIdx_value <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_sqIdx_value <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_singleStep <= '1;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_debug_sim_trig <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_valid <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_instr <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_pc <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_0 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_1 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_2 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_3 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_12 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_20 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_22 <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_isFetchMalAddr <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_hasException <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_trigger <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_preDecodeInfo_isRVC <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_crossPageIPFFix <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_ftqPtr_flag <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_ftqPtr_value <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_ftqOffset <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_ldest <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_fuType <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_fuOpType <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_rfWen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_fpWen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vecWen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_v0Wen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vlWen <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_isXSTrap <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_waitForward <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_blockBackward <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_flushPipe <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vill <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vma <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vta <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vsew <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vlmul <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVill <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVma <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVta <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVsew <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVlmul <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vlsInstr <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_wfflags <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_isMove <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_isVset <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_firstUop <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_lastUop <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_numWB <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_commitType <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_pdest <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_robIdx_flag <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_instrSize <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_dirtyFs <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_dirtyVs <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_traceBlockInPipe_itype <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_traceBlockInPipe_iretire <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_traceBlockInPipe_ilastsize <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_eliminatedMove <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_snapshot <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_lqIdx_value <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_sqIdx_value <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_singleStep <= '1;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_debug_sim_trig <= '1;

    end
    else if(drv_mode==tcnt_dec_base::DRV_X) begin
        vif.drv_mp.drv_cb.clock <= 'x;
        vif.drv_mp.drv_cb.reset <= 'x;
        vif.drv_mp.drv_cb.io_hartId <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_valid <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_instr <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_pc <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_0 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_1 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_2 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_3 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_12 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_20 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_22 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_isFetchMalAddr <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_hasException <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_trigger <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_preDecodeInfo_isRVC <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_crossPageIPFFix <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_ftqPtr_flag <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_ftqPtr_value <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_ftqOffset <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_ldest <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_fuType <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_fuOpType <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_rfWen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_fpWen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vecWen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_v0Wen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vlWen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_isXSTrap <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_waitForward <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_blockBackward <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_flushPipe <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vill <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vma <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vta <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vsew <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vlmul <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVill <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVma <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVta <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVsew <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVlmul <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vlsInstr <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_wfflags <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_isMove <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_isVset <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_firstUop <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_lastUop <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_numWB <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_commitType <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_pdest <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_robIdx_flag <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_instrSize <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_dirtyFs <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_dirtyVs <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_traceBlockInPipe_itype <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_traceBlockInPipe_iretire <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_traceBlockInPipe_ilastsize <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_eliminatedMove <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_snapshot <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_lqIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_sqIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_singleStep <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_debug_sim_trig <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_valid <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_instr <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_pc <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_0 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_1 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_2 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_3 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_12 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_20 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_22 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_isFetchMalAddr <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_hasException <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_trigger <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_preDecodeInfo_isRVC <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_crossPageIPFFix <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_ftqPtr_flag <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_ftqPtr_value <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_ftqOffset <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_ldest <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_fuType <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_fuOpType <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_rfWen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_fpWen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vecWen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_v0Wen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vlWen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_isXSTrap <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_waitForward <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_blockBackward <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_flushPipe <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vill <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vma <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vta <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vsew <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vlmul <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVill <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVma <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVta <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVsew <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVlmul <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vlsInstr <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_wfflags <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_isMove <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_isVset <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_firstUop <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_lastUop <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_numWB <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_commitType <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_pdest <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_robIdx_flag <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_instrSize <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_dirtyFs <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_dirtyVs <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_traceBlockInPipe_itype <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_traceBlockInPipe_iretire <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_traceBlockInPipe_ilastsize <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_eliminatedMove <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_snapshot <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_lqIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_sqIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_singleStep <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_debug_sim_trig <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_valid <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_instr <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_pc <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_0 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_1 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_2 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_3 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_12 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_20 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_22 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_isFetchMalAddr <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_hasException <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_trigger <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_preDecodeInfo_isRVC <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_crossPageIPFFix <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_ftqPtr_flag <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_ftqPtr_value <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_ftqOffset <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_ldest <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_fuType <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_fuOpType <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_rfWen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_fpWen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vecWen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_v0Wen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vlWen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_isXSTrap <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_waitForward <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_blockBackward <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_flushPipe <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vill <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vma <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vta <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vsew <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vlmul <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVill <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVma <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVta <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVsew <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVlmul <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vlsInstr <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_wfflags <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_isMove <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_isVset <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_firstUop <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_lastUop <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_numWB <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_commitType <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_pdest <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_robIdx_flag <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_instrSize <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_dirtyFs <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_dirtyVs <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_traceBlockInPipe_itype <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_traceBlockInPipe_iretire <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_traceBlockInPipe_ilastsize <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_eliminatedMove <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_snapshot <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_lqIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_sqIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_singleStep <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_debug_sim_trig <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_valid <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_instr <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_pc <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_0 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_1 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_2 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_3 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_12 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_20 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_22 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_isFetchMalAddr <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_hasException <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_trigger <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_preDecodeInfo_isRVC <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_crossPageIPFFix <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_ftqPtr_flag <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_ftqPtr_value <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_ftqOffset <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_ldest <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_fuType <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_fuOpType <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_rfWen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_fpWen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vecWen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_v0Wen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vlWen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_isXSTrap <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_waitForward <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_blockBackward <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_flushPipe <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vill <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vma <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vta <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vsew <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vlmul <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVill <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVma <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVta <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVsew <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVlmul <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vlsInstr <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_wfflags <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_isMove <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_isVset <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_firstUop <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_lastUop <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_numWB <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_commitType <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_pdest <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_robIdx_flag <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_instrSize <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_dirtyFs <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_dirtyVs <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_traceBlockInPipe_itype <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_traceBlockInPipe_iretire <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_traceBlockInPipe_ilastsize <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_eliminatedMove <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_snapshot <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_lqIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_sqIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_singleStep <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_debug_sim_trig <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_valid <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_instr <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_pc <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_0 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_1 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_2 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_3 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_12 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_20 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_22 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_isFetchMalAddr <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_hasException <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_trigger <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_preDecodeInfo_isRVC <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_crossPageIPFFix <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_ftqPtr_flag <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_ftqPtr_value <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_ftqOffset <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_ldest <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_fuType <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_fuOpType <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_rfWen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_fpWen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vecWen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_v0Wen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vlWen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_isXSTrap <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_waitForward <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_blockBackward <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_flushPipe <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vill <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vma <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vta <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vsew <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vlmul <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVill <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVma <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVta <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVsew <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVlmul <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vlsInstr <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_wfflags <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_isMove <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_isVset <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_firstUop <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_lastUop <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_numWB <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_commitType <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_pdest <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_robIdx_flag <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_instrSize <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_dirtyFs <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_dirtyVs <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_traceBlockInPipe_itype <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_traceBlockInPipe_iretire <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_traceBlockInPipe_ilastsize <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_eliminatedMove <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_snapshot <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_lqIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_sqIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_singleStep <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_debug_sim_trig <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_valid <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_instr <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_pc <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_0 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_1 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_2 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_3 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_12 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_20 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_22 <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_isFetchMalAddr <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_hasException <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_trigger <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_preDecodeInfo_isRVC <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_crossPageIPFFix <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_ftqPtr_flag <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_ftqPtr_value <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_ftqOffset <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_ldest <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_fuType <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_fuOpType <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_rfWen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_fpWen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vecWen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_v0Wen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vlWen <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_isXSTrap <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_waitForward <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_blockBackward <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_flushPipe <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vill <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vma <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vta <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vsew <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vlmul <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVill <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVma <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVta <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVsew <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVlmul <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vlsInstr <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_wfflags <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_isMove <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_isVset <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_firstUop <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_lastUop <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_numWB <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_commitType <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_pdest <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_robIdx_flag <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_instrSize <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_dirtyFs <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_dirtyVs <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_traceBlockInPipe_itype <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_traceBlockInPipe_iretire <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_traceBlockInPipe_ilastsize <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_eliminatedMove <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_snapshot <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_lqIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_sqIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_singleStep <= 'x;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_debug_sim_trig <= 'x;

    end
    else if(drv_mode==tcnt_dec_base::DRV_RAND) begin
        vif.drv_mp.drv_cb.clock <= $urandom;
        vif.drv_mp.drv_cb.reset <= $urandom;
        vif.drv_mp.drv_cb.io_hartId <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_valid <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_instr <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_pc <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_0 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_1 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_2 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_3 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_12 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_20 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_22 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_isFetchMalAddr <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_hasException <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_trigger <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_preDecodeInfo_isRVC <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_crossPageIPFFix <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_ftqPtr_flag <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_ftqPtr_value <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_ftqOffset <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_ldest <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_fuType <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_fuOpType <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_rfWen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_fpWen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vecWen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_v0Wen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vlWen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_isXSTrap <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_waitForward <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_blockBackward <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_flushPipe <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vill <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vma <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vta <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vsew <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vlmul <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVill <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVma <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVta <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVsew <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVlmul <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vlsInstr <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_wfflags <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_isMove <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_isVset <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_firstUop <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_lastUop <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_numWB <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_commitType <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_pdest <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_robIdx_flag <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_instrSize <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_dirtyFs <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_dirtyVs <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_traceBlockInPipe_itype <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_traceBlockInPipe_iretire <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_traceBlockInPipe_ilastsize <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_eliminatedMove <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_snapshot <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_lqIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_sqIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_singleStep <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_debug_sim_trig <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_valid <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_instr <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_pc <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_0 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_1 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_2 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_3 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_12 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_20 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_22 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_isFetchMalAddr <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_hasException <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_trigger <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_preDecodeInfo_isRVC <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_crossPageIPFFix <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_ftqPtr_flag <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_ftqPtr_value <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_ftqOffset <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_ldest <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_fuType <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_fuOpType <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_rfWen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_fpWen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vecWen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_v0Wen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vlWen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_isXSTrap <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_waitForward <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_blockBackward <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_flushPipe <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vill <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vma <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vta <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vsew <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vlmul <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVill <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVma <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVta <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVsew <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVlmul <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vlsInstr <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_wfflags <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_isMove <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_isVset <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_firstUop <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_lastUop <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_numWB <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_commitType <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_pdest <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_robIdx_flag <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_instrSize <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_dirtyFs <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_dirtyVs <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_traceBlockInPipe_itype <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_traceBlockInPipe_iretire <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_traceBlockInPipe_ilastsize <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_eliminatedMove <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_snapshot <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_lqIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_sqIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_singleStep <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_debug_sim_trig <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_valid <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_instr <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_pc <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_0 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_1 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_2 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_3 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_12 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_20 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_22 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_isFetchMalAddr <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_hasException <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_trigger <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_preDecodeInfo_isRVC <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_crossPageIPFFix <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_ftqPtr_flag <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_ftqPtr_value <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_ftqOffset <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_ldest <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_fuType <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_fuOpType <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_rfWen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_fpWen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vecWen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_v0Wen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vlWen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_isXSTrap <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_waitForward <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_blockBackward <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_flushPipe <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vill <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vma <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vta <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vsew <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vlmul <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVill <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVma <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVta <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVsew <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVlmul <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vlsInstr <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_wfflags <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_isMove <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_isVset <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_firstUop <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_lastUop <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_numWB <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_commitType <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_pdest <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_robIdx_flag <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_instrSize <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_dirtyFs <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_dirtyVs <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_traceBlockInPipe_itype <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_traceBlockInPipe_iretire <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_traceBlockInPipe_ilastsize <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_eliminatedMove <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_snapshot <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_lqIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_sqIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_singleStep <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_debug_sim_trig <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_valid <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_instr <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_pc <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_0 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_1 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_2 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_3 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_12 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_20 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_22 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_isFetchMalAddr <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_hasException <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_trigger <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_preDecodeInfo_isRVC <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_crossPageIPFFix <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_ftqPtr_flag <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_ftqPtr_value <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_ftqOffset <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_ldest <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_fuType <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_fuOpType <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_rfWen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_fpWen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vecWen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_v0Wen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vlWen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_isXSTrap <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_waitForward <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_blockBackward <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_flushPipe <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vill <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vma <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vta <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vsew <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vlmul <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVill <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVma <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVta <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVsew <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVlmul <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vlsInstr <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_wfflags <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_isMove <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_isVset <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_firstUop <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_lastUop <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_numWB <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_commitType <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_pdest <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_robIdx_flag <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_instrSize <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_dirtyFs <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_dirtyVs <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_traceBlockInPipe_itype <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_traceBlockInPipe_iretire <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_traceBlockInPipe_ilastsize <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_eliminatedMove <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_snapshot <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_lqIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_sqIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_singleStep <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_debug_sim_trig <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_valid <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_instr <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_pc <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_0 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_1 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_2 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_3 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_12 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_20 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_22 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_isFetchMalAddr <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_hasException <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_trigger <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_preDecodeInfo_isRVC <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_crossPageIPFFix <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_ftqPtr_flag <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_ftqPtr_value <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_ftqOffset <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_ldest <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_fuType <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_fuOpType <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_rfWen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_fpWen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vecWen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_v0Wen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vlWen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_isXSTrap <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_waitForward <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_blockBackward <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_flushPipe <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vill <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vma <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vta <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vsew <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vlmul <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVill <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVma <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVta <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVsew <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVlmul <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vlsInstr <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_wfflags <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_isMove <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_isVset <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_firstUop <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_lastUop <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_numWB <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_commitType <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_pdest <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_robIdx_flag <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_instrSize <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_dirtyFs <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_dirtyVs <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_traceBlockInPipe_itype <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_traceBlockInPipe_iretire <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_traceBlockInPipe_ilastsize <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_eliminatedMove <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_snapshot <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_lqIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_sqIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_singleStep <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_debug_sim_trig <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_valid <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_instr <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_pc <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_0 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_1 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_2 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_3 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_12 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_20 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_22 <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_isFetchMalAddr <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_hasException <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_trigger <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_preDecodeInfo_isRVC <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_crossPageIPFFix <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_ftqPtr_flag <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_ftqPtr_value <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_ftqOffset <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_ldest <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_fuType <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_fuOpType <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_rfWen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_fpWen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vecWen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_v0Wen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vlWen <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_isXSTrap <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_waitForward <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_blockBackward <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_flushPipe <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vill <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vma <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vta <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vsew <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vlmul <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVill <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVma <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVta <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVsew <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVlmul <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vlsInstr <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_wfflags <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_isMove <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_isVset <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_firstUop <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_lastUop <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_numWB <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_commitType <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_pdest <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_robIdx_flag <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_instrSize <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_dirtyFs <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_dirtyVs <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_traceBlockInPipe_itype <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_traceBlockInPipe_iretire <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_traceBlockInPipe_ilastsize <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_eliminatedMove <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_snapshot <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_lqIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_sqIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_singleStep <= $urandom;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_debug_sim_trig <= $urandom;

    end
    else if(drv_mode==tcnt_dec_base::DRV_LST) begin
        vif.drv_mp.drv_cb.clock <= '0;
        vif.drv_mp.drv_cb.reset <= '0;
        vif.drv_mp.drv_cb.io_hartId <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_valid <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_instr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_pc <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_0 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_1 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_3 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_12 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_20 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_exceptionVec_22 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_isFetchMalAddr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_hasException <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_trigger <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_preDecodeInfo_isRVC <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_crossPageIPFFix <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_ftqPtr_flag <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_ftqPtr_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_ftqOffset <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_ldest <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_fuType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_fuOpType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_rfWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_fpWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vlWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_isXSTrap <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_waitForward <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_blockBackward <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_flushPipe <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vill <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vma <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vta <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vsew <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_vlmul <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVill <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVma <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVta <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVsew <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vpu_specVlmul <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_vlsInstr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_wfflags <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_isMove <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_isVset <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_firstUop <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_lastUop <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_numWB <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_commitType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_instrSize <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_dirtyFs <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_dirtyVs <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_traceBlockInPipe_itype <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_traceBlockInPipe_iretire <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_traceBlockInPipe_ilastsize <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_snapshot <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_lqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_sqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_singleStep <= '0;
        vif.drv_mp.drv_cb.io_enq_req_0_bits_debug_sim_trig <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_valid <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_instr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_pc <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_0 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_1 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_3 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_12 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_20 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_exceptionVec_22 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_isFetchMalAddr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_hasException <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_trigger <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_preDecodeInfo_isRVC <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_crossPageIPFFix <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_ftqPtr_flag <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_ftqPtr_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_ftqOffset <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_ldest <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_fuType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_fuOpType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_rfWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_fpWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vlWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_isXSTrap <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_waitForward <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_blockBackward <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_flushPipe <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vill <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vma <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vta <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vsew <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_vlmul <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVill <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVma <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVta <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVsew <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vpu_specVlmul <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_vlsInstr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_wfflags <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_isMove <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_isVset <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_firstUop <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_lastUop <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_numWB <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_commitType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_instrSize <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_dirtyFs <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_dirtyVs <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_traceBlockInPipe_itype <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_traceBlockInPipe_iretire <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_traceBlockInPipe_ilastsize <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_snapshot <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_lqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_sqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_singleStep <= '0;
        vif.drv_mp.drv_cb.io_enq_req_1_bits_debug_sim_trig <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_valid <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_instr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_pc <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_0 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_1 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_3 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_12 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_20 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_exceptionVec_22 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_isFetchMalAddr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_hasException <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_trigger <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_preDecodeInfo_isRVC <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_crossPageIPFFix <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_ftqPtr_flag <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_ftqPtr_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_ftqOffset <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_ldest <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_fuType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_fuOpType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_rfWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_fpWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vlWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_isXSTrap <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_waitForward <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_blockBackward <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_flushPipe <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vill <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vma <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vta <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vsew <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_vlmul <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVill <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVma <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVta <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVsew <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vpu_specVlmul <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_vlsInstr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_wfflags <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_isMove <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_isVset <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_firstUop <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_lastUop <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_numWB <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_commitType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_instrSize <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_dirtyFs <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_dirtyVs <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_traceBlockInPipe_itype <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_traceBlockInPipe_iretire <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_traceBlockInPipe_ilastsize <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_snapshot <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_lqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_sqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_singleStep <= '0;
        vif.drv_mp.drv_cb.io_enq_req_2_bits_debug_sim_trig <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_valid <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_instr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_pc <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_0 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_1 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_3 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_12 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_20 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_exceptionVec_22 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_isFetchMalAddr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_hasException <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_trigger <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_preDecodeInfo_isRVC <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_crossPageIPFFix <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_ftqPtr_flag <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_ftqPtr_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_ftqOffset <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_ldest <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_fuType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_fuOpType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_rfWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_fpWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vlWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_isXSTrap <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_waitForward <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_blockBackward <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_flushPipe <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vill <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vma <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vta <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vsew <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_vlmul <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVill <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVma <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVta <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVsew <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vpu_specVlmul <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_vlsInstr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_wfflags <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_isMove <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_isVset <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_firstUop <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_lastUop <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_numWB <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_commitType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_instrSize <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_dirtyFs <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_dirtyVs <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_traceBlockInPipe_itype <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_traceBlockInPipe_iretire <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_traceBlockInPipe_ilastsize <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_snapshot <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_lqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_sqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_singleStep <= '0;
        vif.drv_mp.drv_cb.io_enq_req_3_bits_debug_sim_trig <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_valid <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_instr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_pc <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_0 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_1 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_3 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_12 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_20 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_exceptionVec_22 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_isFetchMalAddr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_hasException <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_trigger <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_preDecodeInfo_isRVC <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_crossPageIPFFix <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_ftqPtr_flag <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_ftqPtr_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_ftqOffset <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_ldest <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_fuType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_fuOpType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_rfWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_fpWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vlWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_isXSTrap <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_waitForward <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_blockBackward <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_flushPipe <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vill <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vma <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vta <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vsew <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_vlmul <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVill <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVma <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVta <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVsew <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vpu_specVlmul <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_vlsInstr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_wfflags <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_isMove <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_isVset <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_firstUop <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_lastUop <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_numWB <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_commitType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_instrSize <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_dirtyFs <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_dirtyVs <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_traceBlockInPipe_itype <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_traceBlockInPipe_iretire <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_traceBlockInPipe_ilastsize <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_snapshot <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_lqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_sqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_singleStep <= '0;
        vif.drv_mp.drv_cb.io_enq_req_4_bits_debug_sim_trig <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_valid <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_instr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_pc <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_0 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_1 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_3 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_12 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_20 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_exceptionVec_22 <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_isFetchMalAddr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_hasException <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_trigger <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_preDecodeInfo_isRVC <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_crossPageIPFFix <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_ftqPtr_flag <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_ftqPtr_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_ftqOffset <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_ldest <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_fuType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_fuOpType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_rfWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_fpWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vlWen <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_isXSTrap <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_waitForward <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_blockBackward <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_flushPipe <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vill <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vma <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vta <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vsew <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_vlmul <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVill <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVma <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVta <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVsew <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vpu_specVlmul <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_vlsInstr <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_wfflags <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_isMove <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_isVset <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_firstUop <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_lastUop <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_numWB <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_commitType <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_instrSize <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_dirtyFs <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_dirtyVs <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_traceBlockInPipe_itype <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_traceBlockInPipe_iretire <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_traceBlockInPipe_ilastsize <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_snapshot <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_lqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_sqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_singleStep <= '0;
        vif.drv_mp.drv_cb.io_enq_req_5_bits_debug_sim_trig <= '0;

    end

endtask:drive_idle

`endif


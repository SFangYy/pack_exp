//=========================================================
//File name    : Rob_output_agent_pkg.sv
//Author       : nanyunhao
//Module name  : Rob_output_agent_pkg
//Discribution : Rob_output_agent_pkg : package
//Date         : 2026-01-22
//=========================================================
`ifndef ROB_OUTPUT_AGENT_PKG__SV
`define ROB_OUTPUT_AGENT_PKG__SV

`ifndef TCNT_HAD_INCLUDE_UVM_MACROS
`define TCNT_HAD_INCLUDE_UVM_MACROS
    `include "uvm_macros.svh"
`endif

`include "Rob_output_agent_dec.sv"
`include "Rob_output_agent_interface.sv"
package Rob_output_agent_pkg;

    import uvm_pkg::*;
    import tcnt_realtime::*;
    import tcnt_dec_base::*;
    import tcnt_common_method::*;
    import tcnt_base_pkg::*;

    import Rob_output_agent_dec::*;

    `include "Rob_output_agent_cfg.sv"
    `include "Rob_output_agent_xaction.sv"
    `include "Rob_output_agent_default_sequence.sv"
    `include "Rob_output_agent_driver.sv"
    `include "Rob_output_agent_monitor.sv"
    `include "Rob_output_agent_sequencer.sv"
    `include "Rob_output_agent.sv"

endpackage

import Rob_output_agent_pkg::*;

`endif


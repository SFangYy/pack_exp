`ifndef SV_MAIN__SV
`define SV_MAIN__SV

module sv_main;
    // Import top_tb module
    `include "top_tb.sv"
endmodule

`endif
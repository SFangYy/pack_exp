//=========================================================
//File name    : Rob_output_agent_monitor.sv
//Author       : nanyunhao
//Module name  : Rob_output_agent_monitor
//Discribution : Rob_output_agent_monitor : monitor
//Date         : 2026-01-22
//=========================================================
`ifndef ROB_OUTPUT_AGENT_MONITOR__SV
`define ROB_OUTPUT_AGENT_MONITOR__SV

class Rob_output_agent_monitor  extends tcnt_monitor_base#(virtual Rob_output_agent_interface,Rob_output_agent_cfg,Rob_output_agent_xaction);

    `uvm_component_utils(Rob_output_agent_monitor)

    extern function new(string name, uvm_component parent);
    extern virtual function void build_phase(uvm_phase phase);
    extern task run_phase(uvm_phase phase);
    extern task mon_data();
endclass:Rob_output_agent_monitor

function Rob_output_agent_monitor::new(string name, uvm_component parent);
    super.new(name,parent);
endfunction:new

function void Rob_output_agent_monitor::build_phase(uvm_phase phase);
    super.build_phase(phase);
endfunction:build_phase

task Rob_output_agent_monitor::run_phase(uvm_phase phase);
    super.run_phase(phase);
    this.mon_data();
endtask:run_phase

task Rob_output_agent_monitor::mon_data();

    logic         io_enq_canAccept     ;
    logic         io_enq_canAcceptForDispatch;
    logic         io_enq_isEmpty       ;
    logic         io_flushOut_valid    ;
    logic         io_flushOut_bits_isRVC;
    logic         io_flushOut_bits_robIdx_flag;
    logic [7:0]   io_flushOut_bits_robIdx_value;
    logic         io_flushOut_bits_ftqIdx_flag;
    logic [5:0]   io_flushOut_bits_ftqIdx_value;
    logic [3:0]   io_flushOut_bits_ftqOffset;
    logic         io_flushOut_bits_level;
    logic         io_exception_valid   ;
    logic [31:0]  io_exception_bits_instr;
    logic [2:0]   io_exception_bits_commitType;
    logic         io_exception_bits_exceptionVec_0;
    logic         io_exception_bits_exceptionVec_1;
    logic         io_exception_bits_exceptionVec_2;
    logic         io_exception_bits_exceptionVec_3;
    logic         io_exception_bits_exceptionVec_4;
    logic         io_exception_bits_exceptionVec_5;
    logic         io_exception_bits_exceptionVec_6;
    logic         io_exception_bits_exceptionVec_7;
    logic         io_exception_bits_exceptionVec_8;
    logic         io_exception_bits_exceptionVec_9;
    logic         io_exception_bits_exceptionVec_10;
    logic         io_exception_bits_exceptionVec_11;
    logic         io_exception_bits_exceptionVec_12;
    logic         io_exception_bits_exceptionVec_13;
    logic         io_exception_bits_exceptionVec_14;
    logic         io_exception_bits_exceptionVec_15;
    logic         io_exception_bits_exceptionVec_16;
    logic         io_exception_bits_exceptionVec_17;
    logic         io_exception_bits_exceptionVec_18;
    logic         io_exception_bits_exceptionVec_19;
    logic         io_exception_bits_exceptionVec_20;
    logic         io_exception_bits_exceptionVec_21;
    logic         io_exception_bits_exceptionVec_22;
    logic         io_exception_bits_exceptionVec_23;
    logic         io_exception_bits_isPcBkpt;
    logic         io_exception_bits_isFetchMalAddr;
    logic [63:0]  io_exception_bits_gpaddr;
    logic         io_exception_bits_singleStep;
    logic         io_exception_bits_crossPageIPFFix;
    logic         io_exception_bits_isInterrupt;
    logic         io_exception_bits_isHls;
    logic [3:0]   io_exception_bits_trigger;
    logic         io_exception_bits_isForVSnonLeafPTE;
    logic         io_commits_isCommit  ;
    logic         io_commits_commitValid_0;
    logic         io_commits_commitValid_1;
    logic         io_commits_commitValid_2;
    logic         io_commits_commitValid_3;
    logic         io_commits_commitValid_4;
    logic         io_commits_commitValid_5;
    logic         io_commits_commitValid_6;
    logic         io_commits_commitValid_7;
    logic         io_commits_isWalk    ;
    logic         io_commits_walkValid_0;
    logic         io_commits_walkValid_1;
    logic         io_commits_walkValid_2;
    logic         io_commits_walkValid_3;
    logic         io_commits_walkValid_4;
    logic         io_commits_walkValid_5;
    logic         io_commits_walkValid_6;
    logic         io_commits_walkValid_7;
    logic         io_commits_info_0_walk_v;
    logic         io_commits_info_0_commit_v;
    logic         io_commits_info_0_commit_w;
    logic [6:0]   io_commits_info_0_realDestSize;
    logic         io_commits_info_0_interrupt_safe;
    logic         io_commits_info_0_wflags;
    logic [4:0]   io_commits_info_0_fflags;
    logic         io_commits_info_0_vxsat;
    logic         io_commits_info_0_isRVC;
    logic         io_commits_info_0_isVset;
    logic         io_commits_info_0_isHls;
    logic         io_commits_info_0_isVls;
    logic         io_commits_info_0_vls;
    logic         io_commits_info_0_mmio;
    logic [2:0]   io_commits_info_0_commitType;
    logic         io_commits_info_0_ftqIdx_flag;
    logic [5:0]   io_commits_info_0_ftqIdx_value;
    logic [3:0]   io_commits_info_0_ftqOffset;
    logic [2:0]   io_commits_info_0_instrSize;
    logic         io_commits_info_0_fpWen;
    logic         io_commits_info_0_rfWen;
    logic         io_commits_info_0_needFlush;
    logic [3:0]   io_commits_info_0_traceBlockInPipe_itype;
    logic [3:0]   io_commits_info_0_traceBlockInPipe_iretire;
    logic         io_commits_info_0_traceBlockInPipe_ilastsize;
    logic [49:0]  io_commits_info_0_debug_pc;
    logic [31:0]  io_commits_info_0_debug_instr;
    logic [5:0]   io_commits_info_0_debug_ldest;
    logic [7:0]   io_commits_info_0_debug_pdest;
    logic [7:0]   io_commits_info_0_debug_otherPdest_0;
    logic [7:0]   io_commits_info_0_debug_otherPdest_1;
    logic [7:0]   io_commits_info_0_debug_otherPdest_2;
    logic [7:0]   io_commits_info_0_debug_otherPdest_3;
    logic [7:0]   io_commits_info_0_debug_otherPdest_4;
    logic [7:0]   io_commits_info_0_debug_otherPdest_5;
    logic [7:0]   io_commits_info_0_debug_otherPdest_6;
    logic [34:0]  io_commits_info_0_debug_fuType;
    logic         io_commits_info_0_dirtyFs;
    logic         io_commits_info_0_dirtyVs;
    logic         io_commits_info_1_walk_v;
    logic         io_commits_info_1_commit_v;
    logic         io_commits_info_1_commit_w;
    logic [6:0]   io_commits_info_1_realDestSize;
    logic         io_commits_info_1_interrupt_safe;
    logic         io_commits_info_1_wflags;
    logic [4:0]   io_commits_info_1_fflags;
    logic         io_commits_info_1_vxsat;
    logic         io_commits_info_1_isRVC;
    logic         io_commits_info_1_isVset;
    logic         io_commits_info_1_isHls;
    logic         io_commits_info_1_isVls;
    logic         io_commits_info_1_vls;
    logic         io_commits_info_1_mmio;
    logic [2:0]   io_commits_info_1_commitType;
    logic         io_commits_info_1_ftqIdx_flag;
    logic [5:0]   io_commits_info_1_ftqIdx_value;
    logic [3:0]   io_commits_info_1_ftqOffset;
    logic [2:0]   io_commits_info_1_instrSize;
    logic         io_commits_info_1_fpWen;
    logic         io_commits_info_1_rfWen;
    logic         io_commits_info_1_needFlush;
    logic [3:0]   io_commits_info_1_traceBlockInPipe_itype;
    logic [3:0]   io_commits_info_1_traceBlockInPipe_iretire;
    logic         io_commits_info_1_traceBlockInPipe_ilastsize;
    logic [49:0]  io_commits_info_1_debug_pc;
    logic [31:0]  io_commits_info_1_debug_instr;
    logic [5:0]   io_commits_info_1_debug_ldest;
    logic [7:0]   io_commits_info_1_debug_pdest;
    logic [7:0]   io_commits_info_1_debug_otherPdest_0;
    logic [7:0]   io_commits_info_1_debug_otherPdest_1;
    logic [7:0]   io_commits_info_1_debug_otherPdest_2;
    logic [7:0]   io_commits_info_1_debug_otherPdest_3;
    logic [7:0]   io_commits_info_1_debug_otherPdest_4;
    logic [7:0]   io_commits_info_1_debug_otherPdest_5;
    logic [7:0]   io_commits_info_1_debug_otherPdest_6;
    logic [34:0]  io_commits_info_1_debug_fuType;
    logic         io_commits_info_1_dirtyFs;
    logic         io_commits_info_1_dirtyVs;
    logic         io_commits_info_2_walk_v;
    logic         io_commits_info_2_commit_v;
    logic         io_commits_info_2_commit_w;
    logic [6:0]   io_commits_info_2_realDestSize;
    logic         io_commits_info_2_interrupt_safe;
    logic         io_commits_info_2_wflags;
    logic [4:0]   io_commits_info_2_fflags;
    logic         io_commits_info_2_vxsat;
    logic         io_commits_info_2_isRVC;
    logic         io_commits_info_2_isVset;
    logic         io_commits_info_2_isHls;
    logic         io_commits_info_2_isVls;
    logic         io_commits_info_2_vls;
    logic         io_commits_info_2_mmio;
    logic [2:0]   io_commits_info_2_commitType;
    logic         io_commits_info_2_ftqIdx_flag;
    logic [5:0]   io_commits_info_2_ftqIdx_value;
    logic [3:0]   io_commits_info_2_ftqOffset;
    logic [2:0]   io_commits_info_2_instrSize;
    logic         io_commits_info_2_fpWen;
    logic         io_commits_info_2_rfWen;
    logic         io_commits_info_2_needFlush;
    logic [3:0]   io_commits_info_2_traceBlockInPipe_itype;
    logic [3:0]   io_commits_info_2_traceBlockInPipe_iretire;
    logic         io_commits_info_2_traceBlockInPipe_ilastsize;
    logic [49:0]  io_commits_info_2_debug_pc;
    logic [31:0]  io_commits_info_2_debug_instr;
    logic [5:0]   io_commits_info_2_debug_ldest;
    logic [7:0]   io_commits_info_2_debug_pdest;
    logic [7:0]   io_commits_info_2_debug_otherPdest_0;
    logic [7:0]   io_commits_info_2_debug_otherPdest_1;
    logic [7:0]   io_commits_info_2_debug_otherPdest_2;
    logic [7:0]   io_commits_info_2_debug_otherPdest_3;
    logic [7:0]   io_commits_info_2_debug_otherPdest_4;
    logic [7:0]   io_commits_info_2_debug_otherPdest_5;
    logic [7:0]   io_commits_info_2_debug_otherPdest_6;
    logic [34:0]  io_commits_info_2_debug_fuType;
    logic         io_commits_info_2_dirtyFs;
    logic         io_commits_info_2_dirtyVs;
    logic         io_commits_info_3_walk_v;
    logic         io_commits_info_3_commit_v;
    logic         io_commits_info_3_commit_w;
    logic [6:0]   io_commits_info_3_realDestSize;
    logic         io_commits_info_3_interrupt_safe;
    logic         io_commits_info_3_wflags;
    logic [4:0]   io_commits_info_3_fflags;
    logic         io_commits_info_3_vxsat;
    logic         io_commits_info_3_isRVC;
    logic         io_commits_info_3_isVset;
    logic         io_commits_info_3_isHls;
    logic         io_commits_info_3_isVls;
    logic         io_commits_info_3_vls;
    logic         io_commits_info_3_mmio;
    logic [2:0]   io_commits_info_3_commitType;
    logic         io_commits_info_3_ftqIdx_flag;
    logic [5:0]   io_commits_info_3_ftqIdx_value;
    logic [3:0]   io_commits_info_3_ftqOffset;
    logic [2:0]   io_commits_info_3_instrSize;
    logic         io_commits_info_3_fpWen;
    logic         io_commits_info_3_rfWen;
    logic         io_commits_info_3_needFlush;
    logic [3:0]   io_commits_info_3_traceBlockInPipe_itype;
    logic [3:0]   io_commits_info_3_traceBlockInPipe_iretire;
    logic         io_commits_info_3_traceBlockInPipe_ilastsize;
    logic [49:0]  io_commits_info_3_debug_pc;
    logic [31:0]  io_commits_info_3_debug_instr;
    logic [5:0]   io_commits_info_3_debug_ldest;
    logic [7:0]   io_commits_info_3_debug_pdest;
    logic [7:0]   io_commits_info_3_debug_otherPdest_0;
    logic [7:0]   io_commits_info_3_debug_otherPdest_1;
    logic [7:0]   io_commits_info_3_debug_otherPdest_2;
    logic [7:0]   io_commits_info_3_debug_otherPdest_3;
    logic [7:0]   io_commits_info_3_debug_otherPdest_4;
    logic [7:0]   io_commits_info_3_debug_otherPdest_5;
    logic [7:0]   io_commits_info_3_debug_otherPdest_6;
    logic [34:0]  io_commits_info_3_debug_fuType;
    logic         io_commits_info_3_dirtyFs;
    logic         io_commits_info_3_dirtyVs;
    logic         io_commits_info_4_walk_v;
    logic         io_commits_info_4_commit_v;
    logic         io_commits_info_4_commit_w;
    logic [6:0]   io_commits_info_4_realDestSize;
    logic         io_commits_info_4_interrupt_safe;
    logic         io_commits_info_4_wflags;
    logic [4:0]   io_commits_info_4_fflags;
    logic         io_commits_info_4_vxsat;
    logic         io_commits_info_4_isRVC;
    logic         io_commits_info_4_isVset;
    logic         io_commits_info_4_isHls;
    logic         io_commits_info_4_isVls;
    logic         io_commits_info_4_vls;
    logic         io_commits_info_4_mmio;
    logic [2:0]   io_commits_info_4_commitType;
    logic         io_commits_info_4_ftqIdx_flag;
    logic [5:0]   io_commits_info_4_ftqIdx_value;
    logic [3:0]   io_commits_info_4_ftqOffset;
    logic [2:0]   io_commits_info_4_instrSize;
    logic         io_commits_info_4_fpWen;
    logic         io_commits_info_4_rfWen;
    logic         io_commits_info_4_needFlush;
    logic [3:0]   io_commits_info_4_traceBlockInPipe_itype;
    logic [3:0]   io_commits_info_4_traceBlockInPipe_iretire;
    logic         io_commits_info_4_traceBlockInPipe_ilastsize;
    logic [49:0]  io_commits_info_4_debug_pc;
    logic [31:0]  io_commits_info_4_debug_instr;
    logic [5:0]   io_commits_info_4_debug_ldest;
    logic [7:0]   io_commits_info_4_debug_pdest;
    logic [7:0]   io_commits_info_4_debug_otherPdest_0;
    logic [7:0]   io_commits_info_4_debug_otherPdest_1;
    logic [7:0]   io_commits_info_4_debug_otherPdest_2;
    logic [7:0]   io_commits_info_4_debug_otherPdest_3;
    logic [7:0]   io_commits_info_4_debug_otherPdest_4;
    logic [7:0]   io_commits_info_4_debug_otherPdest_5;
    logic [7:0]   io_commits_info_4_debug_otherPdest_6;
    logic [34:0]  io_commits_info_4_debug_fuType;
    logic         io_commits_info_4_dirtyFs;
    logic         io_commits_info_4_dirtyVs;
    logic         io_commits_info_5_walk_v;
    logic         io_commits_info_5_commit_v;
    logic         io_commits_info_5_commit_w;
    logic [6:0]   io_commits_info_5_realDestSize;
    logic         io_commits_info_5_interrupt_safe;
    logic         io_commits_info_5_wflags;
    logic [4:0]   io_commits_info_5_fflags;
    logic         io_commits_info_5_vxsat;
    logic         io_commits_info_5_isRVC;
    logic         io_commits_info_5_isVset;
    logic         io_commits_info_5_isHls;
    logic         io_commits_info_5_isVls;
    logic         io_commits_info_5_vls;
    logic         io_commits_info_5_mmio;
    logic [2:0]   io_commits_info_5_commitType;
    logic         io_commits_info_5_ftqIdx_flag;
    logic [5:0]   io_commits_info_5_ftqIdx_value;
    logic [3:0]   io_commits_info_5_ftqOffset;
    logic [2:0]   io_commits_info_5_instrSize;
    logic         io_commits_info_5_fpWen;
    logic         io_commits_info_5_rfWen;
    logic         io_commits_info_5_needFlush;
    logic [3:0]   io_commits_info_5_traceBlockInPipe_itype;
    logic [3:0]   io_commits_info_5_traceBlockInPipe_iretire;
    logic         io_commits_info_5_traceBlockInPipe_ilastsize;
    logic [49:0]  io_commits_info_5_debug_pc;
    logic [31:0]  io_commits_info_5_debug_instr;
    logic [5:0]   io_commits_info_5_debug_ldest;
    logic [7:0]   io_commits_info_5_debug_pdest;
    logic [7:0]   io_commits_info_5_debug_otherPdest_0;
    logic [7:0]   io_commits_info_5_debug_otherPdest_1;
    logic [7:0]   io_commits_info_5_debug_otherPdest_2;
    logic [7:0]   io_commits_info_5_debug_otherPdest_3;
    logic [7:0]   io_commits_info_5_debug_otherPdest_4;
    logic [7:0]   io_commits_info_5_debug_otherPdest_5;
    logic [7:0]   io_commits_info_5_debug_otherPdest_6;
    logic [34:0]  io_commits_info_5_debug_fuType;
    logic         io_commits_info_5_dirtyFs;
    logic         io_commits_info_5_dirtyVs;
    logic         io_commits_info_6_walk_v;
    logic         io_commits_info_6_commit_v;
    logic         io_commits_info_6_commit_w;
    logic [6:0]   io_commits_info_6_realDestSize;
    logic         io_commits_info_6_interrupt_safe;
    logic         io_commits_info_6_wflags;
    logic [4:0]   io_commits_info_6_fflags;
    logic         io_commits_info_6_vxsat;
    logic         io_commits_info_6_isRVC;
    logic         io_commits_info_6_isVset;
    logic         io_commits_info_6_isHls;
    logic         io_commits_info_6_isVls;
    logic         io_commits_info_6_vls;
    logic         io_commits_info_6_mmio;
    logic [2:0]   io_commits_info_6_commitType;
    logic         io_commits_info_6_ftqIdx_flag;
    logic [5:0]   io_commits_info_6_ftqIdx_value;
    logic [3:0]   io_commits_info_6_ftqOffset;
    logic [2:0]   io_commits_info_6_instrSize;
    logic         io_commits_info_6_fpWen;
    logic         io_commits_info_6_rfWen;
    logic         io_commits_info_6_needFlush;
    logic [3:0]   io_commits_info_6_traceBlockInPipe_itype;
    logic [3:0]   io_commits_info_6_traceBlockInPipe_iretire;
    logic         io_commits_info_6_traceBlockInPipe_ilastsize;
    logic [49:0]  io_commits_info_6_debug_pc;
    logic [31:0]  io_commits_info_6_debug_instr;
    logic [5:0]   io_commits_info_6_debug_ldest;
    logic [7:0]   io_commits_info_6_debug_pdest;
    logic [7:0]   io_commits_info_6_debug_otherPdest_0;
    logic [7:0]   io_commits_info_6_debug_otherPdest_1;
    logic [7:0]   io_commits_info_6_debug_otherPdest_2;
    logic [7:0]   io_commits_info_6_debug_otherPdest_3;
    logic [7:0]   io_commits_info_6_debug_otherPdest_4;
    logic [7:0]   io_commits_info_6_debug_otherPdest_5;
    logic [7:0]   io_commits_info_6_debug_otherPdest_6;
    logic [34:0]  io_commits_info_6_debug_fuType;
    logic         io_commits_info_6_dirtyFs;
    logic         io_commits_info_6_dirtyVs;
    logic         io_commits_info_7_walk_v;
    logic         io_commits_info_7_commit_v;
    logic         io_commits_info_7_commit_w;
    logic [6:0]   io_commits_info_7_realDestSize;
    logic         io_commits_info_7_interrupt_safe;
    logic         io_commits_info_7_wflags;
    logic [4:0]   io_commits_info_7_fflags;
    logic         io_commits_info_7_vxsat;
    logic         io_commits_info_7_isRVC;
    logic         io_commits_info_7_isVset;
    logic         io_commits_info_7_isHls;
    logic         io_commits_info_7_isVls;
    logic         io_commits_info_7_vls;
    logic         io_commits_info_7_mmio;
    logic [2:0]   io_commits_info_7_commitType;
    logic         io_commits_info_7_ftqIdx_flag;
    logic [5:0]   io_commits_info_7_ftqIdx_value;
    logic [3:0]   io_commits_info_7_ftqOffset;
    logic [2:0]   io_commits_info_7_instrSize;
    logic         io_commits_info_7_fpWen;
    logic         io_commits_info_7_rfWen;
    logic         io_commits_info_7_needFlush;
    logic [3:0]   io_commits_info_7_traceBlockInPipe_itype;
    logic [3:0]   io_commits_info_7_traceBlockInPipe_iretire;
    logic         io_commits_info_7_traceBlockInPipe_ilastsize;
    logic [49:0]  io_commits_info_7_debug_pc;
    logic [31:0]  io_commits_info_7_debug_instr;
    logic [5:0]   io_commits_info_7_debug_ldest;
    logic [7:0]   io_commits_info_7_debug_pdest;
    logic [7:0]   io_commits_info_7_debug_otherPdest_0;
    logic [7:0]   io_commits_info_7_debug_otherPdest_1;
    logic [7:0]   io_commits_info_7_debug_otherPdest_2;
    logic [7:0]   io_commits_info_7_debug_otherPdest_3;
    logic [7:0]   io_commits_info_7_debug_otherPdest_4;
    logic [7:0]   io_commits_info_7_debug_otherPdest_5;
    logic [7:0]   io_commits_info_7_debug_otherPdest_6;
    logic [34:0]  io_commits_info_7_debug_fuType;
    logic         io_commits_info_7_dirtyFs;
    logic         io_commits_info_7_dirtyVs;
    logic         io_commits_robIdx_0_flag;
    logic [7:0]   io_commits_robIdx_0_value;
    logic         io_commits_robIdx_1_flag;
    logic [7:0]   io_commits_robIdx_1_value;
    logic         io_commits_robIdx_2_flag;
    logic [7:0]   io_commits_robIdx_2_value;
    logic         io_commits_robIdx_3_flag;
    logic [7:0]   io_commits_robIdx_3_value;
    logic         io_commits_robIdx_4_flag;
    logic [7:0]   io_commits_robIdx_4_value;
    logic         io_commits_robIdx_5_flag;
    logic [7:0]   io_commits_robIdx_5_value;
    logic         io_commits_robIdx_6_flag;
    logic [7:0]   io_commits_robIdx_6_value;
    logic         io_commits_robIdx_7_flag;
    logic [7:0]   io_commits_robIdx_7_value;
    logic         io_trace_blockCommit ;
    logic         io_trace_traceCommitInfo_blocks_0_valid;
    logic [5:0]   io_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value;
    logic [3:0]   io_trace_traceCommitInfo_blocks_0_bits_ftqOffset;
    logic [3:0]   io_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype;
    logic [3:0]   io_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire;
    logic         io_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize;
    logic         io_trace_traceCommitInfo_blocks_1_valid;
    logic [5:0]   io_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value;
    logic [3:0]   io_trace_traceCommitInfo_blocks_1_bits_ftqOffset;
    logic [3:0]   io_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype;
    logic [3:0]   io_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire;
    logic         io_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize;
    logic         io_trace_traceCommitInfo_blocks_2_valid;
    logic [5:0]   io_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value;
    logic [3:0]   io_trace_traceCommitInfo_blocks_2_bits_ftqOffset;
    logic [3:0]   io_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype;
    logic [3:0]   io_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire;
    logic         io_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize;
    logic         io_trace_traceCommitInfo_blocks_3_valid;
    logic [5:0]   io_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value;
    logic [3:0]   io_trace_traceCommitInfo_blocks_3_bits_ftqOffset;
    logic [3:0]   io_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype;
    logic [3:0]   io_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire;
    logic         io_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize;
    logic         io_trace_traceCommitInfo_blocks_4_valid;
    logic [5:0]   io_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value;
    logic [3:0]   io_trace_traceCommitInfo_blocks_4_bits_ftqOffset;
    logic [3:0]   io_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype;
    logic [3:0]   io_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire;
    logic         io_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize;
    logic         io_trace_traceCommitInfo_blocks_5_valid;
    logic [5:0]   io_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value;
    logic [3:0]   io_trace_traceCommitInfo_blocks_5_bits_ftqOffset;
    logic [3:0]   io_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype;
    logic [3:0]   io_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire;
    logic         io_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize;
    logic         io_trace_traceCommitInfo_blocks_6_valid;
    logic [5:0]   io_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value;
    logic [3:0]   io_trace_traceCommitInfo_blocks_6_bits_ftqOffset;
    logic [3:0]   io_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype;
    logic [3:0]   io_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire;
    logic         io_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize;
    logic         io_trace_traceCommitInfo_blocks_7_valid;
    logic [5:0]   io_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value;
    logic [3:0]   io_trace_traceCommitInfo_blocks_7_bits_ftqOffset;
    logic [3:0]   io_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype;
    logic [3:0]   io_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire;
    logic         io_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize;
    logic         io_rabCommits_isCommit;
    logic         io_rabCommits_commitValid_0;
    logic         io_rabCommits_commitValid_1;
    logic         io_rabCommits_commitValid_2;
    logic         io_rabCommits_commitValid_3;
    logic         io_rabCommits_commitValid_4;
    logic         io_rabCommits_commitValid_5;
    logic         io_rabCommits_isWalk ;
    logic         io_rabCommits_walkValid_0;
    logic         io_rabCommits_walkValid_1;
    logic         io_rabCommits_walkValid_2;
    logic         io_rabCommits_walkValid_3;
    logic         io_rabCommits_walkValid_4;
    logic         io_rabCommits_walkValid_5;
    logic [5:0]   io_rabCommits_info_0_ldest;
    logic [7:0]   io_rabCommits_info_0_pdest;
    logic         io_rabCommits_info_0_rfWen;
    logic         io_rabCommits_info_0_fpWen;
    logic         io_rabCommits_info_0_vecWen;
    logic         io_rabCommits_info_0_v0Wen;
    logic         io_rabCommits_info_0_vlWen;
    logic         io_rabCommits_info_0_isMove;
    logic [5:0]   io_rabCommits_info_1_ldest;
    logic [7:0]   io_rabCommits_info_1_pdest;
    logic         io_rabCommits_info_1_rfWen;
    logic         io_rabCommits_info_1_fpWen;
    logic         io_rabCommits_info_1_vecWen;
    logic         io_rabCommits_info_1_v0Wen;
    logic         io_rabCommits_info_1_vlWen;
    logic         io_rabCommits_info_1_isMove;
    logic [5:0]   io_rabCommits_info_2_ldest;
    logic [7:0]   io_rabCommits_info_2_pdest;
    logic         io_rabCommits_info_2_rfWen;
    logic         io_rabCommits_info_2_fpWen;
    logic         io_rabCommits_info_2_vecWen;
    logic         io_rabCommits_info_2_v0Wen;
    logic         io_rabCommits_info_2_vlWen;
    logic         io_rabCommits_info_2_isMove;
    logic [5:0]   io_rabCommits_info_3_ldest;
    logic [7:0]   io_rabCommits_info_3_pdest;
    logic         io_rabCommits_info_3_rfWen;
    logic         io_rabCommits_info_3_fpWen;
    logic         io_rabCommits_info_3_vecWen;
    logic         io_rabCommits_info_3_v0Wen;
    logic         io_rabCommits_info_3_vlWen;
    logic         io_rabCommits_info_3_isMove;
    logic [5:0]   io_rabCommits_info_4_ldest;
    logic [7:0]   io_rabCommits_info_4_pdest;
    logic         io_rabCommits_info_4_rfWen;
    logic         io_rabCommits_info_4_fpWen;
    logic         io_rabCommits_info_4_vecWen;
    logic         io_rabCommits_info_4_v0Wen;
    logic         io_rabCommits_info_4_vlWen;
    logic         io_rabCommits_info_4_isMove;
    logic [5:0]   io_rabCommits_info_5_ldest;
    logic [7:0]   io_rabCommits_info_5_pdest;
    logic         io_rabCommits_info_5_rfWen;
    logic         io_rabCommits_info_5_fpWen;
    logic         io_rabCommits_info_5_vecWen;
    logic         io_rabCommits_info_5_v0Wen;
    logic         io_rabCommits_info_5_vlWen;
    logic         io_rabCommits_info_5_isMove;
    logic         io_diffCommits_commitValid_0;
    logic         io_diffCommits_commitValid_1;
    logic         io_diffCommits_commitValid_2;
    logic         io_diffCommits_commitValid_3;
    logic         io_diffCommits_commitValid_4;
    logic         io_diffCommits_commitValid_5;
    logic         io_diffCommits_commitValid_6;
    logic         io_diffCommits_commitValid_7;
    logic         io_diffCommits_commitValid_8;
    logic         io_diffCommits_commitValid_9;
    logic         io_diffCommits_commitValid_10;
    logic         io_diffCommits_commitValid_11;
    logic         io_diffCommits_commitValid_12;
    logic         io_diffCommits_commitValid_13;
    logic         io_diffCommits_commitValid_14;
    logic         io_diffCommits_commitValid_15;
    logic         io_diffCommits_commitValid_16;
    logic         io_diffCommits_commitValid_17;
    logic         io_diffCommits_commitValid_18;
    logic         io_diffCommits_commitValid_19;
    logic         io_diffCommits_commitValid_20;
    logic         io_diffCommits_commitValid_21;
    logic         io_diffCommits_commitValid_22;
    logic         io_diffCommits_commitValid_23;
    logic         io_diffCommits_commitValid_24;
    logic         io_diffCommits_commitValid_25;
    logic         io_diffCommits_commitValid_26;
    logic         io_diffCommits_commitValid_27;
    logic         io_diffCommits_commitValid_28;
    logic         io_diffCommits_commitValid_29;
    logic         io_diffCommits_commitValid_30;
    logic         io_diffCommits_commitValid_31;
    logic         io_diffCommits_commitValid_32;
    logic         io_diffCommits_commitValid_33;
    logic         io_diffCommits_commitValid_34;
    logic         io_diffCommits_commitValid_35;
    logic         io_diffCommits_commitValid_36;
    logic         io_diffCommits_commitValid_37;
    logic         io_diffCommits_commitValid_38;
    logic         io_diffCommits_commitValid_39;
    logic         io_diffCommits_commitValid_40;
    logic         io_diffCommits_commitValid_41;
    logic         io_diffCommits_commitValid_42;
    logic         io_diffCommits_commitValid_43;
    logic         io_diffCommits_commitValid_44;
    logic         io_diffCommits_commitValid_45;
    logic         io_diffCommits_commitValid_46;
    logic         io_diffCommits_commitValid_47;
    logic         io_diffCommits_commitValid_48;
    logic         io_diffCommits_commitValid_49;
    logic         io_diffCommits_commitValid_50;
    logic         io_diffCommits_commitValid_51;
    logic         io_diffCommits_commitValid_52;
    logic         io_diffCommits_commitValid_53;
    logic         io_diffCommits_commitValid_54;
    logic         io_diffCommits_commitValid_55;
    logic         io_diffCommits_commitValid_56;
    logic         io_diffCommits_commitValid_57;
    logic         io_diffCommits_commitValid_58;
    logic         io_diffCommits_commitValid_59;
    logic         io_diffCommits_commitValid_60;
    logic         io_diffCommits_commitValid_61;
    logic         io_diffCommits_commitValid_62;
    logic         io_diffCommits_commitValid_63;
    logic         io_diffCommits_commitValid_64;
    logic         io_diffCommits_commitValid_65;
    logic         io_diffCommits_commitValid_66;
    logic         io_diffCommits_commitValid_67;
    logic         io_diffCommits_commitValid_68;
    logic         io_diffCommits_commitValid_69;
    logic         io_diffCommits_commitValid_70;
    logic         io_diffCommits_commitValid_71;
    logic         io_diffCommits_commitValid_72;
    logic         io_diffCommits_commitValid_73;
    logic         io_diffCommits_commitValid_74;
    logic         io_diffCommits_commitValid_75;
    logic         io_diffCommits_commitValid_76;
    logic         io_diffCommits_commitValid_77;
    logic         io_diffCommits_commitValid_78;
    logic         io_diffCommits_commitValid_79;
    logic         io_diffCommits_commitValid_80;
    logic         io_diffCommits_commitValid_81;
    logic         io_diffCommits_commitValid_82;
    logic         io_diffCommits_commitValid_83;
    logic         io_diffCommits_commitValid_84;
    logic         io_diffCommits_commitValid_85;
    logic         io_diffCommits_commitValid_86;
    logic         io_diffCommits_commitValid_87;
    logic         io_diffCommits_commitValid_88;
    logic         io_diffCommits_commitValid_89;
    logic         io_diffCommits_commitValid_90;
    logic         io_diffCommits_commitValid_91;
    logic         io_diffCommits_commitValid_92;
    logic         io_diffCommits_commitValid_93;
    logic         io_diffCommits_commitValid_94;
    logic         io_diffCommits_commitValid_95;
    logic         io_diffCommits_commitValid_96;
    logic         io_diffCommits_commitValid_97;
    logic         io_diffCommits_commitValid_98;
    logic         io_diffCommits_commitValid_99;
    logic         io_diffCommits_commitValid_100;
    logic         io_diffCommits_commitValid_101;
    logic         io_diffCommits_commitValid_102;
    logic         io_diffCommits_commitValid_103;
    logic         io_diffCommits_commitValid_104;
    logic         io_diffCommits_commitValid_105;
    logic         io_diffCommits_commitValid_106;
    logic         io_diffCommits_commitValid_107;
    logic         io_diffCommits_commitValid_108;
    logic         io_diffCommits_commitValid_109;
    logic         io_diffCommits_commitValid_110;
    logic         io_diffCommits_commitValid_111;
    logic         io_diffCommits_commitValid_112;
    logic         io_diffCommits_commitValid_113;
    logic         io_diffCommits_commitValid_114;
    logic         io_diffCommits_commitValid_115;
    logic         io_diffCommits_commitValid_116;
    logic         io_diffCommits_commitValid_117;
    logic         io_diffCommits_commitValid_118;
    logic         io_diffCommits_commitValid_119;
    logic         io_diffCommits_commitValid_120;
    logic         io_diffCommits_commitValid_121;
    logic         io_diffCommits_commitValid_122;
    logic         io_diffCommits_commitValid_123;
    logic         io_diffCommits_commitValid_124;
    logic         io_diffCommits_commitValid_125;
    logic         io_diffCommits_commitValid_126;
    logic         io_diffCommits_commitValid_127;
    logic         io_diffCommits_commitValid_128;
    logic         io_diffCommits_commitValid_129;
    logic         io_diffCommits_commitValid_130;
    logic         io_diffCommits_commitValid_131;
    logic         io_diffCommits_commitValid_132;
    logic         io_diffCommits_commitValid_133;
    logic         io_diffCommits_commitValid_134;
    logic         io_diffCommits_commitValid_135;
    logic         io_diffCommits_commitValid_136;
    logic         io_diffCommits_commitValid_137;
    logic         io_diffCommits_commitValid_138;
    logic         io_diffCommits_commitValid_139;
    logic         io_diffCommits_commitValid_140;
    logic         io_diffCommits_commitValid_141;
    logic         io_diffCommits_commitValid_142;
    logic         io_diffCommits_commitValid_143;
    logic         io_diffCommits_commitValid_144;
    logic         io_diffCommits_commitValid_145;
    logic         io_diffCommits_commitValid_146;
    logic         io_diffCommits_commitValid_147;
    logic         io_diffCommits_commitValid_148;
    logic         io_diffCommits_commitValid_149;
    logic         io_diffCommits_commitValid_150;
    logic         io_diffCommits_commitValid_151;
    logic         io_diffCommits_commitValid_152;
    logic         io_diffCommits_commitValid_153;
    logic         io_diffCommits_commitValid_154;
    logic         io_diffCommits_commitValid_155;
    logic         io_diffCommits_commitValid_156;
    logic         io_diffCommits_commitValid_157;
    logic         io_diffCommits_commitValid_158;
    logic         io_diffCommits_commitValid_159;
    logic         io_diffCommits_commitValid_160;
    logic         io_diffCommits_commitValid_161;
    logic         io_diffCommits_commitValid_162;
    logic         io_diffCommits_commitValid_163;
    logic         io_diffCommits_commitValid_164;
    logic         io_diffCommits_commitValid_165;
    logic         io_diffCommits_commitValid_166;
    logic         io_diffCommits_commitValid_167;
    logic         io_diffCommits_commitValid_168;
    logic         io_diffCommits_commitValid_169;
    logic         io_diffCommits_commitValid_170;
    logic         io_diffCommits_commitValid_171;
    logic         io_diffCommits_commitValid_172;
    logic         io_diffCommits_commitValid_173;
    logic         io_diffCommits_commitValid_174;
    logic         io_diffCommits_commitValid_175;
    logic         io_diffCommits_commitValid_176;
    logic         io_diffCommits_commitValid_177;
    logic         io_diffCommits_commitValid_178;
    logic         io_diffCommits_commitValid_179;
    logic         io_diffCommits_commitValid_180;
    logic         io_diffCommits_commitValid_181;
    logic         io_diffCommits_commitValid_182;
    logic         io_diffCommits_commitValid_183;
    logic         io_diffCommits_commitValid_184;
    logic         io_diffCommits_commitValid_185;
    logic         io_diffCommits_commitValid_186;
    logic         io_diffCommits_commitValid_187;
    logic         io_diffCommits_commitValid_188;
    logic         io_diffCommits_commitValid_189;
    logic         io_diffCommits_commitValid_190;
    logic         io_diffCommits_commitValid_191;
    logic         io_diffCommits_commitValid_192;
    logic         io_diffCommits_commitValid_193;
    logic         io_diffCommits_commitValid_194;
    logic         io_diffCommits_commitValid_195;
    logic         io_diffCommits_commitValid_196;
    logic         io_diffCommits_commitValid_197;
    logic         io_diffCommits_commitValid_198;
    logic         io_diffCommits_commitValid_199;
    logic         io_diffCommits_commitValid_200;
    logic         io_diffCommits_commitValid_201;
    logic         io_diffCommits_commitValid_202;
    logic         io_diffCommits_commitValid_203;
    logic         io_diffCommits_commitValid_204;
    logic         io_diffCommits_commitValid_205;
    logic         io_diffCommits_commitValid_206;
    logic         io_diffCommits_commitValid_207;
    logic         io_diffCommits_commitValid_208;
    logic         io_diffCommits_commitValid_209;
    logic         io_diffCommits_commitValid_210;
    logic         io_diffCommits_commitValid_211;
    logic         io_diffCommits_commitValid_212;
    logic         io_diffCommits_commitValid_213;
    logic         io_diffCommits_commitValid_214;
    logic         io_diffCommits_commitValid_215;
    logic         io_diffCommits_commitValid_216;
    logic         io_diffCommits_commitValid_217;
    logic         io_diffCommits_commitValid_218;
    logic         io_diffCommits_commitValid_219;
    logic         io_diffCommits_commitValid_220;
    logic         io_diffCommits_commitValid_221;
    logic         io_diffCommits_commitValid_222;
    logic         io_diffCommits_commitValid_223;
    logic         io_diffCommits_commitValid_224;
    logic         io_diffCommits_commitValid_225;
    logic         io_diffCommits_commitValid_226;
    logic         io_diffCommits_commitValid_227;
    logic         io_diffCommits_commitValid_228;
    logic         io_diffCommits_commitValid_229;
    logic         io_diffCommits_commitValid_230;
    logic         io_diffCommits_commitValid_231;
    logic         io_diffCommits_commitValid_232;
    logic         io_diffCommits_commitValid_233;
    logic         io_diffCommits_commitValid_234;
    logic         io_diffCommits_commitValid_235;
    logic         io_diffCommits_commitValid_236;
    logic         io_diffCommits_commitValid_237;
    logic         io_diffCommits_commitValid_238;
    logic         io_diffCommits_commitValid_239;
    logic         io_diffCommits_commitValid_240;
    logic         io_diffCommits_commitValid_241;
    logic         io_diffCommits_commitValid_242;
    logic         io_diffCommits_commitValid_243;
    logic         io_diffCommits_commitValid_244;
    logic         io_diffCommits_commitValid_245;
    logic         io_diffCommits_commitValid_246;
    logic         io_diffCommits_commitValid_247;
    logic         io_diffCommits_commitValid_248;
    logic         io_diffCommits_commitValid_249;
    logic         io_diffCommits_commitValid_250;
    logic         io_diffCommits_commitValid_251;
    logic         io_diffCommits_commitValid_252;
    logic         io_diffCommits_commitValid_253;
    logic         io_diffCommits_commitValid_254;
    logic [5:0]   io_diffCommits_info_0_ldest;
    logic [7:0]   io_diffCommits_info_0_pdest;
    logic         io_diffCommits_info_0_rfWen;
    logic         io_diffCommits_info_0_fpWen;
    logic         io_diffCommits_info_0_vecWen;
    logic         io_diffCommits_info_0_v0Wen;
    logic         io_diffCommits_info_0_vlWen;
    logic [5:0]   io_diffCommits_info_1_ldest;
    logic [7:0]   io_diffCommits_info_1_pdest;
    logic         io_diffCommits_info_1_rfWen;
    logic         io_diffCommits_info_1_fpWen;
    logic         io_diffCommits_info_1_vecWen;
    logic         io_diffCommits_info_1_v0Wen;
    logic         io_diffCommits_info_1_vlWen;
    logic [5:0]   io_diffCommits_info_2_ldest;
    logic [7:0]   io_diffCommits_info_2_pdest;
    logic         io_diffCommits_info_2_rfWen;
    logic         io_diffCommits_info_2_fpWen;
    logic         io_diffCommits_info_2_vecWen;
    logic         io_diffCommits_info_2_v0Wen;
    logic         io_diffCommits_info_2_vlWen;
    logic [5:0]   io_diffCommits_info_3_ldest;
    logic [7:0]   io_diffCommits_info_3_pdest;
    logic         io_diffCommits_info_3_rfWen;
    logic         io_diffCommits_info_3_fpWen;
    logic         io_diffCommits_info_3_vecWen;
    logic         io_diffCommits_info_3_v0Wen;
    logic         io_diffCommits_info_3_vlWen;
    logic [5:0]   io_diffCommits_info_4_ldest;
    logic [7:0]   io_diffCommits_info_4_pdest;
    logic         io_diffCommits_info_4_rfWen;
    logic         io_diffCommits_info_4_fpWen;
    logic         io_diffCommits_info_4_vecWen;
    logic         io_diffCommits_info_4_v0Wen;
    logic         io_diffCommits_info_4_vlWen;
    logic [5:0]   io_diffCommits_info_5_ldest;
    logic [7:0]   io_diffCommits_info_5_pdest;
    logic         io_diffCommits_info_5_rfWen;
    logic         io_diffCommits_info_5_fpWen;
    logic         io_diffCommits_info_5_vecWen;
    logic         io_diffCommits_info_5_v0Wen;
    logic         io_diffCommits_info_5_vlWen;
    logic [5:0]   io_diffCommits_info_6_ldest;
    logic [7:0]   io_diffCommits_info_6_pdest;
    logic         io_diffCommits_info_6_rfWen;
    logic         io_diffCommits_info_6_fpWen;
    logic         io_diffCommits_info_6_vecWen;
    logic         io_diffCommits_info_6_v0Wen;
    logic         io_diffCommits_info_6_vlWen;
    logic [5:0]   io_diffCommits_info_7_ldest;
    logic [7:0]   io_diffCommits_info_7_pdest;
    logic         io_diffCommits_info_7_rfWen;
    logic         io_diffCommits_info_7_fpWen;
    logic         io_diffCommits_info_7_vecWen;
    logic         io_diffCommits_info_7_v0Wen;
    logic         io_diffCommits_info_7_vlWen;
    logic [5:0]   io_diffCommits_info_8_ldest;
    logic [7:0]   io_diffCommits_info_8_pdest;
    logic         io_diffCommits_info_8_rfWen;
    logic         io_diffCommits_info_8_fpWen;
    logic         io_diffCommits_info_8_vecWen;
    logic         io_diffCommits_info_8_v0Wen;
    logic         io_diffCommits_info_8_vlWen;
    logic [5:0]   io_diffCommits_info_9_ldest;
    logic [7:0]   io_diffCommits_info_9_pdest;
    logic         io_diffCommits_info_9_rfWen;
    logic         io_diffCommits_info_9_fpWen;
    logic         io_diffCommits_info_9_vecWen;
    logic         io_diffCommits_info_9_v0Wen;
    logic         io_diffCommits_info_9_vlWen;
    logic [5:0]   io_diffCommits_info_10_ldest;
    logic [7:0]   io_diffCommits_info_10_pdest;
    logic         io_diffCommits_info_10_rfWen;
    logic         io_diffCommits_info_10_fpWen;
    logic         io_diffCommits_info_10_vecWen;
    logic         io_diffCommits_info_10_v0Wen;
    logic         io_diffCommits_info_10_vlWen;
    logic [5:0]   io_diffCommits_info_11_ldest;
    logic [7:0]   io_diffCommits_info_11_pdest;
    logic         io_diffCommits_info_11_rfWen;
    logic         io_diffCommits_info_11_fpWen;
    logic         io_diffCommits_info_11_vecWen;
    logic         io_diffCommits_info_11_v0Wen;
    logic         io_diffCommits_info_11_vlWen;
    logic [5:0]   io_diffCommits_info_12_ldest;
    logic [7:0]   io_diffCommits_info_12_pdest;
    logic         io_diffCommits_info_12_rfWen;
    logic         io_diffCommits_info_12_fpWen;
    logic         io_diffCommits_info_12_vecWen;
    logic         io_diffCommits_info_12_v0Wen;
    logic         io_diffCommits_info_12_vlWen;
    logic [5:0]   io_diffCommits_info_13_ldest;
    logic [7:0]   io_diffCommits_info_13_pdest;
    logic         io_diffCommits_info_13_rfWen;
    logic         io_diffCommits_info_13_fpWen;
    logic         io_diffCommits_info_13_vecWen;
    logic         io_diffCommits_info_13_v0Wen;
    logic         io_diffCommits_info_13_vlWen;
    logic [5:0]   io_diffCommits_info_14_ldest;
    logic [7:0]   io_diffCommits_info_14_pdest;
    logic         io_diffCommits_info_14_rfWen;
    logic         io_diffCommits_info_14_fpWen;
    logic         io_diffCommits_info_14_vecWen;
    logic         io_diffCommits_info_14_v0Wen;
    logic         io_diffCommits_info_14_vlWen;
    logic [5:0]   io_diffCommits_info_15_ldest;
    logic [7:0]   io_diffCommits_info_15_pdest;
    logic         io_diffCommits_info_15_rfWen;
    logic         io_diffCommits_info_15_fpWen;
    logic         io_diffCommits_info_15_vecWen;
    logic         io_diffCommits_info_15_v0Wen;
    logic         io_diffCommits_info_15_vlWen;
    logic [5:0]   io_diffCommits_info_16_ldest;
    logic [7:0]   io_diffCommits_info_16_pdest;
    logic         io_diffCommits_info_16_rfWen;
    logic         io_diffCommits_info_16_fpWen;
    logic         io_diffCommits_info_16_vecWen;
    logic         io_diffCommits_info_16_v0Wen;
    logic         io_diffCommits_info_16_vlWen;
    logic [5:0]   io_diffCommits_info_17_ldest;
    logic [7:0]   io_diffCommits_info_17_pdest;
    logic         io_diffCommits_info_17_rfWen;
    logic         io_diffCommits_info_17_fpWen;
    logic         io_diffCommits_info_17_vecWen;
    logic         io_diffCommits_info_17_v0Wen;
    logic         io_diffCommits_info_17_vlWen;
    logic [5:0]   io_diffCommits_info_18_ldest;
    logic [7:0]   io_diffCommits_info_18_pdest;
    logic         io_diffCommits_info_18_rfWen;
    logic         io_diffCommits_info_18_fpWen;
    logic         io_diffCommits_info_18_vecWen;
    logic         io_diffCommits_info_18_v0Wen;
    logic         io_diffCommits_info_18_vlWen;
    logic [5:0]   io_diffCommits_info_19_ldest;
    logic [7:0]   io_diffCommits_info_19_pdest;
    logic         io_diffCommits_info_19_rfWen;
    logic         io_diffCommits_info_19_fpWen;
    logic         io_diffCommits_info_19_vecWen;
    logic         io_diffCommits_info_19_v0Wen;
    logic         io_diffCommits_info_19_vlWen;
    logic [5:0]   io_diffCommits_info_20_ldest;
    logic [7:0]   io_diffCommits_info_20_pdest;
    logic         io_diffCommits_info_20_rfWen;
    logic         io_diffCommits_info_20_fpWen;
    logic         io_diffCommits_info_20_vecWen;
    logic         io_diffCommits_info_20_v0Wen;
    logic         io_diffCommits_info_20_vlWen;
    logic [5:0]   io_diffCommits_info_21_ldest;
    logic [7:0]   io_diffCommits_info_21_pdest;
    logic         io_diffCommits_info_21_rfWen;
    logic         io_diffCommits_info_21_fpWen;
    logic         io_diffCommits_info_21_vecWen;
    logic         io_diffCommits_info_21_v0Wen;
    logic         io_diffCommits_info_21_vlWen;
    logic [5:0]   io_diffCommits_info_22_ldest;
    logic [7:0]   io_diffCommits_info_22_pdest;
    logic         io_diffCommits_info_22_rfWen;
    logic         io_diffCommits_info_22_fpWen;
    logic         io_diffCommits_info_22_vecWen;
    logic         io_diffCommits_info_22_v0Wen;
    logic         io_diffCommits_info_22_vlWen;
    logic [5:0]   io_diffCommits_info_23_ldest;
    logic [7:0]   io_diffCommits_info_23_pdest;
    logic         io_diffCommits_info_23_rfWen;
    logic         io_diffCommits_info_23_fpWen;
    logic         io_diffCommits_info_23_vecWen;
    logic         io_diffCommits_info_23_v0Wen;
    logic         io_diffCommits_info_23_vlWen;
    logic [5:0]   io_diffCommits_info_24_ldest;
    logic [7:0]   io_diffCommits_info_24_pdest;
    logic         io_diffCommits_info_24_rfWen;
    logic         io_diffCommits_info_24_fpWen;
    logic         io_diffCommits_info_24_vecWen;
    logic         io_diffCommits_info_24_v0Wen;
    logic         io_diffCommits_info_24_vlWen;
    logic [5:0]   io_diffCommits_info_25_ldest;
    logic [7:0]   io_diffCommits_info_25_pdest;
    logic         io_diffCommits_info_25_rfWen;
    logic         io_diffCommits_info_25_fpWen;
    logic         io_diffCommits_info_25_vecWen;
    logic         io_diffCommits_info_25_v0Wen;
    logic         io_diffCommits_info_25_vlWen;
    logic [5:0]   io_diffCommits_info_26_ldest;
    logic [7:0]   io_diffCommits_info_26_pdest;
    logic         io_diffCommits_info_26_rfWen;
    logic         io_diffCommits_info_26_fpWen;
    logic         io_diffCommits_info_26_vecWen;
    logic         io_diffCommits_info_26_v0Wen;
    logic         io_diffCommits_info_26_vlWen;
    logic [5:0]   io_diffCommits_info_27_ldest;
    logic [7:0]   io_diffCommits_info_27_pdest;
    logic         io_diffCommits_info_27_rfWen;
    logic         io_diffCommits_info_27_fpWen;
    logic         io_diffCommits_info_27_vecWen;
    logic         io_diffCommits_info_27_v0Wen;
    logic         io_diffCommits_info_27_vlWen;
    logic [5:0]   io_diffCommits_info_28_ldest;
    logic [7:0]   io_diffCommits_info_28_pdest;
    logic         io_diffCommits_info_28_rfWen;
    logic         io_diffCommits_info_28_fpWen;
    logic         io_diffCommits_info_28_vecWen;
    logic         io_diffCommits_info_28_v0Wen;
    logic         io_diffCommits_info_28_vlWen;
    logic [5:0]   io_diffCommits_info_29_ldest;
    logic [7:0]   io_diffCommits_info_29_pdest;
    logic         io_diffCommits_info_29_rfWen;
    logic         io_diffCommits_info_29_fpWen;
    logic         io_diffCommits_info_29_vecWen;
    logic         io_diffCommits_info_29_v0Wen;
    logic         io_diffCommits_info_29_vlWen;
    logic [5:0]   io_diffCommits_info_30_ldest;
    logic [7:0]   io_diffCommits_info_30_pdest;
    logic         io_diffCommits_info_30_rfWen;
    logic         io_diffCommits_info_30_fpWen;
    logic         io_diffCommits_info_30_vecWen;
    logic         io_diffCommits_info_30_v0Wen;
    logic         io_diffCommits_info_30_vlWen;
    logic [5:0]   io_diffCommits_info_31_ldest;
    logic [7:0]   io_diffCommits_info_31_pdest;
    logic         io_diffCommits_info_31_rfWen;
    logic         io_diffCommits_info_31_fpWen;
    logic         io_diffCommits_info_31_vecWen;
    logic         io_diffCommits_info_31_v0Wen;
    logic         io_diffCommits_info_31_vlWen;
    logic [5:0]   io_diffCommits_info_32_ldest;
    logic [7:0]   io_diffCommits_info_32_pdest;
    logic         io_diffCommits_info_32_rfWen;
    logic         io_diffCommits_info_32_fpWen;
    logic         io_diffCommits_info_32_vecWen;
    logic         io_diffCommits_info_32_v0Wen;
    logic         io_diffCommits_info_32_vlWen;
    logic [5:0]   io_diffCommits_info_33_ldest;
    logic [7:0]   io_diffCommits_info_33_pdest;
    logic         io_diffCommits_info_33_rfWen;
    logic         io_diffCommits_info_33_fpWen;
    logic         io_diffCommits_info_33_vecWen;
    logic         io_diffCommits_info_33_v0Wen;
    logic         io_diffCommits_info_33_vlWen;
    logic [5:0]   io_diffCommits_info_34_ldest;
    logic [7:0]   io_diffCommits_info_34_pdest;
    logic         io_diffCommits_info_34_rfWen;
    logic         io_diffCommits_info_34_fpWen;
    logic         io_diffCommits_info_34_vecWen;
    logic         io_diffCommits_info_34_v0Wen;
    logic         io_diffCommits_info_34_vlWen;
    logic [5:0]   io_diffCommits_info_35_ldest;
    logic [7:0]   io_diffCommits_info_35_pdest;
    logic         io_diffCommits_info_35_rfWen;
    logic         io_diffCommits_info_35_fpWen;
    logic         io_diffCommits_info_35_vecWen;
    logic         io_diffCommits_info_35_v0Wen;
    logic         io_diffCommits_info_35_vlWen;
    logic [5:0]   io_diffCommits_info_36_ldest;
    logic [7:0]   io_diffCommits_info_36_pdest;
    logic         io_diffCommits_info_36_rfWen;
    logic         io_diffCommits_info_36_fpWen;
    logic         io_diffCommits_info_36_vecWen;
    logic         io_diffCommits_info_36_v0Wen;
    logic         io_diffCommits_info_36_vlWen;
    logic [5:0]   io_diffCommits_info_37_ldest;
    logic [7:0]   io_diffCommits_info_37_pdest;
    logic         io_diffCommits_info_37_rfWen;
    logic         io_diffCommits_info_37_fpWen;
    logic         io_diffCommits_info_37_vecWen;
    logic         io_diffCommits_info_37_v0Wen;
    logic         io_diffCommits_info_37_vlWen;
    logic [5:0]   io_diffCommits_info_38_ldest;
    logic [7:0]   io_diffCommits_info_38_pdest;
    logic         io_diffCommits_info_38_rfWen;
    logic         io_diffCommits_info_38_fpWen;
    logic         io_diffCommits_info_38_vecWen;
    logic         io_diffCommits_info_38_v0Wen;
    logic         io_diffCommits_info_38_vlWen;
    logic [5:0]   io_diffCommits_info_39_ldest;
    logic [7:0]   io_diffCommits_info_39_pdest;
    logic         io_diffCommits_info_39_rfWen;
    logic         io_diffCommits_info_39_fpWen;
    logic         io_diffCommits_info_39_vecWen;
    logic         io_diffCommits_info_39_v0Wen;
    logic         io_diffCommits_info_39_vlWen;
    logic [5:0]   io_diffCommits_info_40_ldest;
    logic [7:0]   io_diffCommits_info_40_pdest;
    logic         io_diffCommits_info_40_rfWen;
    logic         io_diffCommits_info_40_fpWen;
    logic         io_diffCommits_info_40_vecWen;
    logic         io_diffCommits_info_40_v0Wen;
    logic         io_diffCommits_info_40_vlWen;
    logic [5:0]   io_diffCommits_info_41_ldest;
    logic [7:0]   io_diffCommits_info_41_pdest;
    logic         io_diffCommits_info_41_rfWen;
    logic         io_diffCommits_info_41_fpWen;
    logic         io_diffCommits_info_41_vecWen;
    logic         io_diffCommits_info_41_v0Wen;
    logic         io_diffCommits_info_41_vlWen;
    logic [5:0]   io_diffCommits_info_42_ldest;
    logic [7:0]   io_diffCommits_info_42_pdest;
    logic         io_diffCommits_info_42_rfWen;
    logic         io_diffCommits_info_42_fpWen;
    logic         io_diffCommits_info_42_vecWen;
    logic         io_diffCommits_info_42_v0Wen;
    logic         io_diffCommits_info_42_vlWen;
    logic [5:0]   io_diffCommits_info_43_ldest;
    logic [7:0]   io_diffCommits_info_43_pdest;
    logic         io_diffCommits_info_43_rfWen;
    logic         io_diffCommits_info_43_fpWen;
    logic         io_diffCommits_info_43_vecWen;
    logic         io_diffCommits_info_43_v0Wen;
    logic         io_diffCommits_info_43_vlWen;
    logic [5:0]   io_diffCommits_info_44_ldest;
    logic [7:0]   io_diffCommits_info_44_pdest;
    logic         io_diffCommits_info_44_rfWen;
    logic         io_diffCommits_info_44_fpWen;
    logic         io_diffCommits_info_44_vecWen;
    logic         io_diffCommits_info_44_v0Wen;
    logic         io_diffCommits_info_44_vlWen;
    logic [5:0]   io_diffCommits_info_45_ldest;
    logic [7:0]   io_diffCommits_info_45_pdest;
    logic         io_diffCommits_info_45_rfWen;
    logic         io_diffCommits_info_45_fpWen;
    logic         io_diffCommits_info_45_vecWen;
    logic         io_diffCommits_info_45_v0Wen;
    logic         io_diffCommits_info_45_vlWen;
    logic [5:0]   io_diffCommits_info_46_ldest;
    logic [7:0]   io_diffCommits_info_46_pdest;
    logic         io_diffCommits_info_46_rfWen;
    logic         io_diffCommits_info_46_fpWen;
    logic         io_diffCommits_info_46_vecWen;
    logic         io_diffCommits_info_46_v0Wen;
    logic         io_diffCommits_info_46_vlWen;
    logic [5:0]   io_diffCommits_info_47_ldest;
    logic [7:0]   io_diffCommits_info_47_pdest;
    logic         io_diffCommits_info_47_rfWen;
    logic         io_diffCommits_info_47_fpWen;
    logic         io_diffCommits_info_47_vecWen;
    logic         io_diffCommits_info_47_v0Wen;
    logic         io_diffCommits_info_47_vlWen;
    logic [5:0]   io_diffCommits_info_48_ldest;
    logic [7:0]   io_diffCommits_info_48_pdest;
    logic         io_diffCommits_info_48_rfWen;
    logic         io_diffCommits_info_48_fpWen;
    logic         io_diffCommits_info_48_vecWen;
    logic         io_diffCommits_info_48_v0Wen;
    logic         io_diffCommits_info_48_vlWen;
    logic [5:0]   io_diffCommits_info_49_ldest;
    logic [7:0]   io_diffCommits_info_49_pdest;
    logic         io_diffCommits_info_49_rfWen;
    logic         io_diffCommits_info_49_fpWen;
    logic         io_diffCommits_info_49_vecWen;
    logic         io_diffCommits_info_49_v0Wen;
    logic         io_diffCommits_info_49_vlWen;
    logic [5:0]   io_diffCommits_info_50_ldest;
    logic [7:0]   io_diffCommits_info_50_pdest;
    logic         io_diffCommits_info_50_rfWen;
    logic         io_diffCommits_info_50_fpWen;
    logic         io_diffCommits_info_50_vecWen;
    logic         io_diffCommits_info_50_v0Wen;
    logic         io_diffCommits_info_50_vlWen;
    logic [5:0]   io_diffCommits_info_51_ldest;
    logic [7:0]   io_diffCommits_info_51_pdest;
    logic         io_diffCommits_info_51_rfWen;
    logic         io_diffCommits_info_51_fpWen;
    logic         io_diffCommits_info_51_vecWen;
    logic         io_diffCommits_info_51_v0Wen;
    logic         io_diffCommits_info_51_vlWen;
    logic [5:0]   io_diffCommits_info_52_ldest;
    logic [7:0]   io_diffCommits_info_52_pdest;
    logic         io_diffCommits_info_52_rfWen;
    logic         io_diffCommits_info_52_fpWen;
    logic         io_diffCommits_info_52_vecWen;
    logic         io_diffCommits_info_52_v0Wen;
    logic         io_diffCommits_info_52_vlWen;
    logic [5:0]   io_diffCommits_info_53_ldest;
    logic [7:0]   io_diffCommits_info_53_pdest;
    logic         io_diffCommits_info_53_rfWen;
    logic         io_diffCommits_info_53_fpWen;
    logic         io_diffCommits_info_53_vecWen;
    logic         io_diffCommits_info_53_v0Wen;
    logic         io_diffCommits_info_53_vlWen;
    logic [5:0]   io_diffCommits_info_54_ldest;
    logic [7:0]   io_diffCommits_info_54_pdest;
    logic         io_diffCommits_info_54_rfWen;
    logic         io_diffCommits_info_54_fpWen;
    logic         io_diffCommits_info_54_vecWen;
    logic         io_diffCommits_info_54_v0Wen;
    logic         io_diffCommits_info_54_vlWen;
    logic [5:0]   io_diffCommits_info_55_ldest;
    logic [7:0]   io_diffCommits_info_55_pdest;
    logic         io_diffCommits_info_55_rfWen;
    logic         io_diffCommits_info_55_fpWen;
    logic         io_diffCommits_info_55_vecWen;
    logic         io_diffCommits_info_55_v0Wen;
    logic         io_diffCommits_info_55_vlWen;
    logic [5:0]   io_diffCommits_info_56_ldest;
    logic [7:0]   io_diffCommits_info_56_pdest;
    logic         io_diffCommits_info_56_rfWen;
    logic         io_diffCommits_info_56_fpWen;
    logic         io_diffCommits_info_56_vecWen;
    logic         io_diffCommits_info_56_v0Wen;
    logic         io_diffCommits_info_56_vlWen;
    logic [5:0]   io_diffCommits_info_57_ldest;
    logic [7:0]   io_diffCommits_info_57_pdest;
    logic         io_diffCommits_info_57_rfWen;
    logic         io_diffCommits_info_57_fpWen;
    logic         io_diffCommits_info_57_vecWen;
    logic         io_diffCommits_info_57_v0Wen;
    logic         io_diffCommits_info_57_vlWen;
    logic [5:0]   io_diffCommits_info_58_ldest;
    logic [7:0]   io_diffCommits_info_58_pdest;
    logic         io_diffCommits_info_58_rfWen;
    logic         io_diffCommits_info_58_fpWen;
    logic         io_diffCommits_info_58_vecWen;
    logic         io_diffCommits_info_58_v0Wen;
    logic         io_diffCommits_info_58_vlWen;
    logic [5:0]   io_diffCommits_info_59_ldest;
    logic [7:0]   io_diffCommits_info_59_pdest;
    logic         io_diffCommits_info_59_rfWen;
    logic         io_diffCommits_info_59_fpWen;
    logic         io_diffCommits_info_59_vecWen;
    logic         io_diffCommits_info_59_v0Wen;
    logic         io_diffCommits_info_59_vlWen;
    logic [5:0]   io_diffCommits_info_60_ldest;
    logic [7:0]   io_diffCommits_info_60_pdest;
    logic         io_diffCommits_info_60_rfWen;
    logic         io_diffCommits_info_60_fpWen;
    logic         io_diffCommits_info_60_vecWen;
    logic         io_diffCommits_info_60_v0Wen;
    logic         io_diffCommits_info_60_vlWen;
    logic [5:0]   io_diffCommits_info_61_ldest;
    logic [7:0]   io_diffCommits_info_61_pdest;
    logic         io_diffCommits_info_61_rfWen;
    logic         io_diffCommits_info_61_fpWen;
    logic         io_diffCommits_info_61_vecWen;
    logic         io_diffCommits_info_61_v0Wen;
    logic         io_diffCommits_info_61_vlWen;
    logic [5:0]   io_diffCommits_info_62_ldest;
    logic [7:0]   io_diffCommits_info_62_pdest;
    logic         io_diffCommits_info_62_rfWen;
    logic         io_diffCommits_info_62_fpWen;
    logic         io_diffCommits_info_62_vecWen;
    logic         io_diffCommits_info_62_v0Wen;
    logic         io_diffCommits_info_62_vlWen;
    logic [5:0]   io_diffCommits_info_63_ldest;
    logic [7:0]   io_diffCommits_info_63_pdest;
    logic         io_diffCommits_info_63_rfWen;
    logic         io_diffCommits_info_63_fpWen;
    logic         io_diffCommits_info_63_vecWen;
    logic         io_diffCommits_info_63_v0Wen;
    logic         io_diffCommits_info_63_vlWen;
    logic [5:0]   io_diffCommits_info_64_ldest;
    logic [7:0]   io_diffCommits_info_64_pdest;
    logic         io_diffCommits_info_64_rfWen;
    logic         io_diffCommits_info_64_fpWen;
    logic         io_diffCommits_info_64_vecWen;
    logic         io_diffCommits_info_64_v0Wen;
    logic         io_diffCommits_info_64_vlWen;
    logic [5:0]   io_diffCommits_info_65_ldest;
    logic [7:0]   io_diffCommits_info_65_pdest;
    logic         io_diffCommits_info_65_rfWen;
    logic         io_diffCommits_info_65_fpWen;
    logic         io_diffCommits_info_65_vecWen;
    logic         io_diffCommits_info_65_v0Wen;
    logic         io_diffCommits_info_65_vlWen;
    logic [5:0]   io_diffCommits_info_66_ldest;
    logic [7:0]   io_diffCommits_info_66_pdest;
    logic         io_diffCommits_info_66_rfWen;
    logic         io_diffCommits_info_66_fpWen;
    logic         io_diffCommits_info_66_vecWen;
    logic         io_diffCommits_info_66_v0Wen;
    logic         io_diffCommits_info_66_vlWen;
    logic [5:0]   io_diffCommits_info_67_ldest;
    logic [7:0]   io_diffCommits_info_67_pdest;
    logic         io_diffCommits_info_67_rfWen;
    logic         io_diffCommits_info_67_fpWen;
    logic         io_diffCommits_info_67_vecWen;
    logic         io_diffCommits_info_67_v0Wen;
    logic         io_diffCommits_info_67_vlWen;
    logic [5:0]   io_diffCommits_info_68_ldest;
    logic [7:0]   io_diffCommits_info_68_pdest;
    logic         io_diffCommits_info_68_rfWen;
    logic         io_diffCommits_info_68_fpWen;
    logic         io_diffCommits_info_68_vecWen;
    logic         io_diffCommits_info_68_v0Wen;
    logic         io_diffCommits_info_68_vlWen;
    logic [5:0]   io_diffCommits_info_69_ldest;
    logic [7:0]   io_diffCommits_info_69_pdest;
    logic         io_diffCommits_info_69_rfWen;
    logic         io_diffCommits_info_69_fpWen;
    logic         io_diffCommits_info_69_vecWen;
    logic         io_diffCommits_info_69_v0Wen;
    logic         io_diffCommits_info_69_vlWen;
    logic [5:0]   io_diffCommits_info_70_ldest;
    logic [7:0]   io_diffCommits_info_70_pdest;
    logic         io_diffCommits_info_70_rfWen;
    logic         io_diffCommits_info_70_fpWen;
    logic         io_diffCommits_info_70_vecWen;
    logic         io_diffCommits_info_70_v0Wen;
    logic         io_diffCommits_info_70_vlWen;
    logic [5:0]   io_diffCommits_info_71_ldest;
    logic [7:0]   io_diffCommits_info_71_pdest;
    logic         io_diffCommits_info_71_rfWen;
    logic         io_diffCommits_info_71_fpWen;
    logic         io_diffCommits_info_71_vecWen;
    logic         io_diffCommits_info_71_v0Wen;
    logic         io_diffCommits_info_71_vlWen;
    logic [5:0]   io_diffCommits_info_72_ldest;
    logic [7:0]   io_diffCommits_info_72_pdest;
    logic         io_diffCommits_info_72_rfWen;
    logic         io_diffCommits_info_72_fpWen;
    logic         io_diffCommits_info_72_vecWen;
    logic         io_diffCommits_info_72_v0Wen;
    logic         io_diffCommits_info_72_vlWen;
    logic [5:0]   io_diffCommits_info_73_ldest;
    logic [7:0]   io_diffCommits_info_73_pdest;
    logic         io_diffCommits_info_73_rfWen;
    logic         io_diffCommits_info_73_fpWen;
    logic         io_diffCommits_info_73_vecWen;
    logic         io_diffCommits_info_73_v0Wen;
    logic         io_diffCommits_info_73_vlWen;
    logic [5:0]   io_diffCommits_info_74_ldest;
    logic [7:0]   io_diffCommits_info_74_pdest;
    logic         io_diffCommits_info_74_rfWen;
    logic         io_diffCommits_info_74_fpWen;
    logic         io_diffCommits_info_74_vecWen;
    logic         io_diffCommits_info_74_v0Wen;
    logic         io_diffCommits_info_74_vlWen;
    logic [5:0]   io_diffCommits_info_75_ldest;
    logic [7:0]   io_diffCommits_info_75_pdest;
    logic         io_diffCommits_info_75_rfWen;
    logic         io_diffCommits_info_75_fpWen;
    logic         io_diffCommits_info_75_vecWen;
    logic         io_diffCommits_info_75_v0Wen;
    logic         io_diffCommits_info_75_vlWen;
    logic [5:0]   io_diffCommits_info_76_ldest;
    logic [7:0]   io_diffCommits_info_76_pdest;
    logic         io_diffCommits_info_76_rfWen;
    logic         io_diffCommits_info_76_fpWen;
    logic         io_diffCommits_info_76_vecWen;
    logic         io_diffCommits_info_76_v0Wen;
    logic         io_diffCommits_info_76_vlWen;
    logic [5:0]   io_diffCommits_info_77_ldest;
    logic [7:0]   io_diffCommits_info_77_pdest;
    logic         io_diffCommits_info_77_rfWen;
    logic         io_diffCommits_info_77_fpWen;
    logic         io_diffCommits_info_77_vecWen;
    logic         io_diffCommits_info_77_v0Wen;
    logic         io_diffCommits_info_77_vlWen;
    logic [5:0]   io_diffCommits_info_78_ldest;
    logic [7:0]   io_diffCommits_info_78_pdest;
    logic         io_diffCommits_info_78_rfWen;
    logic         io_diffCommits_info_78_fpWen;
    logic         io_diffCommits_info_78_vecWen;
    logic         io_diffCommits_info_78_v0Wen;
    logic         io_diffCommits_info_78_vlWen;
    logic [5:0]   io_diffCommits_info_79_ldest;
    logic [7:0]   io_diffCommits_info_79_pdest;
    logic         io_diffCommits_info_79_rfWen;
    logic         io_diffCommits_info_79_fpWen;
    logic         io_diffCommits_info_79_vecWen;
    logic         io_diffCommits_info_79_v0Wen;
    logic         io_diffCommits_info_79_vlWen;
    logic [5:0]   io_diffCommits_info_80_ldest;
    logic [7:0]   io_diffCommits_info_80_pdest;
    logic         io_diffCommits_info_80_rfWen;
    logic         io_diffCommits_info_80_fpWen;
    logic         io_diffCommits_info_80_vecWen;
    logic         io_diffCommits_info_80_v0Wen;
    logic         io_diffCommits_info_80_vlWen;
    logic [5:0]   io_diffCommits_info_81_ldest;
    logic [7:0]   io_diffCommits_info_81_pdest;
    logic         io_diffCommits_info_81_rfWen;
    logic         io_diffCommits_info_81_fpWen;
    logic         io_diffCommits_info_81_vecWen;
    logic         io_diffCommits_info_81_v0Wen;
    logic         io_diffCommits_info_81_vlWen;
    logic [5:0]   io_diffCommits_info_82_ldest;
    logic [7:0]   io_diffCommits_info_82_pdest;
    logic         io_diffCommits_info_82_rfWen;
    logic         io_diffCommits_info_82_fpWen;
    logic         io_diffCommits_info_82_vecWen;
    logic         io_diffCommits_info_82_v0Wen;
    logic         io_diffCommits_info_82_vlWen;
    logic [5:0]   io_diffCommits_info_83_ldest;
    logic [7:0]   io_diffCommits_info_83_pdest;
    logic         io_diffCommits_info_83_rfWen;
    logic         io_diffCommits_info_83_fpWen;
    logic         io_diffCommits_info_83_vecWen;
    logic         io_diffCommits_info_83_v0Wen;
    logic         io_diffCommits_info_83_vlWen;
    logic [5:0]   io_diffCommits_info_84_ldest;
    logic [7:0]   io_diffCommits_info_84_pdest;
    logic         io_diffCommits_info_84_rfWen;
    logic         io_diffCommits_info_84_fpWen;
    logic         io_diffCommits_info_84_vecWen;
    logic         io_diffCommits_info_84_v0Wen;
    logic         io_diffCommits_info_84_vlWen;
    logic [5:0]   io_diffCommits_info_85_ldest;
    logic [7:0]   io_diffCommits_info_85_pdest;
    logic         io_diffCommits_info_85_rfWen;
    logic         io_diffCommits_info_85_fpWen;
    logic         io_diffCommits_info_85_vecWen;
    logic         io_diffCommits_info_85_v0Wen;
    logic         io_diffCommits_info_85_vlWen;
    logic [5:0]   io_diffCommits_info_86_ldest;
    logic [7:0]   io_diffCommits_info_86_pdest;
    logic         io_diffCommits_info_86_rfWen;
    logic         io_diffCommits_info_86_fpWen;
    logic         io_diffCommits_info_86_vecWen;
    logic         io_diffCommits_info_86_v0Wen;
    logic         io_diffCommits_info_86_vlWen;
    logic [5:0]   io_diffCommits_info_87_ldest;
    logic [7:0]   io_diffCommits_info_87_pdest;
    logic         io_diffCommits_info_87_rfWen;
    logic         io_diffCommits_info_87_fpWen;
    logic         io_diffCommits_info_87_vecWen;
    logic         io_diffCommits_info_87_v0Wen;
    logic         io_diffCommits_info_87_vlWen;
    logic [5:0]   io_diffCommits_info_88_ldest;
    logic [7:0]   io_diffCommits_info_88_pdest;
    logic         io_diffCommits_info_88_rfWen;
    logic         io_diffCommits_info_88_fpWen;
    logic         io_diffCommits_info_88_vecWen;
    logic         io_diffCommits_info_88_v0Wen;
    logic         io_diffCommits_info_88_vlWen;
    logic [5:0]   io_diffCommits_info_89_ldest;
    logic [7:0]   io_diffCommits_info_89_pdest;
    logic         io_diffCommits_info_89_rfWen;
    logic         io_diffCommits_info_89_fpWen;
    logic         io_diffCommits_info_89_vecWen;
    logic         io_diffCommits_info_89_v0Wen;
    logic         io_diffCommits_info_89_vlWen;
    logic [5:0]   io_diffCommits_info_90_ldest;
    logic [7:0]   io_diffCommits_info_90_pdest;
    logic         io_diffCommits_info_90_rfWen;
    logic         io_diffCommits_info_90_fpWen;
    logic         io_diffCommits_info_90_vecWen;
    logic         io_diffCommits_info_90_v0Wen;
    logic         io_diffCommits_info_90_vlWen;
    logic [5:0]   io_diffCommits_info_91_ldest;
    logic [7:0]   io_diffCommits_info_91_pdest;
    logic         io_diffCommits_info_91_rfWen;
    logic         io_diffCommits_info_91_fpWen;
    logic         io_diffCommits_info_91_vecWen;
    logic         io_diffCommits_info_91_v0Wen;
    logic         io_diffCommits_info_91_vlWen;
    logic [5:0]   io_diffCommits_info_92_ldest;
    logic [7:0]   io_diffCommits_info_92_pdest;
    logic         io_diffCommits_info_92_rfWen;
    logic         io_diffCommits_info_92_fpWen;
    logic         io_diffCommits_info_92_vecWen;
    logic         io_diffCommits_info_92_v0Wen;
    logic         io_diffCommits_info_92_vlWen;
    logic [5:0]   io_diffCommits_info_93_ldest;
    logic [7:0]   io_diffCommits_info_93_pdest;
    logic         io_diffCommits_info_93_rfWen;
    logic         io_diffCommits_info_93_fpWen;
    logic         io_diffCommits_info_93_vecWen;
    logic         io_diffCommits_info_93_v0Wen;
    logic         io_diffCommits_info_93_vlWen;
    logic [5:0]   io_diffCommits_info_94_ldest;
    logic [7:0]   io_diffCommits_info_94_pdest;
    logic         io_diffCommits_info_94_rfWen;
    logic         io_diffCommits_info_94_fpWen;
    logic         io_diffCommits_info_94_vecWen;
    logic         io_diffCommits_info_94_v0Wen;
    logic         io_diffCommits_info_94_vlWen;
    logic [5:0]   io_diffCommits_info_95_ldest;
    logic [7:0]   io_diffCommits_info_95_pdest;
    logic         io_diffCommits_info_95_rfWen;
    logic         io_diffCommits_info_95_fpWen;
    logic         io_diffCommits_info_95_vecWen;
    logic         io_diffCommits_info_95_v0Wen;
    logic         io_diffCommits_info_95_vlWen;
    logic [5:0]   io_diffCommits_info_96_ldest;
    logic [7:0]   io_diffCommits_info_96_pdest;
    logic         io_diffCommits_info_96_rfWen;
    logic         io_diffCommits_info_96_fpWen;
    logic         io_diffCommits_info_96_vecWen;
    logic         io_diffCommits_info_96_v0Wen;
    logic         io_diffCommits_info_96_vlWen;
    logic [5:0]   io_diffCommits_info_97_ldest;
    logic [7:0]   io_diffCommits_info_97_pdest;
    logic         io_diffCommits_info_97_rfWen;
    logic         io_diffCommits_info_97_fpWen;
    logic         io_diffCommits_info_97_vecWen;
    logic         io_diffCommits_info_97_v0Wen;
    logic         io_diffCommits_info_97_vlWen;
    logic [5:0]   io_diffCommits_info_98_ldest;
    logic [7:0]   io_diffCommits_info_98_pdest;
    logic         io_diffCommits_info_98_rfWen;
    logic         io_diffCommits_info_98_fpWen;
    logic         io_diffCommits_info_98_vecWen;
    logic         io_diffCommits_info_98_v0Wen;
    logic         io_diffCommits_info_98_vlWen;
    logic [5:0]   io_diffCommits_info_99_ldest;
    logic [7:0]   io_diffCommits_info_99_pdest;
    logic         io_diffCommits_info_99_rfWen;
    logic         io_diffCommits_info_99_fpWen;
    logic         io_diffCommits_info_99_vecWen;
    logic         io_diffCommits_info_99_v0Wen;
    logic         io_diffCommits_info_99_vlWen;
    logic [5:0]   io_diffCommits_info_100_ldest;
    logic [7:0]   io_diffCommits_info_100_pdest;
    logic         io_diffCommits_info_100_rfWen;
    logic         io_diffCommits_info_100_fpWen;
    logic         io_diffCommits_info_100_vecWen;
    logic         io_diffCommits_info_100_v0Wen;
    logic         io_diffCommits_info_100_vlWen;
    logic [5:0]   io_diffCommits_info_101_ldest;
    logic [7:0]   io_diffCommits_info_101_pdest;
    logic         io_diffCommits_info_101_rfWen;
    logic         io_diffCommits_info_101_fpWen;
    logic         io_diffCommits_info_101_vecWen;
    logic         io_diffCommits_info_101_v0Wen;
    logic         io_diffCommits_info_101_vlWen;
    logic [5:0]   io_diffCommits_info_102_ldest;
    logic [7:0]   io_diffCommits_info_102_pdest;
    logic         io_diffCommits_info_102_rfWen;
    logic         io_diffCommits_info_102_fpWen;
    logic         io_diffCommits_info_102_vecWen;
    logic         io_diffCommits_info_102_v0Wen;
    logic         io_diffCommits_info_102_vlWen;
    logic [5:0]   io_diffCommits_info_103_ldest;
    logic [7:0]   io_diffCommits_info_103_pdest;
    logic         io_diffCommits_info_103_rfWen;
    logic         io_diffCommits_info_103_fpWen;
    logic         io_diffCommits_info_103_vecWen;
    logic         io_diffCommits_info_103_v0Wen;
    logic         io_diffCommits_info_103_vlWen;
    logic [5:0]   io_diffCommits_info_104_ldest;
    logic [7:0]   io_diffCommits_info_104_pdest;
    logic         io_diffCommits_info_104_rfWen;
    logic         io_diffCommits_info_104_fpWen;
    logic         io_diffCommits_info_104_vecWen;
    logic         io_diffCommits_info_104_v0Wen;
    logic         io_diffCommits_info_104_vlWen;
    logic [5:0]   io_diffCommits_info_105_ldest;
    logic [7:0]   io_diffCommits_info_105_pdest;
    logic         io_diffCommits_info_105_rfWen;
    logic         io_diffCommits_info_105_fpWen;
    logic         io_diffCommits_info_105_vecWen;
    logic         io_diffCommits_info_105_v0Wen;
    logic         io_diffCommits_info_105_vlWen;
    logic [5:0]   io_diffCommits_info_106_ldest;
    logic [7:0]   io_diffCommits_info_106_pdest;
    logic         io_diffCommits_info_106_rfWen;
    logic         io_diffCommits_info_106_fpWen;
    logic         io_diffCommits_info_106_vecWen;
    logic         io_diffCommits_info_106_v0Wen;
    logic         io_diffCommits_info_106_vlWen;
    logic [5:0]   io_diffCommits_info_107_ldest;
    logic [7:0]   io_diffCommits_info_107_pdest;
    logic         io_diffCommits_info_107_rfWen;
    logic         io_diffCommits_info_107_fpWen;
    logic         io_diffCommits_info_107_vecWen;
    logic         io_diffCommits_info_107_v0Wen;
    logic         io_diffCommits_info_107_vlWen;
    logic [5:0]   io_diffCommits_info_108_ldest;
    logic [7:0]   io_diffCommits_info_108_pdest;
    logic         io_diffCommits_info_108_rfWen;
    logic         io_diffCommits_info_108_fpWen;
    logic         io_diffCommits_info_108_vecWen;
    logic         io_diffCommits_info_108_v0Wen;
    logic         io_diffCommits_info_108_vlWen;
    logic [5:0]   io_diffCommits_info_109_ldest;
    logic [7:0]   io_diffCommits_info_109_pdest;
    logic         io_diffCommits_info_109_rfWen;
    logic         io_diffCommits_info_109_fpWen;
    logic         io_diffCommits_info_109_vecWen;
    logic         io_diffCommits_info_109_v0Wen;
    logic         io_diffCommits_info_109_vlWen;
    logic [5:0]   io_diffCommits_info_110_ldest;
    logic [7:0]   io_diffCommits_info_110_pdest;
    logic         io_diffCommits_info_110_rfWen;
    logic         io_diffCommits_info_110_fpWen;
    logic         io_diffCommits_info_110_vecWen;
    logic         io_diffCommits_info_110_v0Wen;
    logic         io_diffCommits_info_110_vlWen;
    logic [5:0]   io_diffCommits_info_111_ldest;
    logic [7:0]   io_diffCommits_info_111_pdest;
    logic         io_diffCommits_info_111_rfWen;
    logic         io_diffCommits_info_111_fpWen;
    logic         io_diffCommits_info_111_vecWen;
    logic         io_diffCommits_info_111_v0Wen;
    logic         io_diffCommits_info_111_vlWen;
    logic [5:0]   io_diffCommits_info_112_ldest;
    logic [7:0]   io_diffCommits_info_112_pdest;
    logic         io_diffCommits_info_112_rfWen;
    logic         io_diffCommits_info_112_fpWen;
    logic         io_diffCommits_info_112_vecWen;
    logic         io_diffCommits_info_112_v0Wen;
    logic         io_diffCommits_info_112_vlWen;
    logic [5:0]   io_diffCommits_info_113_ldest;
    logic [7:0]   io_diffCommits_info_113_pdest;
    logic         io_diffCommits_info_113_rfWen;
    logic         io_diffCommits_info_113_fpWen;
    logic         io_diffCommits_info_113_vecWen;
    logic         io_diffCommits_info_113_v0Wen;
    logic         io_diffCommits_info_113_vlWen;
    logic [5:0]   io_diffCommits_info_114_ldest;
    logic [7:0]   io_diffCommits_info_114_pdest;
    logic         io_diffCommits_info_114_rfWen;
    logic         io_diffCommits_info_114_fpWen;
    logic         io_diffCommits_info_114_vecWen;
    logic         io_diffCommits_info_114_v0Wen;
    logic         io_diffCommits_info_114_vlWen;
    logic [5:0]   io_diffCommits_info_115_ldest;
    logic [7:0]   io_diffCommits_info_115_pdest;
    logic         io_diffCommits_info_115_rfWen;
    logic         io_diffCommits_info_115_fpWen;
    logic         io_diffCommits_info_115_vecWen;
    logic         io_diffCommits_info_115_v0Wen;
    logic         io_diffCommits_info_115_vlWen;
    logic [5:0]   io_diffCommits_info_116_ldest;
    logic [7:0]   io_diffCommits_info_116_pdest;
    logic         io_diffCommits_info_116_rfWen;
    logic         io_diffCommits_info_116_fpWen;
    logic         io_diffCommits_info_116_vecWen;
    logic         io_diffCommits_info_116_v0Wen;
    logic         io_diffCommits_info_116_vlWen;
    logic [5:0]   io_diffCommits_info_117_ldest;
    logic [7:0]   io_diffCommits_info_117_pdest;
    logic         io_diffCommits_info_117_rfWen;
    logic         io_diffCommits_info_117_fpWen;
    logic         io_diffCommits_info_117_vecWen;
    logic         io_diffCommits_info_117_v0Wen;
    logic         io_diffCommits_info_117_vlWen;
    logic [5:0]   io_diffCommits_info_118_ldest;
    logic [7:0]   io_diffCommits_info_118_pdest;
    logic         io_diffCommits_info_118_rfWen;
    logic         io_diffCommits_info_118_fpWen;
    logic         io_diffCommits_info_118_vecWen;
    logic         io_diffCommits_info_118_v0Wen;
    logic         io_diffCommits_info_118_vlWen;
    logic [5:0]   io_diffCommits_info_119_ldest;
    logic [7:0]   io_diffCommits_info_119_pdest;
    logic         io_diffCommits_info_119_rfWen;
    logic         io_diffCommits_info_119_fpWen;
    logic         io_diffCommits_info_119_vecWen;
    logic         io_diffCommits_info_119_v0Wen;
    logic         io_diffCommits_info_119_vlWen;
    logic [5:0]   io_diffCommits_info_120_ldest;
    logic [7:0]   io_diffCommits_info_120_pdest;
    logic         io_diffCommits_info_120_rfWen;
    logic         io_diffCommits_info_120_fpWen;
    logic         io_diffCommits_info_120_vecWen;
    logic         io_diffCommits_info_120_v0Wen;
    logic         io_diffCommits_info_120_vlWen;
    logic [5:0]   io_diffCommits_info_121_ldest;
    logic [7:0]   io_diffCommits_info_121_pdest;
    logic         io_diffCommits_info_121_rfWen;
    logic         io_diffCommits_info_121_fpWen;
    logic         io_diffCommits_info_121_vecWen;
    logic         io_diffCommits_info_121_v0Wen;
    logic         io_diffCommits_info_121_vlWen;
    logic [5:0]   io_diffCommits_info_122_ldest;
    logic [7:0]   io_diffCommits_info_122_pdest;
    logic         io_diffCommits_info_122_rfWen;
    logic         io_diffCommits_info_122_fpWen;
    logic         io_diffCommits_info_122_vecWen;
    logic         io_diffCommits_info_122_v0Wen;
    logic         io_diffCommits_info_122_vlWen;
    logic [5:0]   io_diffCommits_info_123_ldest;
    logic [7:0]   io_diffCommits_info_123_pdest;
    logic         io_diffCommits_info_123_rfWen;
    logic         io_diffCommits_info_123_fpWen;
    logic         io_diffCommits_info_123_vecWen;
    logic         io_diffCommits_info_123_v0Wen;
    logic         io_diffCommits_info_123_vlWen;
    logic [5:0]   io_diffCommits_info_124_ldest;
    logic [7:0]   io_diffCommits_info_124_pdest;
    logic         io_diffCommits_info_124_rfWen;
    logic         io_diffCommits_info_124_fpWen;
    logic         io_diffCommits_info_124_vecWen;
    logic         io_diffCommits_info_124_v0Wen;
    logic         io_diffCommits_info_124_vlWen;
    logic [5:0]   io_diffCommits_info_125_ldest;
    logic [7:0]   io_diffCommits_info_125_pdest;
    logic         io_diffCommits_info_125_rfWen;
    logic         io_diffCommits_info_125_fpWen;
    logic         io_diffCommits_info_125_vecWen;
    logic         io_diffCommits_info_125_v0Wen;
    logic         io_diffCommits_info_125_vlWen;
    logic [5:0]   io_diffCommits_info_126_ldest;
    logic [7:0]   io_diffCommits_info_126_pdest;
    logic         io_diffCommits_info_126_rfWen;
    logic         io_diffCommits_info_126_fpWen;
    logic         io_diffCommits_info_126_vecWen;
    logic         io_diffCommits_info_126_v0Wen;
    logic         io_diffCommits_info_126_vlWen;
    logic [5:0]   io_diffCommits_info_127_ldest;
    logic [7:0]   io_diffCommits_info_127_pdest;
    logic         io_diffCommits_info_127_rfWen;
    logic         io_diffCommits_info_127_fpWen;
    logic         io_diffCommits_info_127_vecWen;
    logic         io_diffCommits_info_127_v0Wen;
    logic         io_diffCommits_info_127_vlWen;
    logic [5:0]   io_diffCommits_info_128_ldest;
    logic [7:0]   io_diffCommits_info_128_pdest;
    logic         io_diffCommits_info_128_rfWen;
    logic         io_diffCommits_info_128_fpWen;
    logic         io_diffCommits_info_128_vecWen;
    logic         io_diffCommits_info_128_v0Wen;
    logic         io_diffCommits_info_128_vlWen;
    logic [5:0]   io_diffCommits_info_129_ldest;
    logic [7:0]   io_diffCommits_info_129_pdest;
    logic         io_diffCommits_info_129_rfWen;
    logic         io_diffCommits_info_129_fpWen;
    logic         io_diffCommits_info_129_vecWen;
    logic         io_diffCommits_info_129_v0Wen;
    logic         io_diffCommits_info_129_vlWen;
    logic [5:0]   io_diffCommits_info_130_ldest;
    logic [7:0]   io_diffCommits_info_130_pdest;
    logic         io_diffCommits_info_130_rfWen;
    logic         io_diffCommits_info_130_fpWen;
    logic         io_diffCommits_info_130_vecWen;
    logic         io_diffCommits_info_130_v0Wen;
    logic         io_diffCommits_info_130_vlWen;
    logic [5:0]   io_diffCommits_info_131_ldest;
    logic [7:0]   io_diffCommits_info_131_pdest;
    logic         io_diffCommits_info_131_rfWen;
    logic         io_diffCommits_info_131_fpWen;
    logic         io_diffCommits_info_131_vecWen;
    logic         io_diffCommits_info_131_v0Wen;
    logic         io_diffCommits_info_131_vlWen;
    logic [5:0]   io_diffCommits_info_132_ldest;
    logic [7:0]   io_diffCommits_info_132_pdest;
    logic         io_diffCommits_info_132_rfWen;
    logic         io_diffCommits_info_132_fpWen;
    logic         io_diffCommits_info_132_vecWen;
    logic         io_diffCommits_info_132_v0Wen;
    logic         io_diffCommits_info_132_vlWen;
    logic [5:0]   io_diffCommits_info_133_ldest;
    logic [7:0]   io_diffCommits_info_133_pdest;
    logic         io_diffCommits_info_133_rfWen;
    logic         io_diffCommits_info_133_fpWen;
    logic         io_diffCommits_info_133_vecWen;
    logic         io_diffCommits_info_133_v0Wen;
    logic         io_diffCommits_info_133_vlWen;
    logic [5:0]   io_diffCommits_info_134_ldest;
    logic [7:0]   io_diffCommits_info_134_pdest;
    logic         io_diffCommits_info_134_rfWen;
    logic         io_diffCommits_info_134_fpWen;
    logic         io_diffCommits_info_134_vecWen;
    logic         io_diffCommits_info_134_v0Wen;
    logic         io_diffCommits_info_134_vlWen;
    logic [5:0]   io_diffCommits_info_135_ldest;
    logic [7:0]   io_diffCommits_info_135_pdest;
    logic         io_diffCommits_info_135_rfWen;
    logic         io_diffCommits_info_135_fpWen;
    logic         io_diffCommits_info_135_vecWen;
    logic         io_diffCommits_info_135_v0Wen;
    logic         io_diffCommits_info_135_vlWen;
    logic [5:0]   io_diffCommits_info_136_ldest;
    logic [7:0]   io_diffCommits_info_136_pdest;
    logic         io_diffCommits_info_136_rfWen;
    logic         io_diffCommits_info_136_fpWen;
    logic         io_diffCommits_info_136_vecWen;
    logic         io_diffCommits_info_136_v0Wen;
    logic         io_diffCommits_info_136_vlWen;
    logic [5:0]   io_diffCommits_info_137_ldest;
    logic [7:0]   io_diffCommits_info_137_pdest;
    logic         io_diffCommits_info_137_rfWen;
    logic         io_diffCommits_info_137_fpWen;
    logic         io_diffCommits_info_137_vecWen;
    logic         io_diffCommits_info_137_v0Wen;
    logic         io_diffCommits_info_137_vlWen;
    logic [5:0]   io_diffCommits_info_138_ldest;
    logic [7:0]   io_diffCommits_info_138_pdest;
    logic         io_diffCommits_info_138_rfWen;
    logic         io_diffCommits_info_138_fpWen;
    logic         io_diffCommits_info_138_vecWen;
    logic         io_diffCommits_info_138_v0Wen;
    logic         io_diffCommits_info_138_vlWen;
    logic [5:0]   io_diffCommits_info_139_ldest;
    logic [7:0]   io_diffCommits_info_139_pdest;
    logic         io_diffCommits_info_139_rfWen;
    logic         io_diffCommits_info_139_fpWen;
    logic         io_diffCommits_info_139_vecWen;
    logic         io_diffCommits_info_139_v0Wen;
    logic         io_diffCommits_info_139_vlWen;
    logic [5:0]   io_diffCommits_info_140_ldest;
    logic [7:0]   io_diffCommits_info_140_pdest;
    logic         io_diffCommits_info_140_rfWen;
    logic         io_diffCommits_info_140_fpWen;
    logic         io_diffCommits_info_140_vecWen;
    logic         io_diffCommits_info_140_v0Wen;
    logic         io_diffCommits_info_140_vlWen;
    logic [5:0]   io_diffCommits_info_141_ldest;
    logic [7:0]   io_diffCommits_info_141_pdest;
    logic         io_diffCommits_info_141_rfWen;
    logic         io_diffCommits_info_141_fpWen;
    logic         io_diffCommits_info_141_vecWen;
    logic         io_diffCommits_info_141_v0Wen;
    logic         io_diffCommits_info_141_vlWen;
    logic [5:0]   io_diffCommits_info_142_ldest;
    logic [7:0]   io_diffCommits_info_142_pdest;
    logic         io_diffCommits_info_142_rfWen;
    logic         io_diffCommits_info_142_fpWen;
    logic         io_diffCommits_info_142_vecWen;
    logic         io_diffCommits_info_142_v0Wen;
    logic         io_diffCommits_info_142_vlWen;
    logic [5:0]   io_diffCommits_info_143_ldest;
    logic [7:0]   io_diffCommits_info_143_pdest;
    logic         io_diffCommits_info_143_rfWen;
    logic         io_diffCommits_info_143_fpWen;
    logic         io_diffCommits_info_143_vecWen;
    logic         io_diffCommits_info_143_v0Wen;
    logic         io_diffCommits_info_143_vlWen;
    logic [5:0]   io_diffCommits_info_144_ldest;
    logic [7:0]   io_diffCommits_info_144_pdest;
    logic         io_diffCommits_info_144_rfWen;
    logic         io_diffCommits_info_144_fpWen;
    logic         io_diffCommits_info_144_vecWen;
    logic         io_diffCommits_info_144_v0Wen;
    logic         io_diffCommits_info_144_vlWen;
    logic [5:0]   io_diffCommits_info_145_ldest;
    logic [7:0]   io_diffCommits_info_145_pdest;
    logic         io_diffCommits_info_145_rfWen;
    logic         io_diffCommits_info_145_fpWen;
    logic         io_diffCommits_info_145_vecWen;
    logic         io_diffCommits_info_145_v0Wen;
    logic         io_diffCommits_info_145_vlWen;
    logic [5:0]   io_diffCommits_info_146_ldest;
    logic [7:0]   io_diffCommits_info_146_pdest;
    logic         io_diffCommits_info_146_rfWen;
    logic         io_diffCommits_info_146_fpWen;
    logic         io_diffCommits_info_146_vecWen;
    logic         io_diffCommits_info_146_v0Wen;
    logic         io_diffCommits_info_146_vlWen;
    logic [5:0]   io_diffCommits_info_147_ldest;
    logic [7:0]   io_diffCommits_info_147_pdest;
    logic         io_diffCommits_info_147_rfWen;
    logic         io_diffCommits_info_147_fpWen;
    logic         io_diffCommits_info_147_vecWen;
    logic         io_diffCommits_info_147_v0Wen;
    logic         io_diffCommits_info_147_vlWen;
    logic [5:0]   io_diffCommits_info_148_ldest;
    logic [7:0]   io_diffCommits_info_148_pdest;
    logic         io_diffCommits_info_148_rfWen;
    logic         io_diffCommits_info_148_fpWen;
    logic         io_diffCommits_info_148_vecWen;
    logic         io_diffCommits_info_148_v0Wen;
    logic         io_diffCommits_info_148_vlWen;
    logic [5:0]   io_diffCommits_info_149_ldest;
    logic [7:0]   io_diffCommits_info_149_pdest;
    logic         io_diffCommits_info_149_rfWen;
    logic         io_diffCommits_info_149_fpWen;
    logic         io_diffCommits_info_149_vecWen;
    logic         io_diffCommits_info_149_v0Wen;
    logic         io_diffCommits_info_149_vlWen;
    logic [5:0]   io_diffCommits_info_150_ldest;
    logic [7:0]   io_diffCommits_info_150_pdest;
    logic         io_diffCommits_info_150_rfWen;
    logic         io_diffCommits_info_150_fpWen;
    logic         io_diffCommits_info_150_vecWen;
    logic         io_diffCommits_info_150_v0Wen;
    logic         io_diffCommits_info_150_vlWen;
    logic [5:0]   io_diffCommits_info_151_ldest;
    logic [7:0]   io_diffCommits_info_151_pdest;
    logic         io_diffCommits_info_151_rfWen;
    logic         io_diffCommits_info_151_fpWen;
    logic         io_diffCommits_info_151_vecWen;
    logic         io_diffCommits_info_151_v0Wen;
    logic         io_diffCommits_info_151_vlWen;
    logic [5:0]   io_diffCommits_info_152_ldest;
    logic [7:0]   io_diffCommits_info_152_pdest;
    logic         io_diffCommits_info_152_rfWen;
    logic         io_diffCommits_info_152_fpWen;
    logic         io_diffCommits_info_152_vecWen;
    logic         io_diffCommits_info_152_v0Wen;
    logic         io_diffCommits_info_152_vlWen;
    logic [5:0]   io_diffCommits_info_153_ldest;
    logic [7:0]   io_diffCommits_info_153_pdest;
    logic         io_diffCommits_info_153_rfWen;
    logic         io_diffCommits_info_153_fpWen;
    logic         io_diffCommits_info_153_vecWen;
    logic         io_diffCommits_info_153_v0Wen;
    logic         io_diffCommits_info_153_vlWen;
    logic [5:0]   io_diffCommits_info_154_ldest;
    logic [7:0]   io_diffCommits_info_154_pdest;
    logic         io_diffCommits_info_154_rfWen;
    logic         io_diffCommits_info_154_fpWen;
    logic         io_diffCommits_info_154_vecWen;
    logic         io_diffCommits_info_154_v0Wen;
    logic         io_diffCommits_info_154_vlWen;
    logic [5:0]   io_diffCommits_info_155_ldest;
    logic [7:0]   io_diffCommits_info_155_pdest;
    logic         io_diffCommits_info_155_rfWen;
    logic         io_diffCommits_info_155_fpWen;
    logic         io_diffCommits_info_155_vecWen;
    logic         io_diffCommits_info_155_v0Wen;
    logic         io_diffCommits_info_155_vlWen;
    logic [5:0]   io_diffCommits_info_156_ldest;
    logic [7:0]   io_diffCommits_info_156_pdest;
    logic         io_diffCommits_info_156_rfWen;
    logic         io_diffCommits_info_156_fpWen;
    logic         io_diffCommits_info_156_vecWen;
    logic         io_diffCommits_info_156_v0Wen;
    logic         io_diffCommits_info_156_vlWen;
    logic [5:0]   io_diffCommits_info_157_ldest;
    logic [7:0]   io_diffCommits_info_157_pdest;
    logic         io_diffCommits_info_157_rfWen;
    logic         io_diffCommits_info_157_fpWen;
    logic         io_diffCommits_info_157_vecWen;
    logic         io_diffCommits_info_157_v0Wen;
    logic         io_diffCommits_info_157_vlWen;
    logic [5:0]   io_diffCommits_info_158_ldest;
    logic [7:0]   io_diffCommits_info_158_pdest;
    logic         io_diffCommits_info_158_rfWen;
    logic         io_diffCommits_info_158_fpWen;
    logic         io_diffCommits_info_158_vecWen;
    logic         io_diffCommits_info_158_v0Wen;
    logic         io_diffCommits_info_158_vlWen;
    logic [5:0]   io_diffCommits_info_159_ldest;
    logic [7:0]   io_diffCommits_info_159_pdest;
    logic         io_diffCommits_info_159_rfWen;
    logic         io_diffCommits_info_159_fpWen;
    logic         io_diffCommits_info_159_vecWen;
    logic         io_diffCommits_info_159_v0Wen;
    logic         io_diffCommits_info_159_vlWen;
    logic [5:0]   io_diffCommits_info_160_ldest;
    logic [7:0]   io_diffCommits_info_160_pdest;
    logic         io_diffCommits_info_160_rfWen;
    logic         io_diffCommits_info_160_fpWen;
    logic         io_diffCommits_info_160_vecWen;
    logic         io_diffCommits_info_160_v0Wen;
    logic         io_diffCommits_info_160_vlWen;
    logic [5:0]   io_diffCommits_info_161_ldest;
    logic [7:0]   io_diffCommits_info_161_pdest;
    logic         io_diffCommits_info_161_rfWen;
    logic         io_diffCommits_info_161_fpWen;
    logic         io_diffCommits_info_161_vecWen;
    logic         io_diffCommits_info_161_v0Wen;
    logic         io_diffCommits_info_161_vlWen;
    logic [5:0]   io_diffCommits_info_162_ldest;
    logic [7:0]   io_diffCommits_info_162_pdest;
    logic         io_diffCommits_info_162_rfWen;
    logic         io_diffCommits_info_162_fpWen;
    logic         io_diffCommits_info_162_vecWen;
    logic         io_diffCommits_info_162_v0Wen;
    logic         io_diffCommits_info_162_vlWen;
    logic [5:0]   io_diffCommits_info_163_ldest;
    logic [7:0]   io_diffCommits_info_163_pdest;
    logic         io_diffCommits_info_163_rfWen;
    logic         io_diffCommits_info_163_fpWen;
    logic         io_diffCommits_info_163_vecWen;
    logic         io_diffCommits_info_163_v0Wen;
    logic         io_diffCommits_info_163_vlWen;
    logic [5:0]   io_diffCommits_info_164_ldest;
    logic [7:0]   io_diffCommits_info_164_pdest;
    logic         io_diffCommits_info_164_rfWen;
    logic         io_diffCommits_info_164_fpWen;
    logic         io_diffCommits_info_164_vecWen;
    logic         io_diffCommits_info_164_v0Wen;
    logic         io_diffCommits_info_164_vlWen;
    logic [5:0]   io_diffCommits_info_165_ldest;
    logic [7:0]   io_diffCommits_info_165_pdest;
    logic         io_diffCommits_info_165_rfWen;
    logic         io_diffCommits_info_165_fpWen;
    logic         io_diffCommits_info_165_vecWen;
    logic         io_diffCommits_info_165_v0Wen;
    logic         io_diffCommits_info_165_vlWen;
    logic [5:0]   io_diffCommits_info_166_ldest;
    logic [7:0]   io_diffCommits_info_166_pdest;
    logic         io_diffCommits_info_166_rfWen;
    logic         io_diffCommits_info_166_fpWen;
    logic         io_diffCommits_info_166_vecWen;
    logic         io_diffCommits_info_166_v0Wen;
    logic         io_diffCommits_info_166_vlWen;
    logic [5:0]   io_diffCommits_info_167_ldest;
    logic [7:0]   io_diffCommits_info_167_pdest;
    logic         io_diffCommits_info_167_rfWen;
    logic         io_diffCommits_info_167_fpWen;
    logic         io_diffCommits_info_167_vecWen;
    logic         io_diffCommits_info_167_v0Wen;
    logic         io_diffCommits_info_167_vlWen;
    logic [5:0]   io_diffCommits_info_168_ldest;
    logic [7:0]   io_diffCommits_info_168_pdest;
    logic         io_diffCommits_info_168_rfWen;
    logic         io_diffCommits_info_168_fpWen;
    logic         io_diffCommits_info_168_vecWen;
    logic         io_diffCommits_info_168_v0Wen;
    logic         io_diffCommits_info_168_vlWen;
    logic [5:0]   io_diffCommits_info_169_ldest;
    logic [7:0]   io_diffCommits_info_169_pdest;
    logic         io_diffCommits_info_169_rfWen;
    logic         io_diffCommits_info_169_fpWen;
    logic         io_diffCommits_info_169_vecWen;
    logic         io_diffCommits_info_169_v0Wen;
    logic         io_diffCommits_info_169_vlWen;
    logic [5:0]   io_diffCommits_info_170_ldest;
    logic [7:0]   io_diffCommits_info_170_pdest;
    logic         io_diffCommits_info_170_rfWen;
    logic         io_diffCommits_info_170_fpWen;
    logic         io_diffCommits_info_170_vecWen;
    logic         io_diffCommits_info_170_v0Wen;
    logic         io_diffCommits_info_170_vlWen;
    logic [5:0]   io_diffCommits_info_171_ldest;
    logic [7:0]   io_diffCommits_info_171_pdest;
    logic         io_diffCommits_info_171_rfWen;
    logic         io_diffCommits_info_171_fpWen;
    logic         io_diffCommits_info_171_vecWen;
    logic         io_diffCommits_info_171_v0Wen;
    logic         io_diffCommits_info_171_vlWen;
    logic [5:0]   io_diffCommits_info_172_ldest;
    logic [7:0]   io_diffCommits_info_172_pdest;
    logic         io_diffCommits_info_172_rfWen;
    logic         io_diffCommits_info_172_fpWen;
    logic         io_diffCommits_info_172_vecWen;
    logic         io_diffCommits_info_172_v0Wen;
    logic         io_diffCommits_info_172_vlWen;
    logic [5:0]   io_diffCommits_info_173_ldest;
    logic [7:0]   io_diffCommits_info_173_pdest;
    logic         io_diffCommits_info_173_rfWen;
    logic         io_diffCommits_info_173_fpWen;
    logic         io_diffCommits_info_173_vecWen;
    logic         io_diffCommits_info_173_v0Wen;
    logic         io_diffCommits_info_173_vlWen;
    logic [5:0]   io_diffCommits_info_174_ldest;
    logic [7:0]   io_diffCommits_info_174_pdest;
    logic         io_diffCommits_info_174_rfWen;
    logic         io_diffCommits_info_174_fpWen;
    logic         io_diffCommits_info_174_vecWen;
    logic         io_diffCommits_info_174_v0Wen;
    logic         io_diffCommits_info_174_vlWen;
    logic [5:0]   io_diffCommits_info_175_ldest;
    logic [7:0]   io_diffCommits_info_175_pdest;
    logic         io_diffCommits_info_175_rfWen;
    logic         io_diffCommits_info_175_fpWen;
    logic         io_diffCommits_info_175_vecWen;
    logic         io_diffCommits_info_175_v0Wen;
    logic         io_diffCommits_info_175_vlWen;
    logic [5:0]   io_diffCommits_info_176_ldest;
    logic [7:0]   io_diffCommits_info_176_pdest;
    logic         io_diffCommits_info_176_rfWen;
    logic         io_diffCommits_info_176_fpWen;
    logic         io_diffCommits_info_176_vecWen;
    logic         io_diffCommits_info_176_v0Wen;
    logic         io_diffCommits_info_176_vlWen;
    logic [5:0]   io_diffCommits_info_177_ldest;
    logic [7:0]   io_diffCommits_info_177_pdest;
    logic         io_diffCommits_info_177_rfWen;
    logic         io_diffCommits_info_177_fpWen;
    logic         io_diffCommits_info_177_vecWen;
    logic         io_diffCommits_info_177_v0Wen;
    logic         io_diffCommits_info_177_vlWen;
    logic [5:0]   io_diffCommits_info_178_ldest;
    logic [7:0]   io_diffCommits_info_178_pdest;
    logic         io_diffCommits_info_178_rfWen;
    logic         io_diffCommits_info_178_fpWen;
    logic         io_diffCommits_info_178_vecWen;
    logic         io_diffCommits_info_178_v0Wen;
    logic         io_diffCommits_info_178_vlWen;
    logic [5:0]   io_diffCommits_info_179_ldest;
    logic [7:0]   io_diffCommits_info_179_pdest;
    logic         io_diffCommits_info_179_rfWen;
    logic         io_diffCommits_info_179_fpWen;
    logic         io_diffCommits_info_179_vecWen;
    logic         io_diffCommits_info_179_v0Wen;
    logic         io_diffCommits_info_179_vlWen;
    logic [5:0]   io_diffCommits_info_180_ldest;
    logic [7:0]   io_diffCommits_info_180_pdest;
    logic         io_diffCommits_info_180_rfWen;
    logic         io_diffCommits_info_180_fpWen;
    logic         io_diffCommits_info_180_vecWen;
    logic         io_diffCommits_info_180_v0Wen;
    logic         io_diffCommits_info_180_vlWen;
    logic [5:0]   io_diffCommits_info_181_ldest;
    logic [7:0]   io_diffCommits_info_181_pdest;
    logic         io_diffCommits_info_181_rfWen;
    logic         io_diffCommits_info_181_fpWen;
    logic         io_diffCommits_info_181_vecWen;
    logic         io_diffCommits_info_181_v0Wen;
    logic         io_diffCommits_info_181_vlWen;
    logic [5:0]   io_diffCommits_info_182_ldest;
    logic [7:0]   io_diffCommits_info_182_pdest;
    logic         io_diffCommits_info_182_rfWen;
    logic         io_diffCommits_info_182_fpWen;
    logic         io_diffCommits_info_182_vecWen;
    logic         io_diffCommits_info_182_v0Wen;
    logic         io_diffCommits_info_182_vlWen;
    logic [5:0]   io_diffCommits_info_183_ldest;
    logic [7:0]   io_diffCommits_info_183_pdest;
    logic         io_diffCommits_info_183_rfWen;
    logic         io_diffCommits_info_183_fpWen;
    logic         io_diffCommits_info_183_vecWen;
    logic         io_diffCommits_info_183_v0Wen;
    logic         io_diffCommits_info_183_vlWen;
    logic [5:0]   io_diffCommits_info_184_ldest;
    logic [7:0]   io_diffCommits_info_184_pdest;
    logic         io_diffCommits_info_184_rfWen;
    logic         io_diffCommits_info_184_fpWen;
    logic         io_diffCommits_info_184_vecWen;
    logic         io_diffCommits_info_184_v0Wen;
    logic         io_diffCommits_info_184_vlWen;
    logic [5:0]   io_diffCommits_info_185_ldest;
    logic [7:0]   io_diffCommits_info_185_pdest;
    logic         io_diffCommits_info_185_rfWen;
    logic         io_diffCommits_info_185_fpWen;
    logic         io_diffCommits_info_185_vecWen;
    logic         io_diffCommits_info_185_v0Wen;
    logic         io_diffCommits_info_185_vlWen;
    logic [5:0]   io_diffCommits_info_186_ldest;
    logic [7:0]   io_diffCommits_info_186_pdest;
    logic         io_diffCommits_info_186_rfWen;
    logic         io_diffCommits_info_186_fpWen;
    logic         io_diffCommits_info_186_vecWen;
    logic         io_diffCommits_info_186_v0Wen;
    logic         io_diffCommits_info_186_vlWen;
    logic [5:0]   io_diffCommits_info_187_ldest;
    logic [7:0]   io_diffCommits_info_187_pdest;
    logic         io_diffCommits_info_187_rfWen;
    logic         io_diffCommits_info_187_fpWen;
    logic         io_diffCommits_info_187_vecWen;
    logic         io_diffCommits_info_187_v0Wen;
    logic         io_diffCommits_info_187_vlWen;
    logic [5:0]   io_diffCommits_info_188_ldest;
    logic [7:0]   io_diffCommits_info_188_pdest;
    logic         io_diffCommits_info_188_rfWen;
    logic         io_diffCommits_info_188_fpWen;
    logic         io_diffCommits_info_188_vecWen;
    logic         io_diffCommits_info_188_v0Wen;
    logic         io_diffCommits_info_188_vlWen;
    logic [5:0]   io_diffCommits_info_189_ldest;
    logic [7:0]   io_diffCommits_info_189_pdest;
    logic         io_diffCommits_info_189_rfWen;
    logic         io_diffCommits_info_189_fpWen;
    logic         io_diffCommits_info_189_vecWen;
    logic         io_diffCommits_info_189_v0Wen;
    logic         io_diffCommits_info_189_vlWen;
    logic [5:0]   io_diffCommits_info_190_ldest;
    logic [7:0]   io_diffCommits_info_190_pdest;
    logic         io_diffCommits_info_190_rfWen;
    logic         io_diffCommits_info_190_fpWen;
    logic         io_diffCommits_info_190_vecWen;
    logic         io_diffCommits_info_190_v0Wen;
    logic         io_diffCommits_info_190_vlWen;
    logic [5:0]   io_diffCommits_info_191_ldest;
    logic [7:0]   io_diffCommits_info_191_pdest;
    logic         io_diffCommits_info_191_rfWen;
    logic         io_diffCommits_info_191_fpWen;
    logic         io_diffCommits_info_191_vecWen;
    logic         io_diffCommits_info_191_v0Wen;
    logic         io_diffCommits_info_191_vlWen;
    logic [5:0]   io_diffCommits_info_192_ldest;
    logic [7:0]   io_diffCommits_info_192_pdest;
    logic         io_diffCommits_info_192_rfWen;
    logic         io_diffCommits_info_192_fpWen;
    logic         io_diffCommits_info_192_vecWen;
    logic         io_diffCommits_info_192_v0Wen;
    logic         io_diffCommits_info_192_vlWen;
    logic [5:0]   io_diffCommits_info_193_ldest;
    logic [7:0]   io_diffCommits_info_193_pdest;
    logic         io_diffCommits_info_193_rfWen;
    logic         io_diffCommits_info_193_fpWen;
    logic         io_diffCommits_info_193_vecWen;
    logic         io_diffCommits_info_193_v0Wen;
    logic         io_diffCommits_info_193_vlWen;
    logic [5:0]   io_diffCommits_info_194_ldest;
    logic [7:0]   io_diffCommits_info_194_pdest;
    logic         io_diffCommits_info_194_rfWen;
    logic         io_diffCommits_info_194_fpWen;
    logic         io_diffCommits_info_194_vecWen;
    logic         io_diffCommits_info_194_v0Wen;
    logic         io_diffCommits_info_194_vlWen;
    logic [5:0]   io_diffCommits_info_195_ldest;
    logic [7:0]   io_diffCommits_info_195_pdest;
    logic         io_diffCommits_info_195_rfWen;
    logic         io_diffCommits_info_195_fpWen;
    logic         io_diffCommits_info_195_vecWen;
    logic         io_diffCommits_info_195_v0Wen;
    logic         io_diffCommits_info_195_vlWen;
    logic [5:0]   io_diffCommits_info_196_ldest;
    logic [7:0]   io_diffCommits_info_196_pdest;
    logic         io_diffCommits_info_196_rfWen;
    logic         io_diffCommits_info_196_fpWen;
    logic         io_diffCommits_info_196_vecWen;
    logic         io_diffCommits_info_196_v0Wen;
    logic         io_diffCommits_info_196_vlWen;
    logic [5:0]   io_diffCommits_info_197_ldest;
    logic [7:0]   io_diffCommits_info_197_pdest;
    logic         io_diffCommits_info_197_rfWen;
    logic         io_diffCommits_info_197_fpWen;
    logic         io_diffCommits_info_197_vecWen;
    logic         io_diffCommits_info_197_v0Wen;
    logic         io_diffCommits_info_197_vlWen;
    logic [5:0]   io_diffCommits_info_198_ldest;
    logic [7:0]   io_diffCommits_info_198_pdest;
    logic         io_diffCommits_info_198_rfWen;
    logic         io_diffCommits_info_198_fpWen;
    logic         io_diffCommits_info_198_vecWen;
    logic         io_diffCommits_info_198_v0Wen;
    logic         io_diffCommits_info_198_vlWen;
    logic [5:0]   io_diffCommits_info_199_ldest;
    logic [7:0]   io_diffCommits_info_199_pdest;
    logic         io_diffCommits_info_199_rfWen;
    logic         io_diffCommits_info_199_fpWen;
    logic         io_diffCommits_info_199_vecWen;
    logic         io_diffCommits_info_199_v0Wen;
    logic         io_diffCommits_info_199_vlWen;
    logic [5:0]   io_diffCommits_info_200_ldest;
    logic [7:0]   io_diffCommits_info_200_pdest;
    logic         io_diffCommits_info_200_rfWen;
    logic         io_diffCommits_info_200_fpWen;
    logic         io_diffCommits_info_200_vecWen;
    logic         io_diffCommits_info_200_v0Wen;
    logic         io_diffCommits_info_200_vlWen;
    logic [5:0]   io_diffCommits_info_201_ldest;
    logic [7:0]   io_diffCommits_info_201_pdest;
    logic         io_diffCommits_info_201_rfWen;
    logic         io_diffCommits_info_201_fpWen;
    logic         io_diffCommits_info_201_vecWen;
    logic         io_diffCommits_info_201_v0Wen;
    logic         io_diffCommits_info_201_vlWen;
    logic [5:0]   io_diffCommits_info_202_ldest;
    logic [7:0]   io_diffCommits_info_202_pdest;
    logic         io_diffCommits_info_202_rfWen;
    logic         io_diffCommits_info_202_fpWen;
    logic         io_diffCommits_info_202_vecWen;
    logic         io_diffCommits_info_202_v0Wen;
    logic         io_diffCommits_info_202_vlWen;
    logic [5:0]   io_diffCommits_info_203_ldest;
    logic [7:0]   io_diffCommits_info_203_pdest;
    logic         io_diffCommits_info_203_rfWen;
    logic         io_diffCommits_info_203_fpWen;
    logic         io_diffCommits_info_203_vecWen;
    logic         io_diffCommits_info_203_v0Wen;
    logic         io_diffCommits_info_203_vlWen;
    logic [5:0]   io_diffCommits_info_204_ldest;
    logic [7:0]   io_diffCommits_info_204_pdest;
    logic         io_diffCommits_info_204_rfWen;
    logic         io_diffCommits_info_204_fpWen;
    logic         io_diffCommits_info_204_vecWen;
    logic         io_diffCommits_info_204_v0Wen;
    logic         io_diffCommits_info_204_vlWen;
    logic [5:0]   io_diffCommits_info_205_ldest;
    logic [7:0]   io_diffCommits_info_205_pdest;
    logic         io_diffCommits_info_205_rfWen;
    logic         io_diffCommits_info_205_fpWen;
    logic         io_diffCommits_info_205_vecWen;
    logic         io_diffCommits_info_205_v0Wen;
    logic         io_diffCommits_info_205_vlWen;
    logic [5:0]   io_diffCommits_info_206_ldest;
    logic [7:0]   io_diffCommits_info_206_pdest;
    logic         io_diffCommits_info_206_rfWen;
    logic         io_diffCommits_info_206_fpWen;
    logic         io_diffCommits_info_206_vecWen;
    logic         io_diffCommits_info_206_v0Wen;
    logic         io_diffCommits_info_206_vlWen;
    logic [5:0]   io_diffCommits_info_207_ldest;
    logic [7:0]   io_diffCommits_info_207_pdest;
    logic         io_diffCommits_info_207_rfWen;
    logic         io_diffCommits_info_207_fpWen;
    logic         io_diffCommits_info_207_vecWen;
    logic         io_diffCommits_info_207_v0Wen;
    logic         io_diffCommits_info_207_vlWen;
    logic [5:0]   io_diffCommits_info_208_ldest;
    logic [7:0]   io_diffCommits_info_208_pdest;
    logic         io_diffCommits_info_208_rfWen;
    logic         io_diffCommits_info_208_fpWen;
    logic         io_diffCommits_info_208_vecWen;
    logic         io_diffCommits_info_208_v0Wen;
    logic         io_diffCommits_info_208_vlWen;
    logic [5:0]   io_diffCommits_info_209_ldest;
    logic [7:0]   io_diffCommits_info_209_pdest;
    logic         io_diffCommits_info_209_rfWen;
    logic         io_diffCommits_info_209_fpWen;
    logic         io_diffCommits_info_209_vecWen;
    logic         io_diffCommits_info_209_v0Wen;
    logic         io_diffCommits_info_209_vlWen;
    logic [5:0]   io_diffCommits_info_210_ldest;
    logic [7:0]   io_diffCommits_info_210_pdest;
    logic         io_diffCommits_info_210_rfWen;
    logic         io_diffCommits_info_210_fpWen;
    logic         io_diffCommits_info_210_vecWen;
    logic         io_diffCommits_info_210_v0Wen;
    logic         io_diffCommits_info_210_vlWen;
    logic [5:0]   io_diffCommits_info_211_ldest;
    logic [7:0]   io_diffCommits_info_211_pdest;
    logic         io_diffCommits_info_211_rfWen;
    logic         io_diffCommits_info_211_fpWen;
    logic         io_diffCommits_info_211_vecWen;
    logic         io_diffCommits_info_211_v0Wen;
    logic         io_diffCommits_info_211_vlWen;
    logic [5:0]   io_diffCommits_info_212_ldest;
    logic [7:0]   io_diffCommits_info_212_pdest;
    logic         io_diffCommits_info_212_rfWen;
    logic         io_diffCommits_info_212_fpWen;
    logic         io_diffCommits_info_212_vecWen;
    logic         io_diffCommits_info_212_v0Wen;
    logic         io_diffCommits_info_212_vlWen;
    logic [5:0]   io_diffCommits_info_213_ldest;
    logic [7:0]   io_diffCommits_info_213_pdest;
    logic         io_diffCommits_info_213_rfWen;
    logic         io_diffCommits_info_213_fpWen;
    logic         io_diffCommits_info_213_vecWen;
    logic         io_diffCommits_info_213_v0Wen;
    logic         io_diffCommits_info_213_vlWen;
    logic [5:0]   io_diffCommits_info_214_ldest;
    logic [7:0]   io_diffCommits_info_214_pdest;
    logic         io_diffCommits_info_214_rfWen;
    logic         io_diffCommits_info_214_fpWen;
    logic         io_diffCommits_info_214_vecWen;
    logic         io_diffCommits_info_214_v0Wen;
    logic         io_diffCommits_info_214_vlWen;
    logic [5:0]   io_diffCommits_info_215_ldest;
    logic [7:0]   io_diffCommits_info_215_pdest;
    logic         io_diffCommits_info_215_rfWen;
    logic         io_diffCommits_info_215_fpWen;
    logic         io_diffCommits_info_215_vecWen;
    logic         io_diffCommits_info_215_v0Wen;
    logic         io_diffCommits_info_215_vlWen;
    logic [5:0]   io_diffCommits_info_216_ldest;
    logic [7:0]   io_diffCommits_info_216_pdest;
    logic         io_diffCommits_info_216_rfWen;
    logic         io_diffCommits_info_216_fpWen;
    logic         io_diffCommits_info_216_vecWen;
    logic         io_diffCommits_info_216_v0Wen;
    logic         io_diffCommits_info_216_vlWen;
    logic [5:0]   io_diffCommits_info_217_ldest;
    logic [7:0]   io_diffCommits_info_217_pdest;
    logic         io_diffCommits_info_217_rfWen;
    logic         io_diffCommits_info_217_fpWen;
    logic         io_diffCommits_info_217_vecWen;
    logic         io_diffCommits_info_217_v0Wen;
    logic         io_diffCommits_info_217_vlWen;
    logic [5:0]   io_diffCommits_info_218_ldest;
    logic [7:0]   io_diffCommits_info_218_pdest;
    logic         io_diffCommits_info_218_rfWen;
    logic         io_diffCommits_info_218_fpWen;
    logic         io_diffCommits_info_218_vecWen;
    logic         io_diffCommits_info_218_v0Wen;
    logic         io_diffCommits_info_218_vlWen;
    logic [5:0]   io_diffCommits_info_219_ldest;
    logic [7:0]   io_diffCommits_info_219_pdest;
    logic         io_diffCommits_info_219_rfWen;
    logic         io_diffCommits_info_219_fpWen;
    logic         io_diffCommits_info_219_vecWen;
    logic         io_diffCommits_info_219_v0Wen;
    logic         io_diffCommits_info_219_vlWen;
    logic [5:0]   io_diffCommits_info_220_ldest;
    logic [7:0]   io_diffCommits_info_220_pdest;
    logic         io_diffCommits_info_220_rfWen;
    logic         io_diffCommits_info_220_fpWen;
    logic         io_diffCommits_info_220_vecWen;
    logic         io_diffCommits_info_220_v0Wen;
    logic         io_diffCommits_info_220_vlWen;
    logic [5:0]   io_diffCommits_info_221_ldest;
    logic [7:0]   io_diffCommits_info_221_pdest;
    logic         io_diffCommits_info_221_rfWen;
    logic         io_diffCommits_info_221_fpWen;
    logic         io_diffCommits_info_221_vecWen;
    logic         io_diffCommits_info_221_v0Wen;
    logic         io_diffCommits_info_221_vlWen;
    logic [5:0]   io_diffCommits_info_222_ldest;
    logic [7:0]   io_diffCommits_info_222_pdest;
    logic         io_diffCommits_info_222_rfWen;
    logic         io_diffCommits_info_222_fpWen;
    logic         io_diffCommits_info_222_vecWen;
    logic         io_diffCommits_info_222_v0Wen;
    logic         io_diffCommits_info_222_vlWen;
    logic [5:0]   io_diffCommits_info_223_ldest;
    logic [7:0]   io_diffCommits_info_223_pdest;
    logic         io_diffCommits_info_223_rfWen;
    logic         io_diffCommits_info_223_fpWen;
    logic         io_diffCommits_info_223_vecWen;
    logic         io_diffCommits_info_223_v0Wen;
    logic         io_diffCommits_info_223_vlWen;
    logic [5:0]   io_diffCommits_info_224_ldest;
    logic [7:0]   io_diffCommits_info_224_pdest;
    logic         io_diffCommits_info_224_rfWen;
    logic         io_diffCommits_info_224_fpWen;
    logic         io_diffCommits_info_224_vecWen;
    logic         io_diffCommits_info_224_v0Wen;
    logic         io_diffCommits_info_224_vlWen;
    logic [5:0]   io_diffCommits_info_225_ldest;
    logic [7:0]   io_diffCommits_info_225_pdest;
    logic         io_diffCommits_info_225_rfWen;
    logic         io_diffCommits_info_225_fpWen;
    logic         io_diffCommits_info_225_vecWen;
    logic         io_diffCommits_info_225_v0Wen;
    logic         io_diffCommits_info_225_vlWen;
    logic [5:0]   io_diffCommits_info_226_ldest;
    logic [7:0]   io_diffCommits_info_226_pdest;
    logic         io_diffCommits_info_226_rfWen;
    logic         io_diffCommits_info_226_fpWen;
    logic         io_diffCommits_info_226_vecWen;
    logic         io_diffCommits_info_226_v0Wen;
    logic         io_diffCommits_info_226_vlWen;
    logic [5:0]   io_diffCommits_info_227_ldest;
    logic [7:0]   io_diffCommits_info_227_pdest;
    logic         io_diffCommits_info_227_rfWen;
    logic         io_diffCommits_info_227_fpWen;
    logic         io_diffCommits_info_227_vecWen;
    logic         io_diffCommits_info_227_v0Wen;
    logic         io_diffCommits_info_227_vlWen;
    logic [5:0]   io_diffCommits_info_228_ldest;
    logic [7:0]   io_diffCommits_info_228_pdest;
    logic         io_diffCommits_info_228_rfWen;
    logic         io_diffCommits_info_228_fpWen;
    logic         io_diffCommits_info_228_vecWen;
    logic         io_diffCommits_info_228_v0Wen;
    logic         io_diffCommits_info_228_vlWen;
    logic [5:0]   io_diffCommits_info_229_ldest;
    logic [7:0]   io_diffCommits_info_229_pdest;
    logic         io_diffCommits_info_229_rfWen;
    logic         io_diffCommits_info_229_fpWen;
    logic         io_diffCommits_info_229_vecWen;
    logic         io_diffCommits_info_229_v0Wen;
    logic         io_diffCommits_info_229_vlWen;
    logic [5:0]   io_diffCommits_info_230_ldest;
    logic [7:0]   io_diffCommits_info_230_pdest;
    logic         io_diffCommits_info_230_rfWen;
    logic         io_diffCommits_info_230_fpWen;
    logic         io_diffCommits_info_230_vecWen;
    logic         io_diffCommits_info_230_v0Wen;
    logic         io_diffCommits_info_230_vlWen;
    logic [5:0]   io_diffCommits_info_231_ldest;
    logic [7:0]   io_diffCommits_info_231_pdest;
    logic         io_diffCommits_info_231_rfWen;
    logic         io_diffCommits_info_231_fpWen;
    logic         io_diffCommits_info_231_vecWen;
    logic         io_diffCommits_info_231_v0Wen;
    logic         io_diffCommits_info_231_vlWen;
    logic [5:0]   io_diffCommits_info_232_ldest;
    logic [7:0]   io_diffCommits_info_232_pdest;
    logic         io_diffCommits_info_232_rfWen;
    logic         io_diffCommits_info_232_fpWen;
    logic         io_diffCommits_info_232_vecWen;
    logic         io_diffCommits_info_232_v0Wen;
    logic         io_diffCommits_info_232_vlWen;
    logic [5:0]   io_diffCommits_info_233_ldest;
    logic [7:0]   io_diffCommits_info_233_pdest;
    logic         io_diffCommits_info_233_rfWen;
    logic         io_diffCommits_info_233_fpWen;
    logic         io_diffCommits_info_233_vecWen;
    logic         io_diffCommits_info_233_v0Wen;
    logic         io_diffCommits_info_233_vlWen;
    logic [5:0]   io_diffCommits_info_234_ldest;
    logic [7:0]   io_diffCommits_info_234_pdest;
    logic         io_diffCommits_info_234_rfWen;
    logic         io_diffCommits_info_234_fpWen;
    logic         io_diffCommits_info_234_vecWen;
    logic         io_diffCommits_info_234_v0Wen;
    logic         io_diffCommits_info_234_vlWen;
    logic [5:0]   io_diffCommits_info_235_ldest;
    logic [7:0]   io_diffCommits_info_235_pdest;
    logic         io_diffCommits_info_235_rfWen;
    logic         io_diffCommits_info_235_fpWen;
    logic         io_diffCommits_info_235_vecWen;
    logic         io_diffCommits_info_235_v0Wen;
    logic         io_diffCommits_info_235_vlWen;
    logic [5:0]   io_diffCommits_info_236_ldest;
    logic [7:0]   io_diffCommits_info_236_pdest;
    logic         io_diffCommits_info_236_rfWen;
    logic         io_diffCommits_info_236_fpWen;
    logic         io_diffCommits_info_236_vecWen;
    logic         io_diffCommits_info_236_v0Wen;
    logic         io_diffCommits_info_236_vlWen;
    logic [5:0]   io_diffCommits_info_237_ldest;
    logic [7:0]   io_diffCommits_info_237_pdest;
    logic         io_diffCommits_info_237_rfWen;
    logic         io_diffCommits_info_237_fpWen;
    logic         io_diffCommits_info_237_vecWen;
    logic         io_diffCommits_info_237_v0Wen;
    logic         io_diffCommits_info_237_vlWen;
    logic [5:0]   io_diffCommits_info_238_ldest;
    logic [7:0]   io_diffCommits_info_238_pdest;
    logic         io_diffCommits_info_238_rfWen;
    logic         io_diffCommits_info_238_fpWen;
    logic         io_diffCommits_info_238_vecWen;
    logic         io_diffCommits_info_238_v0Wen;
    logic         io_diffCommits_info_238_vlWen;
    logic [5:0]   io_diffCommits_info_239_ldest;
    logic [7:0]   io_diffCommits_info_239_pdest;
    logic         io_diffCommits_info_239_rfWen;
    logic         io_diffCommits_info_239_fpWen;
    logic         io_diffCommits_info_239_vecWen;
    logic         io_diffCommits_info_239_v0Wen;
    logic         io_diffCommits_info_239_vlWen;
    logic [5:0]   io_diffCommits_info_240_ldest;
    logic [7:0]   io_diffCommits_info_240_pdest;
    logic         io_diffCommits_info_240_rfWen;
    logic         io_diffCommits_info_240_fpWen;
    logic         io_diffCommits_info_240_vecWen;
    logic         io_diffCommits_info_240_v0Wen;
    logic         io_diffCommits_info_240_vlWen;
    logic [5:0]   io_diffCommits_info_241_ldest;
    logic [7:0]   io_diffCommits_info_241_pdest;
    logic         io_diffCommits_info_241_rfWen;
    logic         io_diffCommits_info_241_fpWen;
    logic         io_diffCommits_info_241_vecWen;
    logic         io_diffCommits_info_241_v0Wen;
    logic         io_diffCommits_info_241_vlWen;
    logic [5:0]   io_diffCommits_info_242_ldest;
    logic [7:0]   io_diffCommits_info_242_pdest;
    logic         io_diffCommits_info_242_rfWen;
    logic         io_diffCommits_info_242_fpWen;
    logic         io_diffCommits_info_242_vecWen;
    logic         io_diffCommits_info_242_v0Wen;
    logic         io_diffCommits_info_242_vlWen;
    logic [5:0]   io_diffCommits_info_243_ldest;
    logic [7:0]   io_diffCommits_info_243_pdest;
    logic         io_diffCommits_info_243_rfWen;
    logic         io_diffCommits_info_243_fpWen;
    logic         io_diffCommits_info_243_vecWen;
    logic         io_diffCommits_info_243_v0Wen;
    logic         io_diffCommits_info_243_vlWen;
    logic [5:0]   io_diffCommits_info_244_ldest;
    logic [7:0]   io_diffCommits_info_244_pdest;
    logic         io_diffCommits_info_244_rfWen;
    logic         io_diffCommits_info_244_fpWen;
    logic         io_diffCommits_info_244_vecWen;
    logic         io_diffCommits_info_244_v0Wen;
    logic         io_diffCommits_info_244_vlWen;
    logic [5:0]   io_diffCommits_info_245_ldest;
    logic [7:0]   io_diffCommits_info_245_pdest;
    logic         io_diffCommits_info_245_rfWen;
    logic         io_diffCommits_info_245_fpWen;
    logic         io_diffCommits_info_245_vecWen;
    logic         io_diffCommits_info_245_v0Wen;
    logic         io_diffCommits_info_245_vlWen;
    logic [5:0]   io_diffCommits_info_246_ldest;
    logic [7:0]   io_diffCommits_info_246_pdest;
    logic         io_diffCommits_info_246_rfWen;
    logic         io_diffCommits_info_246_fpWen;
    logic         io_diffCommits_info_246_vecWen;
    logic         io_diffCommits_info_246_v0Wen;
    logic         io_diffCommits_info_246_vlWen;
    logic [5:0]   io_diffCommits_info_247_ldest;
    logic [7:0]   io_diffCommits_info_247_pdest;
    logic         io_diffCommits_info_247_rfWen;
    logic         io_diffCommits_info_247_fpWen;
    logic         io_diffCommits_info_247_vecWen;
    logic         io_diffCommits_info_247_v0Wen;
    logic         io_diffCommits_info_247_vlWen;
    logic [5:0]   io_diffCommits_info_248_ldest;
    logic [7:0]   io_diffCommits_info_248_pdest;
    logic         io_diffCommits_info_248_rfWen;
    logic         io_diffCommits_info_248_fpWen;
    logic         io_diffCommits_info_248_vecWen;
    logic         io_diffCommits_info_248_v0Wen;
    logic         io_diffCommits_info_248_vlWen;
    logic [5:0]   io_diffCommits_info_249_ldest;
    logic [7:0]   io_diffCommits_info_249_pdest;
    logic         io_diffCommits_info_249_rfWen;
    logic         io_diffCommits_info_249_fpWen;
    logic         io_diffCommits_info_249_vecWen;
    logic         io_diffCommits_info_249_v0Wen;
    logic         io_diffCommits_info_249_vlWen;
    logic [5:0]   io_diffCommits_info_250_ldest;
    logic [7:0]   io_diffCommits_info_250_pdest;
    logic         io_diffCommits_info_250_rfWen;
    logic         io_diffCommits_info_250_fpWen;
    logic         io_diffCommits_info_250_vecWen;
    logic         io_diffCommits_info_250_v0Wen;
    logic         io_diffCommits_info_250_vlWen;
    logic [5:0]   io_diffCommits_info_251_ldest;
    logic [7:0]   io_diffCommits_info_251_pdest;
    logic         io_diffCommits_info_251_rfWen;
    logic         io_diffCommits_info_251_fpWen;
    logic         io_diffCommits_info_251_vecWen;
    logic         io_diffCommits_info_251_v0Wen;
    logic         io_diffCommits_info_251_vlWen;
    logic [5:0]   io_diffCommits_info_252_ldest;
    logic [7:0]   io_diffCommits_info_252_pdest;
    logic         io_diffCommits_info_252_rfWen;
    logic         io_diffCommits_info_252_fpWen;
    logic         io_diffCommits_info_252_vecWen;
    logic         io_diffCommits_info_252_v0Wen;
    logic         io_diffCommits_info_252_vlWen;
    logic [5:0]   io_diffCommits_info_253_ldest;
    logic [7:0]   io_diffCommits_info_253_pdest;
    logic         io_diffCommits_info_253_rfWen;
    logic         io_diffCommits_info_253_fpWen;
    logic         io_diffCommits_info_253_vecWen;
    logic         io_diffCommits_info_253_v0Wen;
    logic         io_diffCommits_info_253_vlWen;
    logic [5:0]   io_diffCommits_info_254_ldest;
    logic [7:0]   io_diffCommits_info_254_pdest;
    logic         io_diffCommits_info_254_rfWen;
    logic         io_diffCommits_info_254_fpWen;
    logic         io_diffCommits_info_254_vecWen;
    logic         io_diffCommits_info_254_v0Wen;
    logic         io_diffCommits_info_254_vlWen;
    logic [5:0]   io_diffCommits_info_255_ldest;
    logic [7:0]   io_diffCommits_info_255_pdest;
    logic [5:0]   io_diffCommits_info_256_ldest;
    logic [7:0]   io_diffCommits_info_256_pdest;
    logic [5:0]   io_diffCommits_info_257_ldest;
    logic [7:0]   io_diffCommits_info_257_pdest;
    logic [5:0]   io_diffCommits_info_258_ldest;
    logic [7:0]   io_diffCommits_info_258_pdest;
    logic [5:0]   io_diffCommits_info_259_ldest;
    logic [7:0]   io_diffCommits_info_259_pdest;
    logic [5:0]   io_diffCommits_info_260_ldest;
    logic [7:0]   io_diffCommits_info_260_pdest;
    logic [5:0]   io_diffCommits_info_261_ldest;
    logic [7:0]   io_diffCommits_info_261_pdest;
    logic [5:0]   io_diffCommits_info_262_ldest;
    logic [7:0]   io_diffCommits_info_262_pdest;
    logic [5:0]   io_diffCommits_info_263_ldest;
    logic [7:0]   io_diffCommits_info_263_pdest;
    logic [5:0]   io_diffCommits_info_264_ldest;
    logic [7:0]   io_diffCommits_info_264_pdest;
    logic [5:0]   io_diffCommits_info_265_ldest;
    logic [7:0]   io_diffCommits_info_265_pdest;
    logic [5:0]   io_diffCommits_info_266_ldest;
    logic [7:0]   io_diffCommits_info_266_pdest;
    logic [5:0]   io_diffCommits_info_267_ldest;
    logic [7:0]   io_diffCommits_info_267_pdest;
    logic [5:0]   io_diffCommits_info_268_ldest;
    logic [7:0]   io_diffCommits_info_268_pdest;
    logic [5:0]   io_diffCommits_info_269_ldest;
    logic [7:0]   io_diffCommits_info_269_pdest;
    logic [5:0]   io_diffCommits_info_270_ldest;
    logic [7:0]   io_diffCommits_info_270_pdest;
    logic [5:0]   io_diffCommits_info_271_ldest;
    logic [7:0]   io_diffCommits_info_271_pdest;
    logic [5:0]   io_diffCommits_info_272_ldest;
    logic [7:0]   io_diffCommits_info_272_pdest;
    logic [5:0]   io_diffCommits_info_273_ldest;
    logic [7:0]   io_diffCommits_info_273_pdest;
    logic [5:0]   io_diffCommits_info_274_ldest;
    logic [7:0]   io_diffCommits_info_274_pdest;
    logic [5:0]   io_diffCommits_info_275_ldest;
    logic [7:0]   io_diffCommits_info_275_pdest;
    logic [5:0]   io_diffCommits_info_276_ldest;
    logic [7:0]   io_diffCommits_info_276_pdest;
    logic [5:0]   io_diffCommits_info_277_ldest;
    logic [7:0]   io_diffCommits_info_277_pdest;
    logic [5:0]   io_diffCommits_info_278_ldest;
    logic [7:0]   io_diffCommits_info_278_pdest;
    logic [5:0]   io_diffCommits_info_279_ldest;
    logic [7:0]   io_diffCommits_info_279_pdest;
    logic [5:0]   io_diffCommits_info_280_ldest;
    logic [7:0]   io_diffCommits_info_280_pdest;
    logic [5:0]   io_diffCommits_info_281_ldest;
    logic [7:0]   io_diffCommits_info_281_pdest;
    logic [5:0]   io_diffCommits_info_282_ldest;
    logic [7:0]   io_diffCommits_info_282_pdest;
    logic [5:0]   io_diffCommits_info_283_ldest;
    logic [7:0]   io_diffCommits_info_283_pdest;
    logic [5:0]   io_diffCommits_info_284_ldest;
    logic [7:0]   io_diffCommits_info_284_pdest;
    logic [5:0]   io_diffCommits_info_285_ldest;
    logic [7:0]   io_diffCommits_info_285_pdest;
    logic [5:0]   io_diffCommits_info_286_ldest;
    logic [7:0]   io_diffCommits_info_286_pdest;
    logic [5:0]   io_diffCommits_info_287_ldest;
    logic [7:0]   io_diffCommits_info_287_pdest;
    logic [5:0]   io_diffCommits_info_288_ldest;
    logic [7:0]   io_diffCommits_info_288_pdest;
    logic [5:0]   io_diffCommits_info_289_ldest;
    logic [7:0]   io_diffCommits_info_289_pdest;
    logic [5:0]   io_diffCommits_info_290_ldest;
    logic [7:0]   io_diffCommits_info_290_pdest;
    logic [5:0]   io_diffCommits_info_291_ldest;
    logic [7:0]   io_diffCommits_info_291_pdest;
    logic [5:0]   io_diffCommits_info_292_ldest;
    logic [7:0]   io_diffCommits_info_292_pdest;
    logic [5:0]   io_diffCommits_info_293_ldest;
    logic [7:0]   io_diffCommits_info_293_pdest;
    logic [5:0]   io_diffCommits_info_294_ldest;
    logic [7:0]   io_diffCommits_info_294_pdest;
    logic [5:0]   io_diffCommits_info_295_ldest;
    logic [7:0]   io_diffCommits_info_295_pdest;
    logic [5:0]   io_diffCommits_info_296_ldest;
    logic [7:0]   io_diffCommits_info_296_pdest;
    logic [5:0]   io_diffCommits_info_297_ldest;
    logic [7:0]   io_diffCommits_info_297_pdest;
    logic [5:0]   io_diffCommits_info_298_ldest;
    logic [7:0]   io_diffCommits_info_298_pdest;
    logic [5:0]   io_diffCommits_info_299_ldest;
    logic [7:0]   io_diffCommits_info_299_pdest;
    logic [5:0]   io_diffCommits_info_300_ldest;
    logic [7:0]   io_diffCommits_info_300_pdest;
    logic [5:0]   io_diffCommits_info_301_ldest;
    logic [7:0]   io_diffCommits_info_301_pdest;
    logic [5:0]   io_diffCommits_info_302_ldest;
    logic [7:0]   io_diffCommits_info_302_pdest;
    logic [5:0]   io_diffCommits_info_303_ldest;
    logic [7:0]   io_diffCommits_info_303_pdest;
    logic [5:0]   io_diffCommits_info_304_ldest;
    logic [7:0]   io_diffCommits_info_304_pdest;
    logic [5:0]   io_diffCommits_info_305_ldest;
    logic [7:0]   io_diffCommits_info_305_pdest;
    logic [5:0]   io_diffCommits_info_306_ldest;
    logic [7:0]   io_diffCommits_info_306_pdest;
    logic [5:0]   io_diffCommits_info_307_ldest;
    logic [7:0]   io_diffCommits_info_307_pdest;
    logic [5:0]   io_diffCommits_info_308_ldest;
    logic [7:0]   io_diffCommits_info_308_pdest;
    logic [5:0]   io_diffCommits_info_309_ldest;
    logic [7:0]   io_diffCommits_info_309_pdest;
    logic [5:0]   io_diffCommits_info_310_ldest;
    logic [7:0]   io_diffCommits_info_310_pdest;
    logic [5:0]   io_diffCommits_info_311_ldest;
    logic [7:0]   io_diffCommits_info_311_pdest;
    logic [5:0]   io_diffCommits_info_312_ldest;
    logic [7:0]   io_diffCommits_info_312_pdest;
    logic [5:0]   io_diffCommits_info_313_ldest;
    logic [7:0]   io_diffCommits_info_313_pdest;
    logic [5:0]   io_diffCommits_info_314_ldest;
    logic [7:0]   io_diffCommits_info_314_pdest;
    logic [5:0]   io_diffCommits_info_315_ldest;
    logic [7:0]   io_diffCommits_info_315_pdest;
    logic [5:0]   io_diffCommits_info_316_ldest;
    logic [7:0]   io_diffCommits_info_316_pdest;
    logic [5:0]   io_diffCommits_info_317_ldest;
    logic [7:0]   io_diffCommits_info_317_pdest;
    logic [5:0]   io_diffCommits_info_318_ldest;
    logic [7:0]   io_diffCommits_info_318_pdest;
    logic [5:0]   io_diffCommits_info_319_ldest;
    logic [7:0]   io_diffCommits_info_319_pdest;
    logic [5:0]   io_diffCommits_info_320_ldest;
    logic [7:0]   io_diffCommits_info_320_pdest;
    logic [5:0]   io_diffCommits_info_321_ldest;
    logic [7:0]   io_diffCommits_info_321_pdest;
    logic [5:0]   io_diffCommits_info_322_ldest;
    logic [7:0]   io_diffCommits_info_322_pdest;
    logic [5:0]   io_diffCommits_info_323_ldest;
    logic [7:0]   io_diffCommits_info_323_pdest;
    logic [5:0]   io_diffCommits_info_324_ldest;
    logic [7:0]   io_diffCommits_info_324_pdest;
    logic [5:0]   io_diffCommits_info_325_ldest;
    logic [7:0]   io_diffCommits_info_325_pdest;
    logic [5:0]   io_diffCommits_info_326_ldest;
    logic [7:0]   io_diffCommits_info_326_pdest;
    logic [5:0]   io_diffCommits_info_327_ldest;
    logic [7:0]   io_diffCommits_info_327_pdest;
    logic [5:0]   io_diffCommits_info_328_ldest;
    logic [7:0]   io_diffCommits_info_328_pdest;
    logic [5:0]   io_diffCommits_info_329_ldest;
    logic [7:0]   io_diffCommits_info_329_pdest;
    logic [5:0]   io_diffCommits_info_330_ldest;
    logic [7:0]   io_diffCommits_info_330_pdest;
    logic [5:0]   io_diffCommits_info_331_ldest;
    logic [7:0]   io_diffCommits_info_331_pdest;
    logic [5:0]   io_diffCommits_info_332_ldest;
    logic [7:0]   io_diffCommits_info_332_pdest;
    logic [5:0]   io_diffCommits_info_333_ldest;
    logic [7:0]   io_diffCommits_info_333_pdest;
    logic [5:0]   io_diffCommits_info_334_ldest;
    logic [7:0]   io_diffCommits_info_334_pdest;
    logic [5:0]   io_diffCommits_info_335_ldest;
    logic [7:0]   io_diffCommits_info_335_pdest;
    logic [5:0]   io_diffCommits_info_336_ldest;
    logic [7:0]   io_diffCommits_info_336_pdest;
    logic [5:0]   io_diffCommits_info_337_ldest;
    logic [7:0]   io_diffCommits_info_337_pdest;
    logic [5:0]   io_diffCommits_info_338_ldest;
    logic [7:0]   io_diffCommits_info_338_pdest;
    logic [5:0]   io_diffCommits_info_339_ldest;
    logic [7:0]   io_diffCommits_info_339_pdest;
    logic [5:0]   io_diffCommits_info_340_ldest;
    logic [7:0]   io_diffCommits_info_340_pdest;
    logic [5:0]   io_diffCommits_info_341_ldest;
    logic [7:0]   io_diffCommits_info_341_pdest;
    logic [5:0]   io_diffCommits_info_342_ldest;
    logic [7:0]   io_diffCommits_info_342_pdest;
    logic [5:0]   io_diffCommits_info_343_ldest;
    logic [7:0]   io_diffCommits_info_343_pdest;
    logic [5:0]   io_diffCommits_info_344_ldest;
    logic [7:0]   io_diffCommits_info_344_pdest;
    logic [5:0]   io_diffCommits_info_345_ldest;
    logic [7:0]   io_diffCommits_info_345_pdest;
    logic [5:0]   io_diffCommits_info_346_ldest;
    logic [7:0]   io_diffCommits_info_346_pdest;
    logic [5:0]   io_diffCommits_info_347_ldest;
    logic [7:0]   io_diffCommits_info_347_pdest;
    logic [5:0]   io_diffCommits_info_348_ldest;
    logic [7:0]   io_diffCommits_info_348_pdest;
    logic [5:0]   io_diffCommits_info_349_ldest;
    logic [7:0]   io_diffCommits_info_349_pdest;
    logic [5:0]   io_diffCommits_info_350_ldest;
    logic [7:0]   io_diffCommits_info_350_pdest;
    logic [5:0]   io_diffCommits_info_351_ldest;
    logic [7:0]   io_diffCommits_info_351_pdest;
    logic [5:0]   io_diffCommits_info_352_ldest;
    logic [7:0]   io_diffCommits_info_352_pdest;
    logic [5:0]   io_diffCommits_info_353_ldest;
    logic [7:0]   io_diffCommits_info_353_pdest;
    logic [5:0]   io_diffCommits_info_354_ldest;
    logic [7:0]   io_diffCommits_info_354_pdest;
    logic [5:0]   io_diffCommits_info_355_ldest;
    logic [7:0]   io_diffCommits_info_355_pdest;
    logic [5:0]   io_diffCommits_info_356_ldest;
    logic [7:0]   io_diffCommits_info_356_pdest;
    logic [5:0]   io_diffCommits_info_357_ldest;
    logic [7:0]   io_diffCommits_info_357_pdest;
    logic [5:0]   io_diffCommits_info_358_ldest;
    logic [7:0]   io_diffCommits_info_358_pdest;
    logic [5:0]   io_diffCommits_info_359_ldest;
    logic [7:0]   io_diffCommits_info_359_pdest;
    logic [5:0]   io_diffCommits_info_360_ldest;
    logic [7:0]   io_diffCommits_info_360_pdest;
    logic [5:0]   io_diffCommits_info_361_ldest;
    logic [7:0]   io_diffCommits_info_361_pdest;
    logic [5:0]   io_diffCommits_info_362_ldest;
    logic [7:0]   io_diffCommits_info_362_pdest;
    logic [5:0]   io_diffCommits_info_363_ldest;
    logic [7:0]   io_diffCommits_info_363_pdest;
    logic [5:0]   io_diffCommits_info_364_ldest;
    logic [7:0]   io_diffCommits_info_364_pdest;
    logic [5:0]   io_diffCommits_info_365_ldest;
    logic [7:0]   io_diffCommits_info_365_pdest;
    logic [5:0]   io_diffCommits_info_366_ldest;
    logic [7:0]   io_diffCommits_info_366_pdest;
    logic [5:0]   io_diffCommits_info_367_ldest;
    logic [7:0]   io_diffCommits_info_367_pdest;
    logic [5:0]   io_diffCommits_info_368_ldest;
    logic [7:0]   io_diffCommits_info_368_pdest;
    logic [5:0]   io_diffCommits_info_369_ldest;
    logic [7:0]   io_diffCommits_info_369_pdest;
    logic [5:0]   io_diffCommits_info_370_ldest;
    logic [7:0]   io_diffCommits_info_370_pdest;
    logic [5:0]   io_diffCommits_info_371_ldest;
    logic [7:0]   io_diffCommits_info_371_pdest;
    logic [5:0]   io_diffCommits_info_372_ldest;
    logic [7:0]   io_diffCommits_info_372_pdest;
    logic [5:0]   io_diffCommits_info_373_ldest;
    logic [7:0]   io_diffCommits_info_373_pdest;
    logic [5:0]   io_diffCommits_info_374_ldest;
    logic [7:0]   io_diffCommits_info_374_pdest;
    logic [5:0]   io_diffCommits_info_375_ldest;
    logic [7:0]   io_diffCommits_info_375_pdest;
    logic [5:0]   io_diffCommits_info_376_ldest;
    logic [7:0]   io_diffCommits_info_376_pdest;
    logic [5:0]   io_diffCommits_info_377_ldest;
    logic [7:0]   io_diffCommits_info_377_pdest;
    logic [5:0]   io_diffCommits_info_378_ldest;
    logic [7:0]   io_diffCommits_info_378_pdest;
    logic [5:0]   io_diffCommits_info_379_ldest;
    logic [7:0]   io_diffCommits_info_379_pdest;
    logic [5:0]   io_diffCommits_info_380_ldest;
    logic [7:0]   io_diffCommits_info_380_pdest;
    logic [5:0]   io_diffCommits_info_381_ldest;
    logic [7:0]   io_diffCommits_info_381_pdest;
    logic [5:0]   io_diffCommits_info_382_ldest;
    logic [7:0]   io_diffCommits_info_382_pdest;
    logic [5:0]   io_diffCommits_info_383_ldest;
    logic [7:0]   io_diffCommits_info_383_pdest;
    logic [5:0]   io_diffCommits_info_384_ldest;
    logic [7:0]   io_diffCommits_info_384_pdest;
    logic [5:0]   io_diffCommits_info_385_ldest;
    logic [7:0]   io_diffCommits_info_385_pdest;
    logic [5:0]   io_diffCommits_info_386_ldest;
    logic [7:0]   io_diffCommits_info_386_pdest;
    logic [5:0]   io_diffCommits_info_387_ldest;
    logic [7:0]   io_diffCommits_info_387_pdest;
    logic [5:0]   io_diffCommits_info_388_ldest;
    logic [7:0]   io_diffCommits_info_388_pdest;
    logic [5:0]   io_diffCommits_info_389_ldest;
    logic [7:0]   io_diffCommits_info_389_pdest;
    logic [3:0]   io_lsq_scommit       ;
    logic         io_lsq_pendingMMIOld ;
    logic         io_lsq_pendingst     ;
    logic         io_lsq_pendingPtr_flag;
    logic [7:0]   io_lsq_pendingPtr_value;
    logic         io_robDeqPtr_flag    ;
    logic [7:0]   io_robDeqPtr_value   ;
    logic         io_csr_fflags_valid  ;
    logic [4:0]   io_csr_fflags_bits   ;
    logic         io_csr_vxsat_valid   ;
    logic         io_csr_vxsat_bits    ;
    logic         io_csr_vstart_valid  ;
    logic [63:0]  io_csr_vstart_bits   ;
    logic         io_csr_dirty_fs      ;
    logic         io_csr_dirty_vs      ;
    logic [6:0]   io_csr_perfinfo_retiredInstr;
    logic         io_cpu_halt          ;
    logic         io_wfi_wfiReq        ;
    logic         io_toDecode_isResumeVType;
    logic         io_toDecode_walkToArchVType;
    logic         io_toDecode_walkVType_valid;
    logic         io_toDecode_walkVType_bits_illegal;
    logic         io_toDecode_walkVType_bits_vma;
    logic         io_toDecode_walkVType_bits_vta;
    logic [1:0]   io_toDecode_walkVType_bits_vsew;
    logic [2:0]   io_toDecode_walkVType_bits_vlmul;
    logic         io_toDecode_commitVType_vtype_valid;
    logic         io_toDecode_commitVType_vtype_bits_illegal;
    logic         io_toDecode_commitVType_vtype_bits_vma;
    logic         io_toDecode_commitVType_vtype_bits_vta;
    logic [1:0]   io_toDecode_commitVType_vtype_bits_vsew;
    logic [2:0]   io_toDecode_commitVType_vtype_bits_vlmul;
    logic         io_toDecode_commitVType_hasVsetvl;
    logic         io_readGPAMemAddr_valid;
    logic [5:0]   io_readGPAMemAddr_bits_ftqPtr_value;
    logic [3:0]   io_readGPAMemAddr_bits_ftqOffset;
    logic         io_toVecExcpMod_logicPhyRegMap_0_valid;
    logic [5:0]   io_toVecExcpMod_logicPhyRegMap_0_bits_lreg;
    logic [6:0]   io_toVecExcpMod_logicPhyRegMap_0_bits_preg;
    logic         io_toVecExcpMod_logicPhyRegMap_1_valid;
    logic [5:0]   io_toVecExcpMod_logicPhyRegMap_1_bits_lreg;
    logic [6:0]   io_toVecExcpMod_logicPhyRegMap_1_bits_preg;
    logic         io_toVecExcpMod_logicPhyRegMap_2_valid;
    logic [5:0]   io_toVecExcpMod_logicPhyRegMap_2_bits_lreg;
    logic [6:0]   io_toVecExcpMod_logicPhyRegMap_2_bits_preg;
    logic         io_toVecExcpMod_logicPhyRegMap_3_valid;
    logic [5:0]   io_toVecExcpMod_logicPhyRegMap_3_bits_lreg;
    logic [6:0]   io_toVecExcpMod_logicPhyRegMap_3_bits_preg;
    logic         io_toVecExcpMod_logicPhyRegMap_4_valid;
    logic [5:0]   io_toVecExcpMod_logicPhyRegMap_4_bits_lreg;
    logic [6:0]   io_toVecExcpMod_logicPhyRegMap_4_bits_preg;
    logic         io_toVecExcpMod_logicPhyRegMap_5_valid;
    logic [5:0]   io_toVecExcpMod_logicPhyRegMap_5_bits_lreg;
    logic [6:0]   io_toVecExcpMod_logicPhyRegMap_5_bits_preg;
    logic         io_toVecExcpMod_excpInfo_valid;
    logic [6:0]   io_toVecExcpMod_excpInfo_bits_vstart;
    logic [1:0]   io_toVecExcpMod_excpInfo_bits_vsew;
    logic [1:0]   io_toVecExcpMod_excpInfo_bits_veew;
    logic [2:0]   io_toVecExcpMod_excpInfo_bits_vlmul;
    logic [2:0]   io_toVecExcpMod_excpInfo_bits_nf;
    logic         io_toVecExcpMod_excpInfo_bits_isStride;
    logic         io_toVecExcpMod_excpInfo_bits_isIndexed;
    logic         io_toVecExcpMod_excpInfo_bits_isWhole;
    logic         io_toVecExcpMod_excpInfo_bits_isVlm;
    logic [49:0]  io_storeDebugInfo_1_pc;
    logic [5:0]   io_perf_0_value      ;
    logic [5:0]   io_perf_1_value      ;
    logic [5:0]   io_perf_2_value      ;
    logic [5:0]   io_perf_3_value      ;
    logic [5:0]   io_perf_4_value      ;
    logic [5:0]   io_perf_5_value      ;
    logic [5:0]   io_perf_6_value      ;
    logic [5:0]   io_perf_7_value      ;
    logic [5:0]   io_perf_8_value      ;
    logic [5:0]   io_perf_9_value      ;
    logic [5:0]   io_perf_10_value     ;
    logic [5:0]   io_perf_11_value     ;
    logic [5:0]   io_perf_12_value     ;
    logic [5:0]   io_perf_13_value     ;
    logic [5:0]   io_perf_14_value     ;
    logic [5:0]   io_perf_15_value     ;
    logic [5:0]   io_perf_16_value     ;
    logic [5:0]   io_perf_17_value     ;
    logic         io_error_0           ;

    Rob_output_agent_xaction  mon_tr;
    while(1) begin
        @this.vif.mon_mp.mon_cb;
        io_enq_canAccept = this.vif.mon_mp.mon_cb.io_enq_canAccept;
        io_enq_canAcceptForDispatch = this.vif.mon_mp.mon_cb.io_enq_canAcceptForDispatch;
        io_enq_isEmpty = this.vif.mon_mp.mon_cb.io_enq_isEmpty;
        io_flushOut_valid = this.vif.mon_mp.mon_cb.io_flushOut_valid;
        io_flushOut_bits_isRVC = this.vif.mon_mp.mon_cb.io_flushOut_bits_isRVC;
        io_flushOut_bits_robIdx_flag = this.vif.mon_mp.mon_cb.io_flushOut_bits_robIdx_flag;
        io_flushOut_bits_robIdx_value = this.vif.mon_mp.mon_cb.io_flushOut_bits_robIdx_value;
        io_flushOut_bits_ftqIdx_flag = this.vif.mon_mp.mon_cb.io_flushOut_bits_ftqIdx_flag;
        io_flushOut_bits_ftqIdx_value = this.vif.mon_mp.mon_cb.io_flushOut_bits_ftqIdx_value;
        io_flushOut_bits_ftqOffset = this.vif.mon_mp.mon_cb.io_flushOut_bits_ftqOffset;
        io_flushOut_bits_level = this.vif.mon_mp.mon_cb.io_flushOut_bits_level;
        io_exception_valid = this.vif.mon_mp.mon_cb.io_exception_valid;
        io_exception_bits_instr = this.vif.mon_mp.mon_cb.io_exception_bits_instr;
        io_exception_bits_commitType = this.vif.mon_mp.mon_cb.io_exception_bits_commitType;
        io_exception_bits_exceptionVec_0 = this.vif.mon_mp.mon_cb.io_exception_bits_exceptionVec_0;
        io_exception_bits_exceptionVec_1 = this.vif.mon_mp.mon_cb.io_exception_bits_exceptionVec_1;
        io_exception_bits_exceptionVec_2 = this.vif.mon_mp.mon_cb.io_exception_bits_exceptionVec_2;
        io_exception_bits_exceptionVec_3 = this.vif.mon_mp.mon_cb.io_exception_bits_exceptionVec_3;
        io_exception_bits_exceptionVec_4 = this.vif.mon_mp.mon_cb.io_exception_bits_exceptionVec_4;
        io_exception_bits_exceptionVec_5 = this.vif.mon_mp.mon_cb.io_exception_bits_exceptionVec_5;
        io_exception_bits_exceptionVec_6 = this.vif.mon_mp.mon_cb.io_exception_bits_exceptionVec_6;
        io_exception_bits_exceptionVec_7 = this.vif.mon_mp.mon_cb.io_exception_bits_exceptionVec_7;
        io_exception_bits_exceptionVec_8 = this.vif.mon_mp.mon_cb.io_exception_bits_exceptionVec_8;
        io_exception_bits_exceptionVec_9 = this.vif.mon_mp.mon_cb.io_exception_bits_exceptionVec_9;
        io_exception_bits_exceptionVec_10 = this.vif.mon_mp.mon_cb.io_exception_bits_exceptionVec_10;
        io_exception_bits_exceptionVec_11 = this.vif.mon_mp.mon_cb.io_exception_bits_exceptionVec_11;
        io_exception_bits_exceptionVec_12 = this.vif.mon_mp.mon_cb.io_exception_bits_exceptionVec_12;
        io_exception_bits_exceptionVec_13 = this.vif.mon_mp.mon_cb.io_exception_bits_exceptionVec_13;
        io_exception_bits_exceptionVec_14 = this.vif.mon_mp.mon_cb.io_exception_bits_exceptionVec_14;
        io_exception_bits_exceptionVec_15 = this.vif.mon_mp.mon_cb.io_exception_bits_exceptionVec_15;
        io_exception_bits_exceptionVec_16 = this.vif.mon_mp.mon_cb.io_exception_bits_exceptionVec_16;
        io_exception_bits_exceptionVec_17 = this.vif.mon_mp.mon_cb.io_exception_bits_exceptionVec_17;
        io_exception_bits_exceptionVec_18 = this.vif.mon_mp.mon_cb.io_exception_bits_exceptionVec_18;
        io_exception_bits_exceptionVec_19 = this.vif.mon_mp.mon_cb.io_exception_bits_exceptionVec_19;
        io_exception_bits_exceptionVec_20 = this.vif.mon_mp.mon_cb.io_exception_bits_exceptionVec_20;
        io_exception_bits_exceptionVec_21 = this.vif.mon_mp.mon_cb.io_exception_bits_exceptionVec_21;
        io_exception_bits_exceptionVec_22 = this.vif.mon_mp.mon_cb.io_exception_bits_exceptionVec_22;
        io_exception_bits_exceptionVec_23 = this.vif.mon_mp.mon_cb.io_exception_bits_exceptionVec_23;
        io_exception_bits_isPcBkpt = this.vif.mon_mp.mon_cb.io_exception_bits_isPcBkpt;
        io_exception_bits_isFetchMalAddr = this.vif.mon_mp.mon_cb.io_exception_bits_isFetchMalAddr;
        io_exception_bits_gpaddr = this.vif.mon_mp.mon_cb.io_exception_bits_gpaddr;
        io_exception_bits_singleStep = this.vif.mon_mp.mon_cb.io_exception_bits_singleStep;
        io_exception_bits_crossPageIPFFix = this.vif.mon_mp.mon_cb.io_exception_bits_crossPageIPFFix;
        io_exception_bits_isInterrupt = this.vif.mon_mp.mon_cb.io_exception_bits_isInterrupt;
        io_exception_bits_isHls = this.vif.mon_mp.mon_cb.io_exception_bits_isHls;
        io_exception_bits_trigger = this.vif.mon_mp.mon_cb.io_exception_bits_trigger;
        io_exception_bits_isForVSnonLeafPTE = this.vif.mon_mp.mon_cb.io_exception_bits_isForVSnonLeafPTE;
        io_commits_isCommit = this.vif.mon_mp.mon_cb.io_commits_isCommit;
        io_commits_commitValid_0 = this.vif.mon_mp.mon_cb.io_commits_commitValid_0;
        io_commits_commitValid_1 = this.vif.mon_mp.mon_cb.io_commits_commitValid_1;
        io_commits_commitValid_2 = this.vif.mon_mp.mon_cb.io_commits_commitValid_2;
        io_commits_commitValid_3 = this.vif.mon_mp.mon_cb.io_commits_commitValid_3;
        io_commits_commitValid_4 = this.vif.mon_mp.mon_cb.io_commits_commitValid_4;
        io_commits_commitValid_5 = this.vif.mon_mp.mon_cb.io_commits_commitValid_5;
        io_commits_commitValid_6 = this.vif.mon_mp.mon_cb.io_commits_commitValid_6;
        io_commits_commitValid_7 = this.vif.mon_mp.mon_cb.io_commits_commitValid_7;
        io_commits_isWalk = this.vif.mon_mp.mon_cb.io_commits_isWalk;
        io_commits_walkValid_0 = this.vif.mon_mp.mon_cb.io_commits_walkValid_0;
        io_commits_walkValid_1 = this.vif.mon_mp.mon_cb.io_commits_walkValid_1;
        io_commits_walkValid_2 = this.vif.mon_mp.mon_cb.io_commits_walkValid_2;
        io_commits_walkValid_3 = this.vif.mon_mp.mon_cb.io_commits_walkValid_3;
        io_commits_walkValid_4 = this.vif.mon_mp.mon_cb.io_commits_walkValid_4;
        io_commits_walkValid_5 = this.vif.mon_mp.mon_cb.io_commits_walkValid_5;
        io_commits_walkValid_6 = this.vif.mon_mp.mon_cb.io_commits_walkValid_6;
        io_commits_walkValid_7 = this.vif.mon_mp.mon_cb.io_commits_walkValid_7;
        io_commits_info_0_walk_v = this.vif.mon_mp.mon_cb.io_commits_info_0_walk_v;
        io_commits_info_0_commit_v = this.vif.mon_mp.mon_cb.io_commits_info_0_commit_v;
        io_commits_info_0_commit_w = this.vif.mon_mp.mon_cb.io_commits_info_0_commit_w;
        io_commits_info_0_realDestSize = this.vif.mon_mp.mon_cb.io_commits_info_0_realDestSize;
        io_commits_info_0_interrupt_safe = this.vif.mon_mp.mon_cb.io_commits_info_0_interrupt_safe;
        io_commits_info_0_wflags = this.vif.mon_mp.mon_cb.io_commits_info_0_wflags;
        io_commits_info_0_fflags = this.vif.mon_mp.mon_cb.io_commits_info_0_fflags;
        io_commits_info_0_vxsat = this.vif.mon_mp.mon_cb.io_commits_info_0_vxsat;
        io_commits_info_0_isRVC = this.vif.mon_mp.mon_cb.io_commits_info_0_isRVC;
        io_commits_info_0_isVset = this.vif.mon_mp.mon_cb.io_commits_info_0_isVset;
        io_commits_info_0_isHls = this.vif.mon_mp.mon_cb.io_commits_info_0_isHls;
        io_commits_info_0_isVls = this.vif.mon_mp.mon_cb.io_commits_info_0_isVls;
        io_commits_info_0_vls = this.vif.mon_mp.mon_cb.io_commits_info_0_vls;
        io_commits_info_0_mmio = this.vif.mon_mp.mon_cb.io_commits_info_0_mmio;
        io_commits_info_0_commitType = this.vif.mon_mp.mon_cb.io_commits_info_0_commitType;
        io_commits_info_0_ftqIdx_flag = this.vif.mon_mp.mon_cb.io_commits_info_0_ftqIdx_flag;
        io_commits_info_0_ftqIdx_value = this.vif.mon_mp.mon_cb.io_commits_info_0_ftqIdx_value;
        io_commits_info_0_ftqOffset = this.vif.mon_mp.mon_cb.io_commits_info_0_ftqOffset;
        io_commits_info_0_instrSize = this.vif.mon_mp.mon_cb.io_commits_info_0_instrSize;
        io_commits_info_0_fpWen = this.vif.mon_mp.mon_cb.io_commits_info_0_fpWen;
        io_commits_info_0_rfWen = this.vif.mon_mp.mon_cb.io_commits_info_0_rfWen;
        io_commits_info_0_needFlush = this.vif.mon_mp.mon_cb.io_commits_info_0_needFlush;
        io_commits_info_0_traceBlockInPipe_itype = this.vif.mon_mp.mon_cb.io_commits_info_0_traceBlockInPipe_itype;
        io_commits_info_0_traceBlockInPipe_iretire = this.vif.mon_mp.mon_cb.io_commits_info_0_traceBlockInPipe_iretire;
        io_commits_info_0_traceBlockInPipe_ilastsize = this.vif.mon_mp.mon_cb.io_commits_info_0_traceBlockInPipe_ilastsize;
        io_commits_info_0_debug_pc = this.vif.mon_mp.mon_cb.io_commits_info_0_debug_pc;
        io_commits_info_0_debug_instr = this.vif.mon_mp.mon_cb.io_commits_info_0_debug_instr;
        io_commits_info_0_debug_ldest = this.vif.mon_mp.mon_cb.io_commits_info_0_debug_ldest;
        io_commits_info_0_debug_pdest = this.vif.mon_mp.mon_cb.io_commits_info_0_debug_pdest;
        io_commits_info_0_debug_otherPdest_0 = this.vif.mon_mp.mon_cb.io_commits_info_0_debug_otherPdest_0;
        io_commits_info_0_debug_otherPdest_1 = this.vif.mon_mp.mon_cb.io_commits_info_0_debug_otherPdest_1;
        io_commits_info_0_debug_otherPdest_2 = this.vif.mon_mp.mon_cb.io_commits_info_0_debug_otherPdest_2;
        io_commits_info_0_debug_otherPdest_3 = this.vif.mon_mp.mon_cb.io_commits_info_0_debug_otherPdest_3;
        io_commits_info_0_debug_otherPdest_4 = this.vif.mon_mp.mon_cb.io_commits_info_0_debug_otherPdest_4;
        io_commits_info_0_debug_otherPdest_5 = this.vif.mon_mp.mon_cb.io_commits_info_0_debug_otherPdest_5;
        io_commits_info_0_debug_otherPdest_6 = this.vif.mon_mp.mon_cb.io_commits_info_0_debug_otherPdest_6;
        io_commits_info_0_debug_fuType = this.vif.mon_mp.mon_cb.io_commits_info_0_debug_fuType;
        io_commits_info_0_dirtyFs = this.vif.mon_mp.mon_cb.io_commits_info_0_dirtyFs;
        io_commits_info_0_dirtyVs = this.vif.mon_mp.mon_cb.io_commits_info_0_dirtyVs;
        io_commits_info_1_walk_v = this.vif.mon_mp.mon_cb.io_commits_info_1_walk_v;
        io_commits_info_1_commit_v = this.vif.mon_mp.mon_cb.io_commits_info_1_commit_v;
        io_commits_info_1_commit_w = this.vif.mon_mp.mon_cb.io_commits_info_1_commit_w;
        io_commits_info_1_realDestSize = this.vif.mon_mp.mon_cb.io_commits_info_1_realDestSize;
        io_commits_info_1_interrupt_safe = this.vif.mon_mp.mon_cb.io_commits_info_1_interrupt_safe;
        io_commits_info_1_wflags = this.vif.mon_mp.mon_cb.io_commits_info_1_wflags;
        io_commits_info_1_fflags = this.vif.mon_mp.mon_cb.io_commits_info_1_fflags;
        io_commits_info_1_vxsat = this.vif.mon_mp.mon_cb.io_commits_info_1_vxsat;
        io_commits_info_1_isRVC = this.vif.mon_mp.mon_cb.io_commits_info_1_isRVC;
        io_commits_info_1_isVset = this.vif.mon_mp.mon_cb.io_commits_info_1_isVset;
        io_commits_info_1_isHls = this.vif.mon_mp.mon_cb.io_commits_info_1_isHls;
        io_commits_info_1_isVls = this.vif.mon_mp.mon_cb.io_commits_info_1_isVls;
        io_commits_info_1_vls = this.vif.mon_mp.mon_cb.io_commits_info_1_vls;
        io_commits_info_1_mmio = this.vif.mon_mp.mon_cb.io_commits_info_1_mmio;
        io_commits_info_1_commitType = this.vif.mon_mp.mon_cb.io_commits_info_1_commitType;
        io_commits_info_1_ftqIdx_flag = this.vif.mon_mp.mon_cb.io_commits_info_1_ftqIdx_flag;
        io_commits_info_1_ftqIdx_value = this.vif.mon_mp.mon_cb.io_commits_info_1_ftqIdx_value;
        io_commits_info_1_ftqOffset = this.vif.mon_mp.mon_cb.io_commits_info_1_ftqOffset;
        io_commits_info_1_instrSize = this.vif.mon_mp.mon_cb.io_commits_info_1_instrSize;
        io_commits_info_1_fpWen = this.vif.mon_mp.mon_cb.io_commits_info_1_fpWen;
        io_commits_info_1_rfWen = this.vif.mon_mp.mon_cb.io_commits_info_1_rfWen;
        io_commits_info_1_needFlush = this.vif.mon_mp.mon_cb.io_commits_info_1_needFlush;
        io_commits_info_1_traceBlockInPipe_itype = this.vif.mon_mp.mon_cb.io_commits_info_1_traceBlockInPipe_itype;
        io_commits_info_1_traceBlockInPipe_iretire = this.vif.mon_mp.mon_cb.io_commits_info_1_traceBlockInPipe_iretire;
        io_commits_info_1_traceBlockInPipe_ilastsize = this.vif.mon_mp.mon_cb.io_commits_info_1_traceBlockInPipe_ilastsize;
        io_commits_info_1_debug_pc = this.vif.mon_mp.mon_cb.io_commits_info_1_debug_pc;
        io_commits_info_1_debug_instr = this.vif.mon_mp.mon_cb.io_commits_info_1_debug_instr;
        io_commits_info_1_debug_ldest = this.vif.mon_mp.mon_cb.io_commits_info_1_debug_ldest;
        io_commits_info_1_debug_pdest = this.vif.mon_mp.mon_cb.io_commits_info_1_debug_pdest;
        io_commits_info_1_debug_otherPdest_0 = this.vif.mon_mp.mon_cb.io_commits_info_1_debug_otherPdest_0;
        io_commits_info_1_debug_otherPdest_1 = this.vif.mon_mp.mon_cb.io_commits_info_1_debug_otherPdest_1;
        io_commits_info_1_debug_otherPdest_2 = this.vif.mon_mp.mon_cb.io_commits_info_1_debug_otherPdest_2;
        io_commits_info_1_debug_otherPdest_3 = this.vif.mon_mp.mon_cb.io_commits_info_1_debug_otherPdest_3;
        io_commits_info_1_debug_otherPdest_4 = this.vif.mon_mp.mon_cb.io_commits_info_1_debug_otherPdest_4;
        io_commits_info_1_debug_otherPdest_5 = this.vif.mon_mp.mon_cb.io_commits_info_1_debug_otherPdest_5;
        io_commits_info_1_debug_otherPdest_6 = this.vif.mon_mp.mon_cb.io_commits_info_1_debug_otherPdest_6;
        io_commits_info_1_debug_fuType = this.vif.mon_mp.mon_cb.io_commits_info_1_debug_fuType;
        io_commits_info_1_dirtyFs = this.vif.mon_mp.mon_cb.io_commits_info_1_dirtyFs;
        io_commits_info_1_dirtyVs = this.vif.mon_mp.mon_cb.io_commits_info_1_dirtyVs;
        io_commits_info_2_walk_v = this.vif.mon_mp.mon_cb.io_commits_info_2_walk_v;
        io_commits_info_2_commit_v = this.vif.mon_mp.mon_cb.io_commits_info_2_commit_v;
        io_commits_info_2_commit_w = this.vif.mon_mp.mon_cb.io_commits_info_2_commit_w;
        io_commits_info_2_realDestSize = this.vif.mon_mp.mon_cb.io_commits_info_2_realDestSize;
        io_commits_info_2_interrupt_safe = this.vif.mon_mp.mon_cb.io_commits_info_2_interrupt_safe;
        io_commits_info_2_wflags = this.vif.mon_mp.mon_cb.io_commits_info_2_wflags;
        io_commits_info_2_fflags = this.vif.mon_mp.mon_cb.io_commits_info_2_fflags;
        io_commits_info_2_vxsat = this.vif.mon_mp.mon_cb.io_commits_info_2_vxsat;
        io_commits_info_2_isRVC = this.vif.mon_mp.mon_cb.io_commits_info_2_isRVC;
        io_commits_info_2_isVset = this.vif.mon_mp.mon_cb.io_commits_info_2_isVset;
        io_commits_info_2_isHls = this.vif.mon_mp.mon_cb.io_commits_info_2_isHls;
        io_commits_info_2_isVls = this.vif.mon_mp.mon_cb.io_commits_info_2_isVls;
        io_commits_info_2_vls = this.vif.mon_mp.mon_cb.io_commits_info_2_vls;
        io_commits_info_2_mmio = this.vif.mon_mp.mon_cb.io_commits_info_2_mmio;
        io_commits_info_2_commitType = this.vif.mon_mp.mon_cb.io_commits_info_2_commitType;
        io_commits_info_2_ftqIdx_flag = this.vif.mon_mp.mon_cb.io_commits_info_2_ftqIdx_flag;
        io_commits_info_2_ftqIdx_value = this.vif.mon_mp.mon_cb.io_commits_info_2_ftqIdx_value;
        io_commits_info_2_ftqOffset = this.vif.mon_mp.mon_cb.io_commits_info_2_ftqOffset;
        io_commits_info_2_instrSize = this.vif.mon_mp.mon_cb.io_commits_info_2_instrSize;
        io_commits_info_2_fpWen = this.vif.mon_mp.mon_cb.io_commits_info_2_fpWen;
        io_commits_info_2_rfWen = this.vif.mon_mp.mon_cb.io_commits_info_2_rfWen;
        io_commits_info_2_needFlush = this.vif.mon_mp.mon_cb.io_commits_info_2_needFlush;
        io_commits_info_2_traceBlockInPipe_itype = this.vif.mon_mp.mon_cb.io_commits_info_2_traceBlockInPipe_itype;
        io_commits_info_2_traceBlockInPipe_iretire = this.vif.mon_mp.mon_cb.io_commits_info_2_traceBlockInPipe_iretire;
        io_commits_info_2_traceBlockInPipe_ilastsize = this.vif.mon_mp.mon_cb.io_commits_info_2_traceBlockInPipe_ilastsize;
        io_commits_info_2_debug_pc = this.vif.mon_mp.mon_cb.io_commits_info_2_debug_pc;
        io_commits_info_2_debug_instr = this.vif.mon_mp.mon_cb.io_commits_info_2_debug_instr;
        io_commits_info_2_debug_ldest = this.vif.mon_mp.mon_cb.io_commits_info_2_debug_ldest;
        io_commits_info_2_debug_pdest = this.vif.mon_mp.mon_cb.io_commits_info_2_debug_pdest;
        io_commits_info_2_debug_otherPdest_0 = this.vif.mon_mp.mon_cb.io_commits_info_2_debug_otherPdest_0;
        io_commits_info_2_debug_otherPdest_1 = this.vif.mon_mp.mon_cb.io_commits_info_2_debug_otherPdest_1;
        io_commits_info_2_debug_otherPdest_2 = this.vif.mon_mp.mon_cb.io_commits_info_2_debug_otherPdest_2;
        io_commits_info_2_debug_otherPdest_3 = this.vif.mon_mp.mon_cb.io_commits_info_2_debug_otherPdest_3;
        io_commits_info_2_debug_otherPdest_4 = this.vif.mon_mp.mon_cb.io_commits_info_2_debug_otherPdest_4;
        io_commits_info_2_debug_otherPdest_5 = this.vif.mon_mp.mon_cb.io_commits_info_2_debug_otherPdest_5;
        io_commits_info_2_debug_otherPdest_6 = this.vif.mon_mp.mon_cb.io_commits_info_2_debug_otherPdest_6;
        io_commits_info_2_debug_fuType = this.vif.mon_mp.mon_cb.io_commits_info_2_debug_fuType;
        io_commits_info_2_dirtyFs = this.vif.mon_mp.mon_cb.io_commits_info_2_dirtyFs;
        io_commits_info_2_dirtyVs = this.vif.mon_mp.mon_cb.io_commits_info_2_dirtyVs;
        io_commits_info_3_walk_v = this.vif.mon_mp.mon_cb.io_commits_info_3_walk_v;
        io_commits_info_3_commit_v = this.vif.mon_mp.mon_cb.io_commits_info_3_commit_v;
        io_commits_info_3_commit_w = this.vif.mon_mp.mon_cb.io_commits_info_3_commit_w;
        io_commits_info_3_realDestSize = this.vif.mon_mp.mon_cb.io_commits_info_3_realDestSize;
        io_commits_info_3_interrupt_safe = this.vif.mon_mp.mon_cb.io_commits_info_3_interrupt_safe;
        io_commits_info_3_wflags = this.vif.mon_mp.mon_cb.io_commits_info_3_wflags;
        io_commits_info_3_fflags = this.vif.mon_mp.mon_cb.io_commits_info_3_fflags;
        io_commits_info_3_vxsat = this.vif.mon_mp.mon_cb.io_commits_info_3_vxsat;
        io_commits_info_3_isRVC = this.vif.mon_mp.mon_cb.io_commits_info_3_isRVC;
        io_commits_info_3_isVset = this.vif.mon_mp.mon_cb.io_commits_info_3_isVset;
        io_commits_info_3_isHls = this.vif.mon_mp.mon_cb.io_commits_info_3_isHls;
        io_commits_info_3_isVls = this.vif.mon_mp.mon_cb.io_commits_info_3_isVls;
        io_commits_info_3_vls = this.vif.mon_mp.mon_cb.io_commits_info_3_vls;
        io_commits_info_3_mmio = this.vif.mon_mp.mon_cb.io_commits_info_3_mmio;
        io_commits_info_3_commitType = this.vif.mon_mp.mon_cb.io_commits_info_3_commitType;
        io_commits_info_3_ftqIdx_flag = this.vif.mon_mp.mon_cb.io_commits_info_3_ftqIdx_flag;
        io_commits_info_3_ftqIdx_value = this.vif.mon_mp.mon_cb.io_commits_info_3_ftqIdx_value;
        io_commits_info_3_ftqOffset = this.vif.mon_mp.mon_cb.io_commits_info_3_ftqOffset;
        io_commits_info_3_instrSize = this.vif.mon_mp.mon_cb.io_commits_info_3_instrSize;
        io_commits_info_3_fpWen = this.vif.mon_mp.mon_cb.io_commits_info_3_fpWen;
        io_commits_info_3_rfWen = this.vif.mon_mp.mon_cb.io_commits_info_3_rfWen;
        io_commits_info_3_needFlush = this.vif.mon_mp.mon_cb.io_commits_info_3_needFlush;
        io_commits_info_3_traceBlockInPipe_itype = this.vif.mon_mp.mon_cb.io_commits_info_3_traceBlockInPipe_itype;
        io_commits_info_3_traceBlockInPipe_iretire = this.vif.mon_mp.mon_cb.io_commits_info_3_traceBlockInPipe_iretire;
        io_commits_info_3_traceBlockInPipe_ilastsize = this.vif.mon_mp.mon_cb.io_commits_info_3_traceBlockInPipe_ilastsize;
        io_commits_info_3_debug_pc = this.vif.mon_mp.mon_cb.io_commits_info_3_debug_pc;
        io_commits_info_3_debug_instr = this.vif.mon_mp.mon_cb.io_commits_info_3_debug_instr;
        io_commits_info_3_debug_ldest = this.vif.mon_mp.mon_cb.io_commits_info_3_debug_ldest;
        io_commits_info_3_debug_pdest = this.vif.mon_mp.mon_cb.io_commits_info_3_debug_pdest;
        io_commits_info_3_debug_otherPdest_0 = this.vif.mon_mp.mon_cb.io_commits_info_3_debug_otherPdest_0;
        io_commits_info_3_debug_otherPdest_1 = this.vif.mon_mp.mon_cb.io_commits_info_3_debug_otherPdest_1;
        io_commits_info_3_debug_otherPdest_2 = this.vif.mon_mp.mon_cb.io_commits_info_3_debug_otherPdest_2;
        io_commits_info_3_debug_otherPdest_3 = this.vif.mon_mp.mon_cb.io_commits_info_3_debug_otherPdest_3;
        io_commits_info_3_debug_otherPdest_4 = this.vif.mon_mp.mon_cb.io_commits_info_3_debug_otherPdest_4;
        io_commits_info_3_debug_otherPdest_5 = this.vif.mon_mp.mon_cb.io_commits_info_3_debug_otherPdest_5;
        io_commits_info_3_debug_otherPdest_6 = this.vif.mon_mp.mon_cb.io_commits_info_3_debug_otherPdest_6;
        io_commits_info_3_debug_fuType = this.vif.mon_mp.mon_cb.io_commits_info_3_debug_fuType;
        io_commits_info_3_dirtyFs = this.vif.mon_mp.mon_cb.io_commits_info_3_dirtyFs;
        io_commits_info_3_dirtyVs = this.vif.mon_mp.mon_cb.io_commits_info_3_dirtyVs;
        io_commits_info_4_walk_v = this.vif.mon_mp.mon_cb.io_commits_info_4_walk_v;
        io_commits_info_4_commit_v = this.vif.mon_mp.mon_cb.io_commits_info_4_commit_v;
        io_commits_info_4_commit_w = this.vif.mon_mp.mon_cb.io_commits_info_4_commit_w;
        io_commits_info_4_realDestSize = this.vif.mon_mp.mon_cb.io_commits_info_4_realDestSize;
        io_commits_info_4_interrupt_safe = this.vif.mon_mp.mon_cb.io_commits_info_4_interrupt_safe;
        io_commits_info_4_wflags = this.vif.mon_mp.mon_cb.io_commits_info_4_wflags;
        io_commits_info_4_fflags = this.vif.mon_mp.mon_cb.io_commits_info_4_fflags;
        io_commits_info_4_vxsat = this.vif.mon_mp.mon_cb.io_commits_info_4_vxsat;
        io_commits_info_4_isRVC = this.vif.mon_mp.mon_cb.io_commits_info_4_isRVC;
        io_commits_info_4_isVset = this.vif.mon_mp.mon_cb.io_commits_info_4_isVset;
        io_commits_info_4_isHls = this.vif.mon_mp.mon_cb.io_commits_info_4_isHls;
        io_commits_info_4_isVls = this.vif.mon_mp.mon_cb.io_commits_info_4_isVls;
        io_commits_info_4_vls = this.vif.mon_mp.mon_cb.io_commits_info_4_vls;
        io_commits_info_4_mmio = this.vif.mon_mp.mon_cb.io_commits_info_4_mmio;
        io_commits_info_4_commitType = this.vif.mon_mp.mon_cb.io_commits_info_4_commitType;
        io_commits_info_4_ftqIdx_flag = this.vif.mon_mp.mon_cb.io_commits_info_4_ftqIdx_flag;
        io_commits_info_4_ftqIdx_value = this.vif.mon_mp.mon_cb.io_commits_info_4_ftqIdx_value;
        io_commits_info_4_ftqOffset = this.vif.mon_mp.mon_cb.io_commits_info_4_ftqOffset;
        io_commits_info_4_instrSize = this.vif.mon_mp.mon_cb.io_commits_info_4_instrSize;
        io_commits_info_4_fpWen = this.vif.mon_mp.mon_cb.io_commits_info_4_fpWen;
        io_commits_info_4_rfWen = this.vif.mon_mp.mon_cb.io_commits_info_4_rfWen;
        io_commits_info_4_needFlush = this.vif.mon_mp.mon_cb.io_commits_info_4_needFlush;
        io_commits_info_4_traceBlockInPipe_itype = this.vif.mon_mp.mon_cb.io_commits_info_4_traceBlockInPipe_itype;
        io_commits_info_4_traceBlockInPipe_iretire = this.vif.mon_mp.mon_cb.io_commits_info_4_traceBlockInPipe_iretire;
        io_commits_info_4_traceBlockInPipe_ilastsize = this.vif.mon_mp.mon_cb.io_commits_info_4_traceBlockInPipe_ilastsize;
        io_commits_info_4_debug_pc = this.vif.mon_mp.mon_cb.io_commits_info_4_debug_pc;
        io_commits_info_4_debug_instr = this.vif.mon_mp.mon_cb.io_commits_info_4_debug_instr;
        io_commits_info_4_debug_ldest = this.vif.mon_mp.mon_cb.io_commits_info_4_debug_ldest;
        io_commits_info_4_debug_pdest = this.vif.mon_mp.mon_cb.io_commits_info_4_debug_pdest;
        io_commits_info_4_debug_otherPdest_0 = this.vif.mon_mp.mon_cb.io_commits_info_4_debug_otherPdest_0;
        io_commits_info_4_debug_otherPdest_1 = this.vif.mon_mp.mon_cb.io_commits_info_4_debug_otherPdest_1;
        io_commits_info_4_debug_otherPdest_2 = this.vif.mon_mp.mon_cb.io_commits_info_4_debug_otherPdest_2;
        io_commits_info_4_debug_otherPdest_3 = this.vif.mon_mp.mon_cb.io_commits_info_4_debug_otherPdest_3;
        io_commits_info_4_debug_otherPdest_4 = this.vif.mon_mp.mon_cb.io_commits_info_4_debug_otherPdest_4;
        io_commits_info_4_debug_otherPdest_5 = this.vif.mon_mp.mon_cb.io_commits_info_4_debug_otherPdest_5;
        io_commits_info_4_debug_otherPdest_6 = this.vif.mon_mp.mon_cb.io_commits_info_4_debug_otherPdest_6;
        io_commits_info_4_debug_fuType = this.vif.mon_mp.mon_cb.io_commits_info_4_debug_fuType;
        io_commits_info_4_dirtyFs = this.vif.mon_mp.mon_cb.io_commits_info_4_dirtyFs;
        io_commits_info_4_dirtyVs = this.vif.mon_mp.mon_cb.io_commits_info_4_dirtyVs;
        io_commits_info_5_walk_v = this.vif.mon_mp.mon_cb.io_commits_info_5_walk_v;
        io_commits_info_5_commit_v = this.vif.mon_mp.mon_cb.io_commits_info_5_commit_v;
        io_commits_info_5_commit_w = this.vif.mon_mp.mon_cb.io_commits_info_5_commit_w;
        io_commits_info_5_realDestSize = this.vif.mon_mp.mon_cb.io_commits_info_5_realDestSize;
        io_commits_info_5_interrupt_safe = this.vif.mon_mp.mon_cb.io_commits_info_5_interrupt_safe;
        io_commits_info_5_wflags = this.vif.mon_mp.mon_cb.io_commits_info_5_wflags;
        io_commits_info_5_fflags = this.vif.mon_mp.mon_cb.io_commits_info_5_fflags;
        io_commits_info_5_vxsat = this.vif.mon_mp.mon_cb.io_commits_info_5_vxsat;
        io_commits_info_5_isRVC = this.vif.mon_mp.mon_cb.io_commits_info_5_isRVC;
        io_commits_info_5_isVset = this.vif.mon_mp.mon_cb.io_commits_info_5_isVset;
        io_commits_info_5_isHls = this.vif.mon_mp.mon_cb.io_commits_info_5_isHls;
        io_commits_info_5_isVls = this.vif.mon_mp.mon_cb.io_commits_info_5_isVls;
        io_commits_info_5_vls = this.vif.mon_mp.mon_cb.io_commits_info_5_vls;
        io_commits_info_5_mmio = this.vif.mon_mp.mon_cb.io_commits_info_5_mmio;
        io_commits_info_5_commitType = this.vif.mon_mp.mon_cb.io_commits_info_5_commitType;
        io_commits_info_5_ftqIdx_flag = this.vif.mon_mp.mon_cb.io_commits_info_5_ftqIdx_flag;
        io_commits_info_5_ftqIdx_value = this.vif.mon_mp.mon_cb.io_commits_info_5_ftqIdx_value;
        io_commits_info_5_ftqOffset = this.vif.mon_mp.mon_cb.io_commits_info_5_ftqOffset;
        io_commits_info_5_instrSize = this.vif.mon_mp.mon_cb.io_commits_info_5_instrSize;
        io_commits_info_5_fpWen = this.vif.mon_mp.mon_cb.io_commits_info_5_fpWen;
        io_commits_info_5_rfWen = this.vif.mon_mp.mon_cb.io_commits_info_5_rfWen;
        io_commits_info_5_needFlush = this.vif.mon_mp.mon_cb.io_commits_info_5_needFlush;
        io_commits_info_5_traceBlockInPipe_itype = this.vif.mon_mp.mon_cb.io_commits_info_5_traceBlockInPipe_itype;
        io_commits_info_5_traceBlockInPipe_iretire = this.vif.mon_mp.mon_cb.io_commits_info_5_traceBlockInPipe_iretire;
        io_commits_info_5_traceBlockInPipe_ilastsize = this.vif.mon_mp.mon_cb.io_commits_info_5_traceBlockInPipe_ilastsize;
        io_commits_info_5_debug_pc = this.vif.mon_mp.mon_cb.io_commits_info_5_debug_pc;
        io_commits_info_5_debug_instr = this.vif.mon_mp.mon_cb.io_commits_info_5_debug_instr;
        io_commits_info_5_debug_ldest = this.vif.mon_mp.mon_cb.io_commits_info_5_debug_ldest;
        io_commits_info_5_debug_pdest = this.vif.mon_mp.mon_cb.io_commits_info_5_debug_pdest;
        io_commits_info_5_debug_otherPdest_0 = this.vif.mon_mp.mon_cb.io_commits_info_5_debug_otherPdest_0;
        io_commits_info_5_debug_otherPdest_1 = this.vif.mon_mp.mon_cb.io_commits_info_5_debug_otherPdest_1;
        io_commits_info_5_debug_otherPdest_2 = this.vif.mon_mp.mon_cb.io_commits_info_5_debug_otherPdest_2;
        io_commits_info_5_debug_otherPdest_3 = this.vif.mon_mp.mon_cb.io_commits_info_5_debug_otherPdest_3;
        io_commits_info_5_debug_otherPdest_4 = this.vif.mon_mp.mon_cb.io_commits_info_5_debug_otherPdest_4;
        io_commits_info_5_debug_otherPdest_5 = this.vif.mon_mp.mon_cb.io_commits_info_5_debug_otherPdest_5;
        io_commits_info_5_debug_otherPdest_6 = this.vif.mon_mp.mon_cb.io_commits_info_5_debug_otherPdest_6;
        io_commits_info_5_debug_fuType = this.vif.mon_mp.mon_cb.io_commits_info_5_debug_fuType;
        io_commits_info_5_dirtyFs = this.vif.mon_mp.mon_cb.io_commits_info_5_dirtyFs;
        io_commits_info_5_dirtyVs = this.vif.mon_mp.mon_cb.io_commits_info_5_dirtyVs;
        io_commits_info_6_walk_v = this.vif.mon_mp.mon_cb.io_commits_info_6_walk_v;
        io_commits_info_6_commit_v = this.vif.mon_mp.mon_cb.io_commits_info_6_commit_v;
        io_commits_info_6_commit_w = this.vif.mon_mp.mon_cb.io_commits_info_6_commit_w;
        io_commits_info_6_realDestSize = this.vif.mon_mp.mon_cb.io_commits_info_6_realDestSize;
        io_commits_info_6_interrupt_safe = this.vif.mon_mp.mon_cb.io_commits_info_6_interrupt_safe;
        io_commits_info_6_wflags = this.vif.mon_mp.mon_cb.io_commits_info_6_wflags;
        io_commits_info_6_fflags = this.vif.mon_mp.mon_cb.io_commits_info_6_fflags;
        io_commits_info_6_vxsat = this.vif.mon_mp.mon_cb.io_commits_info_6_vxsat;
        io_commits_info_6_isRVC = this.vif.mon_mp.mon_cb.io_commits_info_6_isRVC;
        io_commits_info_6_isVset = this.vif.mon_mp.mon_cb.io_commits_info_6_isVset;
        io_commits_info_6_isHls = this.vif.mon_mp.mon_cb.io_commits_info_6_isHls;
        io_commits_info_6_isVls = this.vif.mon_mp.mon_cb.io_commits_info_6_isVls;
        io_commits_info_6_vls = this.vif.mon_mp.mon_cb.io_commits_info_6_vls;
        io_commits_info_6_mmio = this.vif.mon_mp.mon_cb.io_commits_info_6_mmio;
        io_commits_info_6_commitType = this.vif.mon_mp.mon_cb.io_commits_info_6_commitType;
        io_commits_info_6_ftqIdx_flag = this.vif.mon_mp.mon_cb.io_commits_info_6_ftqIdx_flag;
        io_commits_info_6_ftqIdx_value = this.vif.mon_mp.mon_cb.io_commits_info_6_ftqIdx_value;
        io_commits_info_6_ftqOffset = this.vif.mon_mp.mon_cb.io_commits_info_6_ftqOffset;
        io_commits_info_6_instrSize = this.vif.mon_mp.mon_cb.io_commits_info_6_instrSize;
        io_commits_info_6_fpWen = this.vif.mon_mp.mon_cb.io_commits_info_6_fpWen;
        io_commits_info_6_rfWen = this.vif.mon_mp.mon_cb.io_commits_info_6_rfWen;
        io_commits_info_6_needFlush = this.vif.mon_mp.mon_cb.io_commits_info_6_needFlush;
        io_commits_info_6_traceBlockInPipe_itype = this.vif.mon_mp.mon_cb.io_commits_info_6_traceBlockInPipe_itype;
        io_commits_info_6_traceBlockInPipe_iretire = this.vif.mon_mp.mon_cb.io_commits_info_6_traceBlockInPipe_iretire;
        io_commits_info_6_traceBlockInPipe_ilastsize = this.vif.mon_mp.mon_cb.io_commits_info_6_traceBlockInPipe_ilastsize;
        io_commits_info_6_debug_pc = this.vif.mon_mp.mon_cb.io_commits_info_6_debug_pc;
        io_commits_info_6_debug_instr = this.vif.mon_mp.mon_cb.io_commits_info_6_debug_instr;
        io_commits_info_6_debug_ldest = this.vif.mon_mp.mon_cb.io_commits_info_6_debug_ldest;
        io_commits_info_6_debug_pdest = this.vif.mon_mp.mon_cb.io_commits_info_6_debug_pdest;
        io_commits_info_6_debug_otherPdest_0 = this.vif.mon_mp.mon_cb.io_commits_info_6_debug_otherPdest_0;
        io_commits_info_6_debug_otherPdest_1 = this.vif.mon_mp.mon_cb.io_commits_info_6_debug_otherPdest_1;
        io_commits_info_6_debug_otherPdest_2 = this.vif.mon_mp.mon_cb.io_commits_info_6_debug_otherPdest_2;
        io_commits_info_6_debug_otherPdest_3 = this.vif.mon_mp.mon_cb.io_commits_info_6_debug_otherPdest_3;
        io_commits_info_6_debug_otherPdest_4 = this.vif.mon_mp.mon_cb.io_commits_info_6_debug_otherPdest_4;
        io_commits_info_6_debug_otherPdest_5 = this.vif.mon_mp.mon_cb.io_commits_info_6_debug_otherPdest_5;
        io_commits_info_6_debug_otherPdest_6 = this.vif.mon_mp.mon_cb.io_commits_info_6_debug_otherPdest_6;
        io_commits_info_6_debug_fuType = this.vif.mon_mp.mon_cb.io_commits_info_6_debug_fuType;
        io_commits_info_6_dirtyFs = this.vif.mon_mp.mon_cb.io_commits_info_6_dirtyFs;
        io_commits_info_6_dirtyVs = this.vif.mon_mp.mon_cb.io_commits_info_6_dirtyVs;
        io_commits_info_7_walk_v = this.vif.mon_mp.mon_cb.io_commits_info_7_walk_v;
        io_commits_info_7_commit_v = this.vif.mon_mp.mon_cb.io_commits_info_7_commit_v;
        io_commits_info_7_commit_w = this.vif.mon_mp.mon_cb.io_commits_info_7_commit_w;
        io_commits_info_7_realDestSize = this.vif.mon_mp.mon_cb.io_commits_info_7_realDestSize;
        io_commits_info_7_interrupt_safe = this.vif.mon_mp.mon_cb.io_commits_info_7_interrupt_safe;
        io_commits_info_7_wflags = this.vif.mon_mp.mon_cb.io_commits_info_7_wflags;
        io_commits_info_7_fflags = this.vif.mon_mp.mon_cb.io_commits_info_7_fflags;
        io_commits_info_7_vxsat = this.vif.mon_mp.mon_cb.io_commits_info_7_vxsat;
        io_commits_info_7_isRVC = this.vif.mon_mp.mon_cb.io_commits_info_7_isRVC;
        io_commits_info_7_isVset = this.vif.mon_mp.mon_cb.io_commits_info_7_isVset;
        io_commits_info_7_isHls = this.vif.mon_mp.mon_cb.io_commits_info_7_isHls;
        io_commits_info_7_isVls = this.vif.mon_mp.mon_cb.io_commits_info_7_isVls;
        io_commits_info_7_vls = this.vif.mon_mp.mon_cb.io_commits_info_7_vls;
        io_commits_info_7_mmio = this.vif.mon_mp.mon_cb.io_commits_info_7_mmio;
        io_commits_info_7_commitType = this.vif.mon_mp.mon_cb.io_commits_info_7_commitType;
        io_commits_info_7_ftqIdx_flag = this.vif.mon_mp.mon_cb.io_commits_info_7_ftqIdx_flag;
        io_commits_info_7_ftqIdx_value = this.vif.mon_mp.mon_cb.io_commits_info_7_ftqIdx_value;
        io_commits_info_7_ftqOffset = this.vif.mon_mp.mon_cb.io_commits_info_7_ftqOffset;
        io_commits_info_7_instrSize = this.vif.mon_mp.mon_cb.io_commits_info_7_instrSize;
        io_commits_info_7_fpWen = this.vif.mon_mp.mon_cb.io_commits_info_7_fpWen;
        io_commits_info_7_rfWen = this.vif.mon_mp.mon_cb.io_commits_info_7_rfWen;
        io_commits_info_7_needFlush = this.vif.mon_mp.mon_cb.io_commits_info_7_needFlush;
        io_commits_info_7_traceBlockInPipe_itype = this.vif.mon_mp.mon_cb.io_commits_info_7_traceBlockInPipe_itype;
        io_commits_info_7_traceBlockInPipe_iretire = this.vif.mon_mp.mon_cb.io_commits_info_7_traceBlockInPipe_iretire;
        io_commits_info_7_traceBlockInPipe_ilastsize = this.vif.mon_mp.mon_cb.io_commits_info_7_traceBlockInPipe_ilastsize;
        io_commits_info_7_debug_pc = this.vif.mon_mp.mon_cb.io_commits_info_7_debug_pc;
        io_commits_info_7_debug_instr = this.vif.mon_mp.mon_cb.io_commits_info_7_debug_instr;
        io_commits_info_7_debug_ldest = this.vif.mon_mp.mon_cb.io_commits_info_7_debug_ldest;
        io_commits_info_7_debug_pdest = this.vif.mon_mp.mon_cb.io_commits_info_7_debug_pdest;
        io_commits_info_7_debug_otherPdest_0 = this.vif.mon_mp.mon_cb.io_commits_info_7_debug_otherPdest_0;
        io_commits_info_7_debug_otherPdest_1 = this.vif.mon_mp.mon_cb.io_commits_info_7_debug_otherPdest_1;
        io_commits_info_7_debug_otherPdest_2 = this.vif.mon_mp.mon_cb.io_commits_info_7_debug_otherPdest_2;
        io_commits_info_7_debug_otherPdest_3 = this.vif.mon_mp.mon_cb.io_commits_info_7_debug_otherPdest_3;
        io_commits_info_7_debug_otherPdest_4 = this.vif.mon_mp.mon_cb.io_commits_info_7_debug_otherPdest_4;
        io_commits_info_7_debug_otherPdest_5 = this.vif.mon_mp.mon_cb.io_commits_info_7_debug_otherPdest_5;
        io_commits_info_7_debug_otherPdest_6 = this.vif.mon_mp.mon_cb.io_commits_info_7_debug_otherPdest_6;
        io_commits_info_7_debug_fuType = this.vif.mon_mp.mon_cb.io_commits_info_7_debug_fuType;
        io_commits_info_7_dirtyFs = this.vif.mon_mp.mon_cb.io_commits_info_7_dirtyFs;
        io_commits_info_7_dirtyVs = this.vif.mon_mp.mon_cb.io_commits_info_7_dirtyVs;
        io_commits_robIdx_0_flag = this.vif.mon_mp.mon_cb.io_commits_robIdx_0_flag;
        io_commits_robIdx_0_value = this.vif.mon_mp.mon_cb.io_commits_robIdx_0_value;
        io_commits_robIdx_1_flag = this.vif.mon_mp.mon_cb.io_commits_robIdx_1_flag;
        io_commits_robIdx_1_value = this.vif.mon_mp.mon_cb.io_commits_robIdx_1_value;
        io_commits_robIdx_2_flag = this.vif.mon_mp.mon_cb.io_commits_robIdx_2_flag;
        io_commits_robIdx_2_value = this.vif.mon_mp.mon_cb.io_commits_robIdx_2_value;
        io_commits_robIdx_3_flag = this.vif.mon_mp.mon_cb.io_commits_robIdx_3_flag;
        io_commits_robIdx_3_value = this.vif.mon_mp.mon_cb.io_commits_robIdx_3_value;
        io_commits_robIdx_4_flag = this.vif.mon_mp.mon_cb.io_commits_robIdx_4_flag;
        io_commits_robIdx_4_value = this.vif.mon_mp.mon_cb.io_commits_robIdx_4_value;
        io_commits_robIdx_5_flag = this.vif.mon_mp.mon_cb.io_commits_robIdx_5_flag;
        io_commits_robIdx_5_value = this.vif.mon_mp.mon_cb.io_commits_robIdx_5_value;
        io_commits_robIdx_6_flag = this.vif.mon_mp.mon_cb.io_commits_robIdx_6_flag;
        io_commits_robIdx_6_value = this.vif.mon_mp.mon_cb.io_commits_robIdx_6_value;
        io_commits_robIdx_7_flag = this.vif.mon_mp.mon_cb.io_commits_robIdx_7_flag;
        io_commits_robIdx_7_value = this.vif.mon_mp.mon_cb.io_commits_robIdx_7_value;
        io_trace_blockCommit = this.vif.mon_mp.mon_cb.io_trace_blockCommit;
        io_trace_traceCommitInfo_blocks_0_valid = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_0_valid;
        io_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value;
        io_trace_traceCommitInfo_blocks_0_bits_ftqOffset = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_0_bits_ftqOffset;
        io_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype;
        io_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire;
        io_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize;
        io_trace_traceCommitInfo_blocks_1_valid = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_1_valid;
        io_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value;
        io_trace_traceCommitInfo_blocks_1_bits_ftqOffset = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_1_bits_ftqOffset;
        io_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype;
        io_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire;
        io_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize;
        io_trace_traceCommitInfo_blocks_2_valid = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_2_valid;
        io_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value;
        io_trace_traceCommitInfo_blocks_2_bits_ftqOffset = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_2_bits_ftqOffset;
        io_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype;
        io_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire;
        io_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize;
        io_trace_traceCommitInfo_blocks_3_valid = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_3_valid;
        io_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value;
        io_trace_traceCommitInfo_blocks_3_bits_ftqOffset = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_3_bits_ftqOffset;
        io_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype;
        io_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire;
        io_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize;
        io_trace_traceCommitInfo_blocks_4_valid = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_4_valid;
        io_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value;
        io_trace_traceCommitInfo_blocks_4_bits_ftqOffset = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_4_bits_ftqOffset;
        io_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype;
        io_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire;
        io_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize;
        io_trace_traceCommitInfo_blocks_5_valid = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_5_valid;
        io_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value;
        io_trace_traceCommitInfo_blocks_5_bits_ftqOffset = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_5_bits_ftqOffset;
        io_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype;
        io_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire;
        io_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize;
        io_trace_traceCommitInfo_blocks_6_valid = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_6_valid;
        io_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value;
        io_trace_traceCommitInfo_blocks_6_bits_ftqOffset = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_6_bits_ftqOffset;
        io_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype;
        io_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire;
        io_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize;
        io_trace_traceCommitInfo_blocks_7_valid = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_7_valid;
        io_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value;
        io_trace_traceCommitInfo_blocks_7_bits_ftqOffset = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_7_bits_ftqOffset;
        io_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype;
        io_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire;
        io_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize = this.vif.mon_mp.mon_cb.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize;
        io_rabCommits_isCommit = this.vif.mon_mp.mon_cb.io_rabCommits_isCommit;
        io_rabCommits_commitValid_0 = this.vif.mon_mp.mon_cb.io_rabCommits_commitValid_0;
        io_rabCommits_commitValid_1 = this.vif.mon_mp.mon_cb.io_rabCommits_commitValid_1;
        io_rabCommits_commitValid_2 = this.vif.mon_mp.mon_cb.io_rabCommits_commitValid_2;
        io_rabCommits_commitValid_3 = this.vif.mon_mp.mon_cb.io_rabCommits_commitValid_3;
        io_rabCommits_commitValid_4 = this.vif.mon_mp.mon_cb.io_rabCommits_commitValid_4;
        io_rabCommits_commitValid_5 = this.vif.mon_mp.mon_cb.io_rabCommits_commitValid_5;
        io_rabCommits_isWalk = this.vif.mon_mp.mon_cb.io_rabCommits_isWalk;
        io_rabCommits_walkValid_0 = this.vif.mon_mp.mon_cb.io_rabCommits_walkValid_0;
        io_rabCommits_walkValid_1 = this.vif.mon_mp.mon_cb.io_rabCommits_walkValid_1;
        io_rabCommits_walkValid_2 = this.vif.mon_mp.mon_cb.io_rabCommits_walkValid_2;
        io_rabCommits_walkValid_3 = this.vif.mon_mp.mon_cb.io_rabCommits_walkValid_3;
        io_rabCommits_walkValid_4 = this.vif.mon_mp.mon_cb.io_rabCommits_walkValid_4;
        io_rabCommits_walkValid_5 = this.vif.mon_mp.mon_cb.io_rabCommits_walkValid_5;
        io_rabCommits_info_0_ldest = this.vif.mon_mp.mon_cb.io_rabCommits_info_0_ldest;
        io_rabCommits_info_0_pdest = this.vif.mon_mp.mon_cb.io_rabCommits_info_0_pdest;
        io_rabCommits_info_0_rfWen = this.vif.mon_mp.mon_cb.io_rabCommits_info_0_rfWen;
        io_rabCommits_info_0_fpWen = this.vif.mon_mp.mon_cb.io_rabCommits_info_0_fpWen;
        io_rabCommits_info_0_vecWen = this.vif.mon_mp.mon_cb.io_rabCommits_info_0_vecWen;
        io_rabCommits_info_0_v0Wen = this.vif.mon_mp.mon_cb.io_rabCommits_info_0_v0Wen;
        io_rabCommits_info_0_vlWen = this.vif.mon_mp.mon_cb.io_rabCommits_info_0_vlWen;
        io_rabCommits_info_0_isMove = this.vif.mon_mp.mon_cb.io_rabCommits_info_0_isMove;
        io_rabCommits_info_1_ldest = this.vif.mon_mp.mon_cb.io_rabCommits_info_1_ldest;
        io_rabCommits_info_1_pdest = this.vif.mon_mp.mon_cb.io_rabCommits_info_1_pdest;
        io_rabCommits_info_1_rfWen = this.vif.mon_mp.mon_cb.io_rabCommits_info_1_rfWen;
        io_rabCommits_info_1_fpWen = this.vif.mon_mp.mon_cb.io_rabCommits_info_1_fpWen;
        io_rabCommits_info_1_vecWen = this.vif.mon_mp.mon_cb.io_rabCommits_info_1_vecWen;
        io_rabCommits_info_1_v0Wen = this.vif.mon_mp.mon_cb.io_rabCommits_info_1_v0Wen;
        io_rabCommits_info_1_vlWen = this.vif.mon_mp.mon_cb.io_rabCommits_info_1_vlWen;
        io_rabCommits_info_1_isMove = this.vif.mon_mp.mon_cb.io_rabCommits_info_1_isMove;
        io_rabCommits_info_2_ldest = this.vif.mon_mp.mon_cb.io_rabCommits_info_2_ldest;
        io_rabCommits_info_2_pdest = this.vif.mon_mp.mon_cb.io_rabCommits_info_2_pdest;
        io_rabCommits_info_2_rfWen = this.vif.mon_mp.mon_cb.io_rabCommits_info_2_rfWen;
        io_rabCommits_info_2_fpWen = this.vif.mon_mp.mon_cb.io_rabCommits_info_2_fpWen;
        io_rabCommits_info_2_vecWen = this.vif.mon_mp.mon_cb.io_rabCommits_info_2_vecWen;
        io_rabCommits_info_2_v0Wen = this.vif.mon_mp.mon_cb.io_rabCommits_info_2_v0Wen;
        io_rabCommits_info_2_vlWen = this.vif.mon_mp.mon_cb.io_rabCommits_info_2_vlWen;
        io_rabCommits_info_2_isMove = this.vif.mon_mp.mon_cb.io_rabCommits_info_2_isMove;
        io_rabCommits_info_3_ldest = this.vif.mon_mp.mon_cb.io_rabCommits_info_3_ldest;
        io_rabCommits_info_3_pdest = this.vif.mon_mp.mon_cb.io_rabCommits_info_3_pdest;
        io_rabCommits_info_3_rfWen = this.vif.mon_mp.mon_cb.io_rabCommits_info_3_rfWen;
        io_rabCommits_info_3_fpWen = this.vif.mon_mp.mon_cb.io_rabCommits_info_3_fpWen;
        io_rabCommits_info_3_vecWen = this.vif.mon_mp.mon_cb.io_rabCommits_info_3_vecWen;
        io_rabCommits_info_3_v0Wen = this.vif.mon_mp.mon_cb.io_rabCommits_info_3_v0Wen;
        io_rabCommits_info_3_vlWen = this.vif.mon_mp.mon_cb.io_rabCommits_info_3_vlWen;
        io_rabCommits_info_3_isMove = this.vif.mon_mp.mon_cb.io_rabCommits_info_3_isMove;
        io_rabCommits_info_4_ldest = this.vif.mon_mp.mon_cb.io_rabCommits_info_4_ldest;
        io_rabCommits_info_4_pdest = this.vif.mon_mp.mon_cb.io_rabCommits_info_4_pdest;
        io_rabCommits_info_4_rfWen = this.vif.mon_mp.mon_cb.io_rabCommits_info_4_rfWen;
        io_rabCommits_info_4_fpWen = this.vif.mon_mp.mon_cb.io_rabCommits_info_4_fpWen;
        io_rabCommits_info_4_vecWen = this.vif.mon_mp.mon_cb.io_rabCommits_info_4_vecWen;
        io_rabCommits_info_4_v0Wen = this.vif.mon_mp.mon_cb.io_rabCommits_info_4_v0Wen;
        io_rabCommits_info_4_vlWen = this.vif.mon_mp.mon_cb.io_rabCommits_info_4_vlWen;
        io_rabCommits_info_4_isMove = this.vif.mon_mp.mon_cb.io_rabCommits_info_4_isMove;
        io_rabCommits_info_5_ldest = this.vif.mon_mp.mon_cb.io_rabCommits_info_5_ldest;
        io_rabCommits_info_5_pdest = this.vif.mon_mp.mon_cb.io_rabCommits_info_5_pdest;
        io_rabCommits_info_5_rfWen = this.vif.mon_mp.mon_cb.io_rabCommits_info_5_rfWen;
        io_rabCommits_info_5_fpWen = this.vif.mon_mp.mon_cb.io_rabCommits_info_5_fpWen;
        io_rabCommits_info_5_vecWen = this.vif.mon_mp.mon_cb.io_rabCommits_info_5_vecWen;
        io_rabCommits_info_5_v0Wen = this.vif.mon_mp.mon_cb.io_rabCommits_info_5_v0Wen;
        io_rabCommits_info_5_vlWen = this.vif.mon_mp.mon_cb.io_rabCommits_info_5_vlWen;
        io_rabCommits_info_5_isMove = this.vif.mon_mp.mon_cb.io_rabCommits_info_5_isMove;
        io_diffCommits_commitValid_0 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_0;
        io_diffCommits_commitValid_1 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_1;
        io_diffCommits_commitValid_2 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_2;
        io_diffCommits_commitValid_3 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_3;
        io_diffCommits_commitValid_4 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_4;
        io_diffCommits_commitValid_5 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_5;
        io_diffCommits_commitValid_6 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_6;
        io_diffCommits_commitValid_7 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_7;
        io_diffCommits_commitValid_8 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_8;
        io_diffCommits_commitValid_9 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_9;
        io_diffCommits_commitValid_10 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_10;
        io_diffCommits_commitValid_11 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_11;
        io_diffCommits_commitValid_12 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_12;
        io_diffCommits_commitValid_13 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_13;
        io_diffCommits_commitValid_14 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_14;
        io_diffCommits_commitValid_15 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_15;
        io_diffCommits_commitValid_16 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_16;
        io_diffCommits_commitValid_17 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_17;
        io_diffCommits_commitValid_18 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_18;
        io_diffCommits_commitValid_19 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_19;
        io_diffCommits_commitValid_20 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_20;
        io_diffCommits_commitValid_21 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_21;
        io_diffCommits_commitValid_22 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_22;
        io_diffCommits_commitValid_23 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_23;
        io_diffCommits_commitValid_24 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_24;
        io_diffCommits_commitValid_25 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_25;
        io_diffCommits_commitValid_26 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_26;
        io_diffCommits_commitValid_27 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_27;
        io_diffCommits_commitValid_28 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_28;
        io_diffCommits_commitValid_29 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_29;
        io_diffCommits_commitValid_30 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_30;
        io_diffCommits_commitValid_31 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_31;
        io_diffCommits_commitValid_32 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_32;
        io_diffCommits_commitValid_33 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_33;
        io_diffCommits_commitValid_34 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_34;
        io_diffCommits_commitValid_35 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_35;
        io_diffCommits_commitValid_36 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_36;
        io_diffCommits_commitValid_37 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_37;
        io_diffCommits_commitValid_38 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_38;
        io_diffCommits_commitValid_39 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_39;
        io_diffCommits_commitValid_40 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_40;
        io_diffCommits_commitValid_41 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_41;
        io_diffCommits_commitValid_42 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_42;
        io_diffCommits_commitValid_43 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_43;
        io_diffCommits_commitValid_44 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_44;
        io_diffCommits_commitValid_45 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_45;
        io_diffCommits_commitValid_46 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_46;
        io_diffCommits_commitValid_47 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_47;
        io_diffCommits_commitValid_48 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_48;
        io_diffCommits_commitValid_49 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_49;
        io_diffCommits_commitValid_50 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_50;
        io_diffCommits_commitValid_51 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_51;
        io_diffCommits_commitValid_52 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_52;
        io_diffCommits_commitValid_53 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_53;
        io_diffCommits_commitValid_54 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_54;
        io_diffCommits_commitValid_55 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_55;
        io_diffCommits_commitValid_56 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_56;
        io_diffCommits_commitValid_57 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_57;
        io_diffCommits_commitValid_58 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_58;
        io_diffCommits_commitValid_59 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_59;
        io_diffCommits_commitValid_60 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_60;
        io_diffCommits_commitValid_61 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_61;
        io_diffCommits_commitValid_62 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_62;
        io_diffCommits_commitValid_63 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_63;
        io_diffCommits_commitValid_64 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_64;
        io_diffCommits_commitValid_65 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_65;
        io_diffCommits_commitValid_66 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_66;
        io_diffCommits_commitValid_67 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_67;
        io_diffCommits_commitValid_68 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_68;
        io_diffCommits_commitValid_69 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_69;
        io_diffCommits_commitValid_70 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_70;
        io_diffCommits_commitValid_71 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_71;
        io_diffCommits_commitValid_72 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_72;
        io_diffCommits_commitValid_73 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_73;
        io_diffCommits_commitValid_74 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_74;
        io_diffCommits_commitValid_75 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_75;
        io_diffCommits_commitValid_76 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_76;
        io_diffCommits_commitValid_77 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_77;
        io_diffCommits_commitValid_78 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_78;
        io_diffCommits_commitValid_79 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_79;
        io_diffCommits_commitValid_80 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_80;
        io_diffCommits_commitValid_81 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_81;
        io_diffCommits_commitValid_82 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_82;
        io_diffCommits_commitValid_83 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_83;
        io_diffCommits_commitValid_84 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_84;
        io_diffCommits_commitValid_85 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_85;
        io_diffCommits_commitValid_86 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_86;
        io_diffCommits_commitValid_87 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_87;
        io_diffCommits_commitValid_88 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_88;
        io_diffCommits_commitValid_89 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_89;
        io_diffCommits_commitValid_90 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_90;
        io_diffCommits_commitValid_91 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_91;
        io_diffCommits_commitValid_92 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_92;
        io_diffCommits_commitValid_93 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_93;
        io_diffCommits_commitValid_94 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_94;
        io_diffCommits_commitValid_95 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_95;
        io_diffCommits_commitValid_96 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_96;
        io_diffCommits_commitValid_97 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_97;
        io_diffCommits_commitValid_98 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_98;
        io_diffCommits_commitValid_99 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_99;
        io_diffCommits_commitValid_100 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_100;
        io_diffCommits_commitValid_101 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_101;
        io_diffCommits_commitValid_102 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_102;
        io_diffCommits_commitValid_103 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_103;
        io_diffCommits_commitValid_104 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_104;
        io_diffCommits_commitValid_105 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_105;
        io_diffCommits_commitValid_106 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_106;
        io_diffCommits_commitValid_107 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_107;
        io_diffCommits_commitValid_108 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_108;
        io_diffCommits_commitValid_109 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_109;
        io_diffCommits_commitValid_110 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_110;
        io_diffCommits_commitValid_111 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_111;
        io_diffCommits_commitValid_112 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_112;
        io_diffCommits_commitValid_113 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_113;
        io_diffCommits_commitValid_114 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_114;
        io_diffCommits_commitValid_115 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_115;
        io_diffCommits_commitValid_116 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_116;
        io_diffCommits_commitValid_117 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_117;
        io_diffCommits_commitValid_118 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_118;
        io_diffCommits_commitValid_119 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_119;
        io_diffCommits_commitValid_120 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_120;
        io_diffCommits_commitValid_121 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_121;
        io_diffCommits_commitValid_122 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_122;
        io_diffCommits_commitValid_123 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_123;
        io_diffCommits_commitValid_124 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_124;
        io_diffCommits_commitValid_125 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_125;
        io_diffCommits_commitValid_126 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_126;
        io_diffCommits_commitValid_127 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_127;
        io_diffCommits_commitValid_128 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_128;
        io_diffCommits_commitValid_129 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_129;
        io_diffCommits_commitValid_130 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_130;
        io_diffCommits_commitValid_131 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_131;
        io_diffCommits_commitValid_132 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_132;
        io_diffCommits_commitValid_133 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_133;
        io_diffCommits_commitValid_134 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_134;
        io_diffCommits_commitValid_135 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_135;
        io_diffCommits_commitValid_136 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_136;
        io_diffCommits_commitValid_137 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_137;
        io_diffCommits_commitValid_138 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_138;
        io_diffCommits_commitValid_139 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_139;
        io_diffCommits_commitValid_140 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_140;
        io_diffCommits_commitValid_141 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_141;
        io_diffCommits_commitValid_142 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_142;
        io_diffCommits_commitValid_143 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_143;
        io_diffCommits_commitValid_144 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_144;
        io_diffCommits_commitValid_145 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_145;
        io_diffCommits_commitValid_146 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_146;
        io_diffCommits_commitValid_147 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_147;
        io_diffCommits_commitValid_148 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_148;
        io_diffCommits_commitValid_149 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_149;
        io_diffCommits_commitValid_150 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_150;
        io_diffCommits_commitValid_151 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_151;
        io_diffCommits_commitValid_152 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_152;
        io_diffCommits_commitValid_153 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_153;
        io_diffCommits_commitValid_154 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_154;
        io_diffCommits_commitValid_155 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_155;
        io_diffCommits_commitValid_156 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_156;
        io_diffCommits_commitValid_157 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_157;
        io_diffCommits_commitValid_158 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_158;
        io_diffCommits_commitValid_159 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_159;
        io_diffCommits_commitValid_160 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_160;
        io_diffCommits_commitValid_161 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_161;
        io_diffCommits_commitValid_162 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_162;
        io_diffCommits_commitValid_163 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_163;
        io_diffCommits_commitValid_164 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_164;
        io_diffCommits_commitValid_165 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_165;
        io_diffCommits_commitValid_166 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_166;
        io_diffCommits_commitValid_167 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_167;
        io_diffCommits_commitValid_168 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_168;
        io_diffCommits_commitValid_169 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_169;
        io_diffCommits_commitValid_170 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_170;
        io_diffCommits_commitValid_171 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_171;
        io_diffCommits_commitValid_172 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_172;
        io_diffCommits_commitValid_173 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_173;
        io_diffCommits_commitValid_174 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_174;
        io_diffCommits_commitValid_175 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_175;
        io_diffCommits_commitValid_176 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_176;
        io_diffCommits_commitValid_177 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_177;
        io_diffCommits_commitValid_178 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_178;
        io_diffCommits_commitValid_179 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_179;
        io_diffCommits_commitValid_180 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_180;
        io_diffCommits_commitValid_181 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_181;
        io_diffCommits_commitValid_182 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_182;
        io_diffCommits_commitValid_183 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_183;
        io_diffCommits_commitValid_184 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_184;
        io_diffCommits_commitValid_185 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_185;
        io_diffCommits_commitValid_186 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_186;
        io_diffCommits_commitValid_187 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_187;
        io_diffCommits_commitValid_188 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_188;
        io_diffCommits_commitValid_189 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_189;
        io_diffCommits_commitValid_190 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_190;
        io_diffCommits_commitValid_191 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_191;
        io_diffCommits_commitValid_192 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_192;
        io_diffCommits_commitValid_193 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_193;
        io_diffCommits_commitValid_194 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_194;
        io_diffCommits_commitValid_195 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_195;
        io_diffCommits_commitValid_196 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_196;
        io_diffCommits_commitValid_197 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_197;
        io_diffCommits_commitValid_198 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_198;
        io_diffCommits_commitValid_199 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_199;
        io_diffCommits_commitValid_200 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_200;
        io_diffCommits_commitValid_201 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_201;
        io_diffCommits_commitValid_202 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_202;
        io_diffCommits_commitValid_203 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_203;
        io_diffCommits_commitValid_204 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_204;
        io_diffCommits_commitValid_205 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_205;
        io_diffCommits_commitValid_206 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_206;
        io_diffCommits_commitValid_207 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_207;
        io_diffCommits_commitValid_208 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_208;
        io_diffCommits_commitValid_209 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_209;
        io_diffCommits_commitValid_210 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_210;
        io_diffCommits_commitValid_211 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_211;
        io_diffCommits_commitValid_212 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_212;
        io_diffCommits_commitValid_213 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_213;
        io_diffCommits_commitValid_214 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_214;
        io_diffCommits_commitValid_215 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_215;
        io_diffCommits_commitValid_216 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_216;
        io_diffCommits_commitValid_217 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_217;
        io_diffCommits_commitValid_218 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_218;
        io_diffCommits_commitValid_219 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_219;
        io_diffCommits_commitValid_220 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_220;
        io_diffCommits_commitValid_221 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_221;
        io_diffCommits_commitValid_222 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_222;
        io_diffCommits_commitValid_223 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_223;
        io_diffCommits_commitValid_224 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_224;
        io_diffCommits_commitValid_225 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_225;
        io_diffCommits_commitValid_226 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_226;
        io_diffCommits_commitValid_227 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_227;
        io_diffCommits_commitValid_228 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_228;
        io_diffCommits_commitValid_229 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_229;
        io_diffCommits_commitValid_230 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_230;
        io_diffCommits_commitValid_231 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_231;
        io_diffCommits_commitValid_232 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_232;
        io_diffCommits_commitValid_233 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_233;
        io_diffCommits_commitValid_234 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_234;
        io_diffCommits_commitValid_235 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_235;
        io_diffCommits_commitValid_236 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_236;
        io_diffCommits_commitValid_237 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_237;
        io_diffCommits_commitValid_238 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_238;
        io_diffCommits_commitValid_239 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_239;
        io_diffCommits_commitValid_240 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_240;
        io_diffCommits_commitValid_241 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_241;
        io_diffCommits_commitValid_242 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_242;
        io_diffCommits_commitValid_243 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_243;
        io_diffCommits_commitValid_244 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_244;
        io_diffCommits_commitValid_245 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_245;
        io_diffCommits_commitValid_246 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_246;
        io_diffCommits_commitValid_247 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_247;
        io_diffCommits_commitValid_248 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_248;
        io_diffCommits_commitValid_249 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_249;
        io_diffCommits_commitValid_250 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_250;
        io_diffCommits_commitValid_251 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_251;
        io_diffCommits_commitValid_252 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_252;
        io_diffCommits_commitValid_253 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_253;
        io_diffCommits_commitValid_254 = this.vif.mon_mp.mon_cb.io_diffCommits_commitValid_254;
        io_diffCommits_info_0_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_0_ldest;
        io_diffCommits_info_0_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_0_pdest;
        io_diffCommits_info_0_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_0_rfWen;
        io_diffCommits_info_0_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_0_fpWen;
        io_diffCommits_info_0_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_0_vecWen;
        io_diffCommits_info_0_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_0_v0Wen;
        io_diffCommits_info_0_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_0_vlWen;
        io_diffCommits_info_1_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_1_ldest;
        io_diffCommits_info_1_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_1_pdest;
        io_diffCommits_info_1_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_1_rfWen;
        io_diffCommits_info_1_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_1_fpWen;
        io_diffCommits_info_1_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_1_vecWen;
        io_diffCommits_info_1_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_1_v0Wen;
        io_diffCommits_info_1_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_1_vlWen;
        io_diffCommits_info_2_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_2_ldest;
        io_diffCommits_info_2_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_2_pdest;
        io_diffCommits_info_2_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_2_rfWen;
        io_diffCommits_info_2_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_2_fpWen;
        io_diffCommits_info_2_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_2_vecWen;
        io_diffCommits_info_2_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_2_v0Wen;
        io_diffCommits_info_2_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_2_vlWen;
        io_diffCommits_info_3_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_3_ldest;
        io_diffCommits_info_3_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_3_pdest;
        io_diffCommits_info_3_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_3_rfWen;
        io_diffCommits_info_3_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_3_fpWen;
        io_diffCommits_info_3_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_3_vecWen;
        io_diffCommits_info_3_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_3_v0Wen;
        io_diffCommits_info_3_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_3_vlWen;
        io_diffCommits_info_4_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_4_ldest;
        io_diffCommits_info_4_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_4_pdest;
        io_diffCommits_info_4_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_4_rfWen;
        io_diffCommits_info_4_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_4_fpWen;
        io_diffCommits_info_4_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_4_vecWen;
        io_diffCommits_info_4_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_4_v0Wen;
        io_diffCommits_info_4_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_4_vlWen;
        io_diffCommits_info_5_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_5_ldest;
        io_diffCommits_info_5_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_5_pdest;
        io_diffCommits_info_5_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_5_rfWen;
        io_diffCommits_info_5_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_5_fpWen;
        io_diffCommits_info_5_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_5_vecWen;
        io_diffCommits_info_5_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_5_v0Wen;
        io_diffCommits_info_5_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_5_vlWen;
        io_diffCommits_info_6_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_6_ldest;
        io_diffCommits_info_6_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_6_pdest;
        io_diffCommits_info_6_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_6_rfWen;
        io_diffCommits_info_6_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_6_fpWen;
        io_diffCommits_info_6_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_6_vecWen;
        io_diffCommits_info_6_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_6_v0Wen;
        io_diffCommits_info_6_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_6_vlWen;
        io_diffCommits_info_7_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_7_ldest;
        io_diffCommits_info_7_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_7_pdest;
        io_diffCommits_info_7_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_7_rfWen;
        io_diffCommits_info_7_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_7_fpWen;
        io_diffCommits_info_7_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_7_vecWen;
        io_diffCommits_info_7_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_7_v0Wen;
        io_diffCommits_info_7_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_7_vlWen;
        io_diffCommits_info_8_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_8_ldest;
        io_diffCommits_info_8_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_8_pdest;
        io_diffCommits_info_8_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_8_rfWen;
        io_diffCommits_info_8_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_8_fpWen;
        io_diffCommits_info_8_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_8_vecWen;
        io_diffCommits_info_8_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_8_v0Wen;
        io_diffCommits_info_8_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_8_vlWen;
        io_diffCommits_info_9_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_9_ldest;
        io_diffCommits_info_9_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_9_pdest;
        io_diffCommits_info_9_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_9_rfWen;
        io_diffCommits_info_9_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_9_fpWen;
        io_diffCommits_info_9_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_9_vecWen;
        io_diffCommits_info_9_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_9_v0Wen;
        io_diffCommits_info_9_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_9_vlWen;
        io_diffCommits_info_10_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_10_ldest;
        io_diffCommits_info_10_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_10_pdest;
        io_diffCommits_info_10_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_10_rfWen;
        io_diffCommits_info_10_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_10_fpWen;
        io_diffCommits_info_10_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_10_vecWen;
        io_diffCommits_info_10_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_10_v0Wen;
        io_diffCommits_info_10_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_10_vlWen;
        io_diffCommits_info_11_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_11_ldest;
        io_diffCommits_info_11_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_11_pdest;
        io_diffCommits_info_11_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_11_rfWen;
        io_diffCommits_info_11_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_11_fpWen;
        io_diffCommits_info_11_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_11_vecWen;
        io_diffCommits_info_11_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_11_v0Wen;
        io_diffCommits_info_11_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_11_vlWen;
        io_diffCommits_info_12_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_12_ldest;
        io_diffCommits_info_12_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_12_pdest;
        io_diffCommits_info_12_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_12_rfWen;
        io_diffCommits_info_12_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_12_fpWen;
        io_diffCommits_info_12_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_12_vecWen;
        io_diffCommits_info_12_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_12_v0Wen;
        io_diffCommits_info_12_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_12_vlWen;
        io_diffCommits_info_13_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_13_ldest;
        io_diffCommits_info_13_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_13_pdest;
        io_diffCommits_info_13_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_13_rfWen;
        io_diffCommits_info_13_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_13_fpWen;
        io_diffCommits_info_13_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_13_vecWen;
        io_diffCommits_info_13_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_13_v0Wen;
        io_diffCommits_info_13_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_13_vlWen;
        io_diffCommits_info_14_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_14_ldest;
        io_diffCommits_info_14_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_14_pdest;
        io_diffCommits_info_14_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_14_rfWen;
        io_diffCommits_info_14_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_14_fpWen;
        io_diffCommits_info_14_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_14_vecWen;
        io_diffCommits_info_14_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_14_v0Wen;
        io_diffCommits_info_14_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_14_vlWen;
        io_diffCommits_info_15_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_15_ldest;
        io_diffCommits_info_15_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_15_pdest;
        io_diffCommits_info_15_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_15_rfWen;
        io_diffCommits_info_15_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_15_fpWen;
        io_diffCommits_info_15_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_15_vecWen;
        io_diffCommits_info_15_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_15_v0Wen;
        io_diffCommits_info_15_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_15_vlWen;
        io_diffCommits_info_16_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_16_ldest;
        io_diffCommits_info_16_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_16_pdest;
        io_diffCommits_info_16_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_16_rfWen;
        io_diffCommits_info_16_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_16_fpWen;
        io_diffCommits_info_16_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_16_vecWen;
        io_diffCommits_info_16_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_16_v0Wen;
        io_diffCommits_info_16_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_16_vlWen;
        io_diffCommits_info_17_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_17_ldest;
        io_diffCommits_info_17_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_17_pdest;
        io_diffCommits_info_17_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_17_rfWen;
        io_diffCommits_info_17_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_17_fpWen;
        io_diffCommits_info_17_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_17_vecWen;
        io_diffCommits_info_17_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_17_v0Wen;
        io_diffCommits_info_17_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_17_vlWen;
        io_diffCommits_info_18_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_18_ldest;
        io_diffCommits_info_18_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_18_pdest;
        io_diffCommits_info_18_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_18_rfWen;
        io_diffCommits_info_18_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_18_fpWen;
        io_diffCommits_info_18_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_18_vecWen;
        io_diffCommits_info_18_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_18_v0Wen;
        io_diffCommits_info_18_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_18_vlWen;
        io_diffCommits_info_19_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_19_ldest;
        io_diffCommits_info_19_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_19_pdest;
        io_diffCommits_info_19_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_19_rfWen;
        io_diffCommits_info_19_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_19_fpWen;
        io_diffCommits_info_19_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_19_vecWen;
        io_diffCommits_info_19_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_19_v0Wen;
        io_diffCommits_info_19_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_19_vlWen;
        io_diffCommits_info_20_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_20_ldest;
        io_diffCommits_info_20_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_20_pdest;
        io_diffCommits_info_20_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_20_rfWen;
        io_diffCommits_info_20_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_20_fpWen;
        io_diffCommits_info_20_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_20_vecWen;
        io_diffCommits_info_20_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_20_v0Wen;
        io_diffCommits_info_20_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_20_vlWen;
        io_diffCommits_info_21_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_21_ldest;
        io_diffCommits_info_21_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_21_pdest;
        io_diffCommits_info_21_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_21_rfWen;
        io_diffCommits_info_21_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_21_fpWen;
        io_diffCommits_info_21_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_21_vecWen;
        io_diffCommits_info_21_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_21_v0Wen;
        io_diffCommits_info_21_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_21_vlWen;
        io_diffCommits_info_22_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_22_ldest;
        io_diffCommits_info_22_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_22_pdest;
        io_diffCommits_info_22_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_22_rfWen;
        io_diffCommits_info_22_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_22_fpWen;
        io_diffCommits_info_22_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_22_vecWen;
        io_diffCommits_info_22_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_22_v0Wen;
        io_diffCommits_info_22_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_22_vlWen;
        io_diffCommits_info_23_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_23_ldest;
        io_diffCommits_info_23_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_23_pdest;
        io_diffCommits_info_23_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_23_rfWen;
        io_diffCommits_info_23_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_23_fpWen;
        io_diffCommits_info_23_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_23_vecWen;
        io_diffCommits_info_23_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_23_v0Wen;
        io_diffCommits_info_23_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_23_vlWen;
        io_diffCommits_info_24_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_24_ldest;
        io_diffCommits_info_24_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_24_pdest;
        io_diffCommits_info_24_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_24_rfWen;
        io_diffCommits_info_24_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_24_fpWen;
        io_diffCommits_info_24_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_24_vecWen;
        io_diffCommits_info_24_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_24_v0Wen;
        io_diffCommits_info_24_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_24_vlWen;
        io_diffCommits_info_25_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_25_ldest;
        io_diffCommits_info_25_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_25_pdest;
        io_diffCommits_info_25_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_25_rfWen;
        io_diffCommits_info_25_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_25_fpWen;
        io_diffCommits_info_25_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_25_vecWen;
        io_diffCommits_info_25_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_25_v0Wen;
        io_diffCommits_info_25_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_25_vlWen;
        io_diffCommits_info_26_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_26_ldest;
        io_diffCommits_info_26_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_26_pdest;
        io_diffCommits_info_26_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_26_rfWen;
        io_diffCommits_info_26_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_26_fpWen;
        io_diffCommits_info_26_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_26_vecWen;
        io_diffCommits_info_26_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_26_v0Wen;
        io_diffCommits_info_26_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_26_vlWen;
        io_diffCommits_info_27_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_27_ldest;
        io_diffCommits_info_27_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_27_pdest;
        io_diffCommits_info_27_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_27_rfWen;
        io_diffCommits_info_27_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_27_fpWen;
        io_diffCommits_info_27_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_27_vecWen;
        io_diffCommits_info_27_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_27_v0Wen;
        io_diffCommits_info_27_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_27_vlWen;
        io_diffCommits_info_28_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_28_ldest;
        io_diffCommits_info_28_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_28_pdest;
        io_diffCommits_info_28_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_28_rfWen;
        io_diffCommits_info_28_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_28_fpWen;
        io_diffCommits_info_28_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_28_vecWen;
        io_diffCommits_info_28_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_28_v0Wen;
        io_diffCommits_info_28_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_28_vlWen;
        io_diffCommits_info_29_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_29_ldest;
        io_diffCommits_info_29_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_29_pdest;
        io_diffCommits_info_29_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_29_rfWen;
        io_diffCommits_info_29_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_29_fpWen;
        io_diffCommits_info_29_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_29_vecWen;
        io_diffCommits_info_29_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_29_v0Wen;
        io_diffCommits_info_29_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_29_vlWen;
        io_diffCommits_info_30_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_30_ldest;
        io_diffCommits_info_30_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_30_pdest;
        io_diffCommits_info_30_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_30_rfWen;
        io_diffCommits_info_30_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_30_fpWen;
        io_diffCommits_info_30_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_30_vecWen;
        io_diffCommits_info_30_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_30_v0Wen;
        io_diffCommits_info_30_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_30_vlWen;
        io_diffCommits_info_31_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_31_ldest;
        io_diffCommits_info_31_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_31_pdest;
        io_diffCommits_info_31_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_31_rfWen;
        io_diffCommits_info_31_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_31_fpWen;
        io_diffCommits_info_31_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_31_vecWen;
        io_diffCommits_info_31_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_31_v0Wen;
        io_diffCommits_info_31_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_31_vlWen;
        io_diffCommits_info_32_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_32_ldest;
        io_diffCommits_info_32_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_32_pdest;
        io_diffCommits_info_32_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_32_rfWen;
        io_diffCommits_info_32_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_32_fpWen;
        io_diffCommits_info_32_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_32_vecWen;
        io_diffCommits_info_32_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_32_v0Wen;
        io_diffCommits_info_32_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_32_vlWen;
        io_diffCommits_info_33_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_33_ldest;
        io_diffCommits_info_33_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_33_pdest;
        io_diffCommits_info_33_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_33_rfWen;
        io_diffCommits_info_33_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_33_fpWen;
        io_diffCommits_info_33_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_33_vecWen;
        io_diffCommits_info_33_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_33_v0Wen;
        io_diffCommits_info_33_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_33_vlWen;
        io_diffCommits_info_34_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_34_ldest;
        io_diffCommits_info_34_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_34_pdest;
        io_diffCommits_info_34_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_34_rfWen;
        io_diffCommits_info_34_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_34_fpWen;
        io_diffCommits_info_34_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_34_vecWen;
        io_diffCommits_info_34_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_34_v0Wen;
        io_diffCommits_info_34_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_34_vlWen;
        io_diffCommits_info_35_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_35_ldest;
        io_diffCommits_info_35_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_35_pdest;
        io_diffCommits_info_35_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_35_rfWen;
        io_diffCommits_info_35_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_35_fpWen;
        io_diffCommits_info_35_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_35_vecWen;
        io_diffCommits_info_35_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_35_v0Wen;
        io_diffCommits_info_35_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_35_vlWen;
        io_diffCommits_info_36_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_36_ldest;
        io_diffCommits_info_36_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_36_pdest;
        io_diffCommits_info_36_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_36_rfWen;
        io_diffCommits_info_36_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_36_fpWen;
        io_diffCommits_info_36_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_36_vecWen;
        io_diffCommits_info_36_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_36_v0Wen;
        io_diffCommits_info_36_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_36_vlWen;
        io_diffCommits_info_37_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_37_ldest;
        io_diffCommits_info_37_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_37_pdest;
        io_diffCommits_info_37_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_37_rfWen;
        io_diffCommits_info_37_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_37_fpWen;
        io_diffCommits_info_37_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_37_vecWen;
        io_diffCommits_info_37_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_37_v0Wen;
        io_diffCommits_info_37_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_37_vlWen;
        io_diffCommits_info_38_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_38_ldest;
        io_diffCommits_info_38_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_38_pdest;
        io_diffCommits_info_38_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_38_rfWen;
        io_diffCommits_info_38_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_38_fpWen;
        io_diffCommits_info_38_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_38_vecWen;
        io_diffCommits_info_38_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_38_v0Wen;
        io_diffCommits_info_38_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_38_vlWen;
        io_diffCommits_info_39_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_39_ldest;
        io_diffCommits_info_39_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_39_pdest;
        io_diffCommits_info_39_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_39_rfWen;
        io_diffCommits_info_39_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_39_fpWen;
        io_diffCommits_info_39_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_39_vecWen;
        io_diffCommits_info_39_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_39_v0Wen;
        io_diffCommits_info_39_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_39_vlWen;
        io_diffCommits_info_40_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_40_ldest;
        io_diffCommits_info_40_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_40_pdest;
        io_diffCommits_info_40_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_40_rfWen;
        io_diffCommits_info_40_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_40_fpWen;
        io_diffCommits_info_40_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_40_vecWen;
        io_diffCommits_info_40_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_40_v0Wen;
        io_diffCommits_info_40_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_40_vlWen;
        io_diffCommits_info_41_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_41_ldest;
        io_diffCommits_info_41_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_41_pdest;
        io_diffCommits_info_41_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_41_rfWen;
        io_diffCommits_info_41_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_41_fpWen;
        io_diffCommits_info_41_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_41_vecWen;
        io_diffCommits_info_41_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_41_v0Wen;
        io_diffCommits_info_41_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_41_vlWen;
        io_diffCommits_info_42_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_42_ldest;
        io_diffCommits_info_42_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_42_pdest;
        io_diffCommits_info_42_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_42_rfWen;
        io_diffCommits_info_42_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_42_fpWen;
        io_diffCommits_info_42_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_42_vecWen;
        io_diffCommits_info_42_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_42_v0Wen;
        io_diffCommits_info_42_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_42_vlWen;
        io_diffCommits_info_43_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_43_ldest;
        io_diffCommits_info_43_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_43_pdest;
        io_diffCommits_info_43_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_43_rfWen;
        io_diffCommits_info_43_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_43_fpWen;
        io_diffCommits_info_43_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_43_vecWen;
        io_diffCommits_info_43_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_43_v0Wen;
        io_diffCommits_info_43_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_43_vlWen;
        io_diffCommits_info_44_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_44_ldest;
        io_diffCommits_info_44_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_44_pdest;
        io_diffCommits_info_44_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_44_rfWen;
        io_diffCommits_info_44_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_44_fpWen;
        io_diffCommits_info_44_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_44_vecWen;
        io_diffCommits_info_44_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_44_v0Wen;
        io_diffCommits_info_44_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_44_vlWen;
        io_diffCommits_info_45_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_45_ldest;
        io_diffCommits_info_45_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_45_pdest;
        io_diffCommits_info_45_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_45_rfWen;
        io_diffCommits_info_45_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_45_fpWen;
        io_diffCommits_info_45_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_45_vecWen;
        io_diffCommits_info_45_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_45_v0Wen;
        io_diffCommits_info_45_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_45_vlWen;
        io_diffCommits_info_46_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_46_ldest;
        io_diffCommits_info_46_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_46_pdest;
        io_diffCommits_info_46_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_46_rfWen;
        io_diffCommits_info_46_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_46_fpWen;
        io_diffCommits_info_46_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_46_vecWen;
        io_diffCommits_info_46_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_46_v0Wen;
        io_diffCommits_info_46_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_46_vlWen;
        io_diffCommits_info_47_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_47_ldest;
        io_diffCommits_info_47_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_47_pdest;
        io_diffCommits_info_47_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_47_rfWen;
        io_diffCommits_info_47_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_47_fpWen;
        io_diffCommits_info_47_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_47_vecWen;
        io_diffCommits_info_47_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_47_v0Wen;
        io_diffCommits_info_47_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_47_vlWen;
        io_diffCommits_info_48_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_48_ldest;
        io_diffCommits_info_48_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_48_pdest;
        io_diffCommits_info_48_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_48_rfWen;
        io_diffCommits_info_48_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_48_fpWen;
        io_diffCommits_info_48_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_48_vecWen;
        io_diffCommits_info_48_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_48_v0Wen;
        io_diffCommits_info_48_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_48_vlWen;
        io_diffCommits_info_49_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_49_ldest;
        io_diffCommits_info_49_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_49_pdest;
        io_diffCommits_info_49_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_49_rfWen;
        io_diffCommits_info_49_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_49_fpWen;
        io_diffCommits_info_49_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_49_vecWen;
        io_diffCommits_info_49_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_49_v0Wen;
        io_diffCommits_info_49_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_49_vlWen;
        io_diffCommits_info_50_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_50_ldest;
        io_diffCommits_info_50_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_50_pdest;
        io_diffCommits_info_50_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_50_rfWen;
        io_diffCommits_info_50_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_50_fpWen;
        io_diffCommits_info_50_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_50_vecWen;
        io_diffCommits_info_50_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_50_v0Wen;
        io_diffCommits_info_50_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_50_vlWen;
        io_diffCommits_info_51_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_51_ldest;
        io_diffCommits_info_51_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_51_pdest;
        io_diffCommits_info_51_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_51_rfWen;
        io_diffCommits_info_51_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_51_fpWen;
        io_diffCommits_info_51_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_51_vecWen;
        io_diffCommits_info_51_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_51_v0Wen;
        io_diffCommits_info_51_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_51_vlWen;
        io_diffCommits_info_52_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_52_ldest;
        io_diffCommits_info_52_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_52_pdest;
        io_diffCommits_info_52_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_52_rfWen;
        io_diffCommits_info_52_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_52_fpWen;
        io_diffCommits_info_52_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_52_vecWen;
        io_diffCommits_info_52_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_52_v0Wen;
        io_diffCommits_info_52_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_52_vlWen;
        io_diffCommits_info_53_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_53_ldest;
        io_diffCommits_info_53_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_53_pdest;
        io_diffCommits_info_53_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_53_rfWen;
        io_diffCommits_info_53_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_53_fpWen;
        io_diffCommits_info_53_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_53_vecWen;
        io_diffCommits_info_53_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_53_v0Wen;
        io_diffCommits_info_53_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_53_vlWen;
        io_diffCommits_info_54_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_54_ldest;
        io_diffCommits_info_54_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_54_pdest;
        io_diffCommits_info_54_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_54_rfWen;
        io_diffCommits_info_54_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_54_fpWen;
        io_diffCommits_info_54_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_54_vecWen;
        io_diffCommits_info_54_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_54_v0Wen;
        io_diffCommits_info_54_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_54_vlWen;
        io_diffCommits_info_55_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_55_ldest;
        io_diffCommits_info_55_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_55_pdest;
        io_diffCommits_info_55_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_55_rfWen;
        io_diffCommits_info_55_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_55_fpWen;
        io_diffCommits_info_55_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_55_vecWen;
        io_diffCommits_info_55_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_55_v0Wen;
        io_diffCommits_info_55_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_55_vlWen;
        io_diffCommits_info_56_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_56_ldest;
        io_diffCommits_info_56_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_56_pdest;
        io_diffCommits_info_56_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_56_rfWen;
        io_diffCommits_info_56_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_56_fpWen;
        io_diffCommits_info_56_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_56_vecWen;
        io_diffCommits_info_56_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_56_v0Wen;
        io_diffCommits_info_56_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_56_vlWen;
        io_diffCommits_info_57_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_57_ldest;
        io_diffCommits_info_57_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_57_pdest;
        io_diffCommits_info_57_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_57_rfWen;
        io_diffCommits_info_57_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_57_fpWen;
        io_diffCommits_info_57_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_57_vecWen;
        io_diffCommits_info_57_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_57_v0Wen;
        io_diffCommits_info_57_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_57_vlWen;
        io_diffCommits_info_58_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_58_ldest;
        io_diffCommits_info_58_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_58_pdest;
        io_diffCommits_info_58_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_58_rfWen;
        io_diffCommits_info_58_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_58_fpWen;
        io_diffCommits_info_58_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_58_vecWen;
        io_diffCommits_info_58_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_58_v0Wen;
        io_diffCommits_info_58_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_58_vlWen;
        io_diffCommits_info_59_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_59_ldest;
        io_diffCommits_info_59_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_59_pdest;
        io_diffCommits_info_59_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_59_rfWen;
        io_diffCommits_info_59_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_59_fpWen;
        io_diffCommits_info_59_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_59_vecWen;
        io_diffCommits_info_59_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_59_v0Wen;
        io_diffCommits_info_59_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_59_vlWen;
        io_diffCommits_info_60_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_60_ldest;
        io_diffCommits_info_60_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_60_pdest;
        io_diffCommits_info_60_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_60_rfWen;
        io_diffCommits_info_60_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_60_fpWen;
        io_diffCommits_info_60_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_60_vecWen;
        io_diffCommits_info_60_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_60_v0Wen;
        io_diffCommits_info_60_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_60_vlWen;
        io_diffCommits_info_61_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_61_ldest;
        io_diffCommits_info_61_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_61_pdest;
        io_diffCommits_info_61_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_61_rfWen;
        io_diffCommits_info_61_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_61_fpWen;
        io_diffCommits_info_61_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_61_vecWen;
        io_diffCommits_info_61_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_61_v0Wen;
        io_diffCommits_info_61_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_61_vlWen;
        io_diffCommits_info_62_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_62_ldest;
        io_diffCommits_info_62_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_62_pdest;
        io_diffCommits_info_62_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_62_rfWen;
        io_diffCommits_info_62_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_62_fpWen;
        io_diffCommits_info_62_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_62_vecWen;
        io_diffCommits_info_62_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_62_v0Wen;
        io_diffCommits_info_62_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_62_vlWen;
        io_diffCommits_info_63_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_63_ldest;
        io_diffCommits_info_63_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_63_pdest;
        io_diffCommits_info_63_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_63_rfWen;
        io_diffCommits_info_63_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_63_fpWen;
        io_diffCommits_info_63_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_63_vecWen;
        io_diffCommits_info_63_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_63_v0Wen;
        io_diffCommits_info_63_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_63_vlWen;
        io_diffCommits_info_64_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_64_ldest;
        io_diffCommits_info_64_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_64_pdest;
        io_diffCommits_info_64_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_64_rfWen;
        io_diffCommits_info_64_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_64_fpWen;
        io_diffCommits_info_64_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_64_vecWen;
        io_diffCommits_info_64_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_64_v0Wen;
        io_diffCommits_info_64_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_64_vlWen;
        io_diffCommits_info_65_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_65_ldest;
        io_diffCommits_info_65_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_65_pdest;
        io_diffCommits_info_65_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_65_rfWen;
        io_diffCommits_info_65_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_65_fpWen;
        io_diffCommits_info_65_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_65_vecWen;
        io_diffCommits_info_65_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_65_v0Wen;
        io_diffCommits_info_65_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_65_vlWen;
        io_diffCommits_info_66_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_66_ldest;
        io_diffCommits_info_66_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_66_pdest;
        io_diffCommits_info_66_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_66_rfWen;
        io_diffCommits_info_66_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_66_fpWen;
        io_diffCommits_info_66_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_66_vecWen;
        io_diffCommits_info_66_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_66_v0Wen;
        io_diffCommits_info_66_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_66_vlWen;
        io_diffCommits_info_67_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_67_ldest;
        io_diffCommits_info_67_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_67_pdest;
        io_diffCommits_info_67_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_67_rfWen;
        io_diffCommits_info_67_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_67_fpWen;
        io_diffCommits_info_67_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_67_vecWen;
        io_diffCommits_info_67_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_67_v0Wen;
        io_diffCommits_info_67_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_67_vlWen;
        io_diffCommits_info_68_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_68_ldest;
        io_diffCommits_info_68_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_68_pdest;
        io_diffCommits_info_68_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_68_rfWen;
        io_diffCommits_info_68_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_68_fpWen;
        io_diffCommits_info_68_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_68_vecWen;
        io_diffCommits_info_68_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_68_v0Wen;
        io_diffCommits_info_68_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_68_vlWen;
        io_diffCommits_info_69_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_69_ldest;
        io_diffCommits_info_69_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_69_pdest;
        io_diffCommits_info_69_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_69_rfWen;
        io_diffCommits_info_69_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_69_fpWen;
        io_diffCommits_info_69_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_69_vecWen;
        io_diffCommits_info_69_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_69_v0Wen;
        io_diffCommits_info_69_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_69_vlWen;
        io_diffCommits_info_70_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_70_ldest;
        io_diffCommits_info_70_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_70_pdest;
        io_diffCommits_info_70_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_70_rfWen;
        io_diffCommits_info_70_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_70_fpWen;
        io_diffCommits_info_70_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_70_vecWen;
        io_diffCommits_info_70_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_70_v0Wen;
        io_diffCommits_info_70_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_70_vlWen;
        io_diffCommits_info_71_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_71_ldest;
        io_diffCommits_info_71_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_71_pdest;
        io_diffCommits_info_71_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_71_rfWen;
        io_diffCommits_info_71_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_71_fpWen;
        io_diffCommits_info_71_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_71_vecWen;
        io_diffCommits_info_71_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_71_v0Wen;
        io_diffCommits_info_71_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_71_vlWen;
        io_diffCommits_info_72_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_72_ldest;
        io_diffCommits_info_72_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_72_pdest;
        io_diffCommits_info_72_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_72_rfWen;
        io_diffCommits_info_72_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_72_fpWen;
        io_diffCommits_info_72_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_72_vecWen;
        io_diffCommits_info_72_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_72_v0Wen;
        io_diffCommits_info_72_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_72_vlWen;
        io_diffCommits_info_73_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_73_ldest;
        io_diffCommits_info_73_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_73_pdest;
        io_diffCommits_info_73_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_73_rfWen;
        io_diffCommits_info_73_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_73_fpWen;
        io_diffCommits_info_73_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_73_vecWen;
        io_diffCommits_info_73_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_73_v0Wen;
        io_diffCommits_info_73_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_73_vlWen;
        io_diffCommits_info_74_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_74_ldest;
        io_diffCommits_info_74_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_74_pdest;
        io_diffCommits_info_74_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_74_rfWen;
        io_diffCommits_info_74_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_74_fpWen;
        io_diffCommits_info_74_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_74_vecWen;
        io_diffCommits_info_74_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_74_v0Wen;
        io_diffCommits_info_74_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_74_vlWen;
        io_diffCommits_info_75_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_75_ldest;
        io_diffCommits_info_75_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_75_pdest;
        io_diffCommits_info_75_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_75_rfWen;
        io_diffCommits_info_75_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_75_fpWen;
        io_diffCommits_info_75_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_75_vecWen;
        io_diffCommits_info_75_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_75_v0Wen;
        io_diffCommits_info_75_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_75_vlWen;
        io_diffCommits_info_76_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_76_ldest;
        io_diffCommits_info_76_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_76_pdest;
        io_diffCommits_info_76_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_76_rfWen;
        io_diffCommits_info_76_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_76_fpWen;
        io_diffCommits_info_76_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_76_vecWen;
        io_diffCommits_info_76_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_76_v0Wen;
        io_diffCommits_info_76_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_76_vlWen;
        io_diffCommits_info_77_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_77_ldest;
        io_diffCommits_info_77_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_77_pdest;
        io_diffCommits_info_77_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_77_rfWen;
        io_diffCommits_info_77_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_77_fpWen;
        io_diffCommits_info_77_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_77_vecWen;
        io_diffCommits_info_77_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_77_v0Wen;
        io_diffCommits_info_77_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_77_vlWen;
        io_diffCommits_info_78_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_78_ldest;
        io_diffCommits_info_78_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_78_pdest;
        io_diffCommits_info_78_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_78_rfWen;
        io_diffCommits_info_78_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_78_fpWen;
        io_diffCommits_info_78_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_78_vecWen;
        io_diffCommits_info_78_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_78_v0Wen;
        io_diffCommits_info_78_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_78_vlWen;
        io_diffCommits_info_79_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_79_ldest;
        io_diffCommits_info_79_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_79_pdest;
        io_diffCommits_info_79_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_79_rfWen;
        io_diffCommits_info_79_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_79_fpWen;
        io_diffCommits_info_79_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_79_vecWen;
        io_diffCommits_info_79_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_79_v0Wen;
        io_diffCommits_info_79_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_79_vlWen;
        io_diffCommits_info_80_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_80_ldest;
        io_diffCommits_info_80_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_80_pdest;
        io_diffCommits_info_80_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_80_rfWen;
        io_diffCommits_info_80_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_80_fpWen;
        io_diffCommits_info_80_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_80_vecWen;
        io_diffCommits_info_80_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_80_v0Wen;
        io_diffCommits_info_80_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_80_vlWen;
        io_diffCommits_info_81_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_81_ldest;
        io_diffCommits_info_81_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_81_pdest;
        io_diffCommits_info_81_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_81_rfWen;
        io_diffCommits_info_81_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_81_fpWen;
        io_diffCommits_info_81_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_81_vecWen;
        io_diffCommits_info_81_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_81_v0Wen;
        io_diffCommits_info_81_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_81_vlWen;
        io_diffCommits_info_82_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_82_ldest;
        io_diffCommits_info_82_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_82_pdest;
        io_diffCommits_info_82_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_82_rfWen;
        io_diffCommits_info_82_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_82_fpWen;
        io_diffCommits_info_82_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_82_vecWen;
        io_diffCommits_info_82_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_82_v0Wen;
        io_diffCommits_info_82_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_82_vlWen;
        io_diffCommits_info_83_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_83_ldest;
        io_diffCommits_info_83_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_83_pdest;
        io_diffCommits_info_83_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_83_rfWen;
        io_diffCommits_info_83_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_83_fpWen;
        io_diffCommits_info_83_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_83_vecWen;
        io_diffCommits_info_83_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_83_v0Wen;
        io_diffCommits_info_83_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_83_vlWen;
        io_diffCommits_info_84_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_84_ldest;
        io_diffCommits_info_84_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_84_pdest;
        io_diffCommits_info_84_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_84_rfWen;
        io_diffCommits_info_84_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_84_fpWen;
        io_diffCommits_info_84_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_84_vecWen;
        io_diffCommits_info_84_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_84_v0Wen;
        io_diffCommits_info_84_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_84_vlWen;
        io_diffCommits_info_85_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_85_ldest;
        io_diffCommits_info_85_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_85_pdest;
        io_diffCommits_info_85_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_85_rfWen;
        io_diffCommits_info_85_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_85_fpWen;
        io_diffCommits_info_85_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_85_vecWen;
        io_diffCommits_info_85_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_85_v0Wen;
        io_diffCommits_info_85_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_85_vlWen;
        io_diffCommits_info_86_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_86_ldest;
        io_diffCommits_info_86_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_86_pdest;
        io_diffCommits_info_86_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_86_rfWen;
        io_diffCommits_info_86_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_86_fpWen;
        io_diffCommits_info_86_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_86_vecWen;
        io_diffCommits_info_86_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_86_v0Wen;
        io_diffCommits_info_86_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_86_vlWen;
        io_diffCommits_info_87_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_87_ldest;
        io_diffCommits_info_87_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_87_pdest;
        io_diffCommits_info_87_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_87_rfWen;
        io_diffCommits_info_87_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_87_fpWen;
        io_diffCommits_info_87_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_87_vecWen;
        io_diffCommits_info_87_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_87_v0Wen;
        io_diffCommits_info_87_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_87_vlWen;
        io_diffCommits_info_88_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_88_ldest;
        io_diffCommits_info_88_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_88_pdest;
        io_diffCommits_info_88_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_88_rfWen;
        io_diffCommits_info_88_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_88_fpWen;
        io_diffCommits_info_88_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_88_vecWen;
        io_diffCommits_info_88_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_88_v0Wen;
        io_diffCommits_info_88_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_88_vlWen;
        io_diffCommits_info_89_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_89_ldest;
        io_diffCommits_info_89_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_89_pdest;
        io_diffCommits_info_89_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_89_rfWen;
        io_diffCommits_info_89_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_89_fpWen;
        io_diffCommits_info_89_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_89_vecWen;
        io_diffCommits_info_89_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_89_v0Wen;
        io_diffCommits_info_89_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_89_vlWen;
        io_diffCommits_info_90_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_90_ldest;
        io_diffCommits_info_90_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_90_pdest;
        io_diffCommits_info_90_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_90_rfWen;
        io_diffCommits_info_90_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_90_fpWen;
        io_diffCommits_info_90_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_90_vecWen;
        io_diffCommits_info_90_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_90_v0Wen;
        io_diffCommits_info_90_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_90_vlWen;
        io_diffCommits_info_91_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_91_ldest;
        io_diffCommits_info_91_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_91_pdest;
        io_diffCommits_info_91_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_91_rfWen;
        io_diffCommits_info_91_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_91_fpWen;
        io_diffCommits_info_91_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_91_vecWen;
        io_diffCommits_info_91_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_91_v0Wen;
        io_diffCommits_info_91_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_91_vlWen;
        io_diffCommits_info_92_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_92_ldest;
        io_diffCommits_info_92_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_92_pdest;
        io_diffCommits_info_92_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_92_rfWen;
        io_diffCommits_info_92_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_92_fpWen;
        io_diffCommits_info_92_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_92_vecWen;
        io_diffCommits_info_92_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_92_v0Wen;
        io_diffCommits_info_92_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_92_vlWen;
        io_diffCommits_info_93_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_93_ldest;
        io_diffCommits_info_93_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_93_pdest;
        io_diffCommits_info_93_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_93_rfWen;
        io_diffCommits_info_93_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_93_fpWen;
        io_diffCommits_info_93_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_93_vecWen;
        io_diffCommits_info_93_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_93_v0Wen;
        io_diffCommits_info_93_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_93_vlWen;
        io_diffCommits_info_94_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_94_ldest;
        io_diffCommits_info_94_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_94_pdest;
        io_diffCommits_info_94_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_94_rfWen;
        io_diffCommits_info_94_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_94_fpWen;
        io_diffCommits_info_94_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_94_vecWen;
        io_diffCommits_info_94_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_94_v0Wen;
        io_diffCommits_info_94_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_94_vlWen;
        io_diffCommits_info_95_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_95_ldest;
        io_diffCommits_info_95_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_95_pdest;
        io_diffCommits_info_95_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_95_rfWen;
        io_diffCommits_info_95_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_95_fpWen;
        io_diffCommits_info_95_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_95_vecWen;
        io_diffCommits_info_95_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_95_v0Wen;
        io_diffCommits_info_95_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_95_vlWen;
        io_diffCommits_info_96_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_96_ldest;
        io_diffCommits_info_96_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_96_pdest;
        io_diffCommits_info_96_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_96_rfWen;
        io_diffCommits_info_96_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_96_fpWen;
        io_diffCommits_info_96_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_96_vecWen;
        io_diffCommits_info_96_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_96_v0Wen;
        io_diffCommits_info_96_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_96_vlWen;
        io_diffCommits_info_97_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_97_ldest;
        io_diffCommits_info_97_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_97_pdest;
        io_diffCommits_info_97_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_97_rfWen;
        io_diffCommits_info_97_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_97_fpWen;
        io_diffCommits_info_97_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_97_vecWen;
        io_diffCommits_info_97_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_97_v0Wen;
        io_diffCommits_info_97_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_97_vlWen;
        io_diffCommits_info_98_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_98_ldest;
        io_diffCommits_info_98_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_98_pdest;
        io_diffCommits_info_98_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_98_rfWen;
        io_diffCommits_info_98_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_98_fpWen;
        io_diffCommits_info_98_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_98_vecWen;
        io_diffCommits_info_98_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_98_v0Wen;
        io_diffCommits_info_98_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_98_vlWen;
        io_diffCommits_info_99_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_99_ldest;
        io_diffCommits_info_99_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_99_pdest;
        io_diffCommits_info_99_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_99_rfWen;
        io_diffCommits_info_99_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_99_fpWen;
        io_diffCommits_info_99_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_99_vecWen;
        io_diffCommits_info_99_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_99_v0Wen;
        io_diffCommits_info_99_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_99_vlWen;
        io_diffCommits_info_100_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_100_ldest;
        io_diffCommits_info_100_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_100_pdest;
        io_diffCommits_info_100_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_100_rfWen;
        io_diffCommits_info_100_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_100_fpWen;
        io_diffCommits_info_100_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_100_vecWen;
        io_diffCommits_info_100_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_100_v0Wen;
        io_diffCommits_info_100_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_100_vlWen;
        io_diffCommits_info_101_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_101_ldest;
        io_diffCommits_info_101_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_101_pdest;
        io_diffCommits_info_101_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_101_rfWen;
        io_diffCommits_info_101_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_101_fpWen;
        io_diffCommits_info_101_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_101_vecWen;
        io_diffCommits_info_101_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_101_v0Wen;
        io_diffCommits_info_101_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_101_vlWen;
        io_diffCommits_info_102_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_102_ldest;
        io_diffCommits_info_102_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_102_pdest;
        io_diffCommits_info_102_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_102_rfWen;
        io_diffCommits_info_102_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_102_fpWen;
        io_diffCommits_info_102_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_102_vecWen;
        io_diffCommits_info_102_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_102_v0Wen;
        io_diffCommits_info_102_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_102_vlWen;
        io_diffCommits_info_103_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_103_ldest;
        io_diffCommits_info_103_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_103_pdest;
        io_diffCommits_info_103_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_103_rfWen;
        io_diffCommits_info_103_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_103_fpWen;
        io_diffCommits_info_103_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_103_vecWen;
        io_diffCommits_info_103_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_103_v0Wen;
        io_diffCommits_info_103_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_103_vlWen;
        io_diffCommits_info_104_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_104_ldest;
        io_diffCommits_info_104_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_104_pdest;
        io_diffCommits_info_104_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_104_rfWen;
        io_diffCommits_info_104_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_104_fpWen;
        io_diffCommits_info_104_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_104_vecWen;
        io_diffCommits_info_104_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_104_v0Wen;
        io_diffCommits_info_104_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_104_vlWen;
        io_diffCommits_info_105_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_105_ldest;
        io_diffCommits_info_105_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_105_pdest;
        io_diffCommits_info_105_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_105_rfWen;
        io_diffCommits_info_105_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_105_fpWen;
        io_diffCommits_info_105_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_105_vecWen;
        io_diffCommits_info_105_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_105_v0Wen;
        io_diffCommits_info_105_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_105_vlWen;
        io_diffCommits_info_106_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_106_ldest;
        io_diffCommits_info_106_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_106_pdest;
        io_diffCommits_info_106_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_106_rfWen;
        io_diffCommits_info_106_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_106_fpWen;
        io_diffCommits_info_106_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_106_vecWen;
        io_diffCommits_info_106_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_106_v0Wen;
        io_diffCommits_info_106_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_106_vlWen;
        io_diffCommits_info_107_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_107_ldest;
        io_diffCommits_info_107_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_107_pdest;
        io_diffCommits_info_107_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_107_rfWen;
        io_diffCommits_info_107_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_107_fpWen;
        io_diffCommits_info_107_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_107_vecWen;
        io_diffCommits_info_107_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_107_v0Wen;
        io_diffCommits_info_107_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_107_vlWen;
        io_diffCommits_info_108_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_108_ldest;
        io_diffCommits_info_108_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_108_pdest;
        io_diffCommits_info_108_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_108_rfWen;
        io_diffCommits_info_108_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_108_fpWen;
        io_diffCommits_info_108_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_108_vecWen;
        io_diffCommits_info_108_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_108_v0Wen;
        io_diffCommits_info_108_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_108_vlWen;
        io_diffCommits_info_109_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_109_ldest;
        io_diffCommits_info_109_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_109_pdest;
        io_diffCommits_info_109_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_109_rfWen;
        io_diffCommits_info_109_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_109_fpWen;
        io_diffCommits_info_109_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_109_vecWen;
        io_diffCommits_info_109_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_109_v0Wen;
        io_diffCommits_info_109_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_109_vlWen;
        io_diffCommits_info_110_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_110_ldest;
        io_diffCommits_info_110_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_110_pdest;
        io_diffCommits_info_110_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_110_rfWen;
        io_diffCommits_info_110_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_110_fpWen;
        io_diffCommits_info_110_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_110_vecWen;
        io_diffCommits_info_110_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_110_v0Wen;
        io_diffCommits_info_110_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_110_vlWen;
        io_diffCommits_info_111_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_111_ldest;
        io_diffCommits_info_111_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_111_pdest;
        io_diffCommits_info_111_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_111_rfWen;
        io_diffCommits_info_111_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_111_fpWen;
        io_diffCommits_info_111_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_111_vecWen;
        io_diffCommits_info_111_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_111_v0Wen;
        io_diffCommits_info_111_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_111_vlWen;
        io_diffCommits_info_112_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_112_ldest;
        io_diffCommits_info_112_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_112_pdest;
        io_diffCommits_info_112_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_112_rfWen;
        io_diffCommits_info_112_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_112_fpWen;
        io_diffCommits_info_112_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_112_vecWen;
        io_diffCommits_info_112_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_112_v0Wen;
        io_diffCommits_info_112_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_112_vlWen;
        io_diffCommits_info_113_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_113_ldest;
        io_diffCommits_info_113_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_113_pdest;
        io_diffCommits_info_113_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_113_rfWen;
        io_diffCommits_info_113_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_113_fpWen;
        io_diffCommits_info_113_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_113_vecWen;
        io_diffCommits_info_113_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_113_v0Wen;
        io_diffCommits_info_113_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_113_vlWen;
        io_diffCommits_info_114_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_114_ldest;
        io_diffCommits_info_114_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_114_pdest;
        io_diffCommits_info_114_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_114_rfWen;
        io_diffCommits_info_114_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_114_fpWen;
        io_diffCommits_info_114_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_114_vecWen;
        io_diffCommits_info_114_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_114_v0Wen;
        io_diffCommits_info_114_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_114_vlWen;
        io_diffCommits_info_115_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_115_ldest;
        io_diffCommits_info_115_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_115_pdest;
        io_diffCommits_info_115_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_115_rfWen;
        io_diffCommits_info_115_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_115_fpWen;
        io_diffCommits_info_115_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_115_vecWen;
        io_diffCommits_info_115_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_115_v0Wen;
        io_diffCommits_info_115_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_115_vlWen;
        io_diffCommits_info_116_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_116_ldest;
        io_diffCommits_info_116_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_116_pdest;
        io_diffCommits_info_116_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_116_rfWen;
        io_diffCommits_info_116_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_116_fpWen;
        io_diffCommits_info_116_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_116_vecWen;
        io_diffCommits_info_116_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_116_v0Wen;
        io_diffCommits_info_116_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_116_vlWen;
        io_diffCommits_info_117_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_117_ldest;
        io_diffCommits_info_117_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_117_pdest;
        io_diffCommits_info_117_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_117_rfWen;
        io_diffCommits_info_117_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_117_fpWen;
        io_diffCommits_info_117_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_117_vecWen;
        io_diffCommits_info_117_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_117_v0Wen;
        io_diffCommits_info_117_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_117_vlWen;
        io_diffCommits_info_118_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_118_ldest;
        io_diffCommits_info_118_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_118_pdest;
        io_diffCommits_info_118_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_118_rfWen;
        io_diffCommits_info_118_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_118_fpWen;
        io_diffCommits_info_118_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_118_vecWen;
        io_diffCommits_info_118_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_118_v0Wen;
        io_diffCommits_info_118_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_118_vlWen;
        io_diffCommits_info_119_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_119_ldest;
        io_diffCommits_info_119_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_119_pdest;
        io_diffCommits_info_119_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_119_rfWen;
        io_diffCommits_info_119_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_119_fpWen;
        io_diffCommits_info_119_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_119_vecWen;
        io_diffCommits_info_119_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_119_v0Wen;
        io_diffCommits_info_119_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_119_vlWen;
        io_diffCommits_info_120_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_120_ldest;
        io_diffCommits_info_120_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_120_pdest;
        io_diffCommits_info_120_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_120_rfWen;
        io_diffCommits_info_120_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_120_fpWen;
        io_diffCommits_info_120_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_120_vecWen;
        io_diffCommits_info_120_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_120_v0Wen;
        io_diffCommits_info_120_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_120_vlWen;
        io_diffCommits_info_121_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_121_ldest;
        io_diffCommits_info_121_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_121_pdest;
        io_diffCommits_info_121_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_121_rfWen;
        io_diffCommits_info_121_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_121_fpWen;
        io_diffCommits_info_121_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_121_vecWen;
        io_diffCommits_info_121_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_121_v0Wen;
        io_diffCommits_info_121_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_121_vlWen;
        io_diffCommits_info_122_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_122_ldest;
        io_diffCommits_info_122_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_122_pdest;
        io_diffCommits_info_122_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_122_rfWen;
        io_diffCommits_info_122_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_122_fpWen;
        io_diffCommits_info_122_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_122_vecWen;
        io_diffCommits_info_122_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_122_v0Wen;
        io_diffCommits_info_122_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_122_vlWen;
        io_diffCommits_info_123_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_123_ldest;
        io_diffCommits_info_123_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_123_pdest;
        io_diffCommits_info_123_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_123_rfWen;
        io_diffCommits_info_123_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_123_fpWen;
        io_diffCommits_info_123_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_123_vecWen;
        io_diffCommits_info_123_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_123_v0Wen;
        io_diffCommits_info_123_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_123_vlWen;
        io_diffCommits_info_124_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_124_ldest;
        io_diffCommits_info_124_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_124_pdest;
        io_diffCommits_info_124_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_124_rfWen;
        io_diffCommits_info_124_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_124_fpWen;
        io_diffCommits_info_124_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_124_vecWen;
        io_diffCommits_info_124_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_124_v0Wen;
        io_diffCommits_info_124_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_124_vlWen;
        io_diffCommits_info_125_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_125_ldest;
        io_diffCommits_info_125_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_125_pdest;
        io_diffCommits_info_125_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_125_rfWen;
        io_diffCommits_info_125_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_125_fpWen;
        io_diffCommits_info_125_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_125_vecWen;
        io_diffCommits_info_125_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_125_v0Wen;
        io_diffCommits_info_125_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_125_vlWen;
        io_diffCommits_info_126_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_126_ldest;
        io_diffCommits_info_126_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_126_pdest;
        io_diffCommits_info_126_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_126_rfWen;
        io_diffCommits_info_126_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_126_fpWen;
        io_diffCommits_info_126_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_126_vecWen;
        io_diffCommits_info_126_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_126_v0Wen;
        io_diffCommits_info_126_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_126_vlWen;
        io_diffCommits_info_127_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_127_ldest;
        io_diffCommits_info_127_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_127_pdest;
        io_diffCommits_info_127_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_127_rfWen;
        io_diffCommits_info_127_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_127_fpWen;
        io_diffCommits_info_127_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_127_vecWen;
        io_diffCommits_info_127_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_127_v0Wen;
        io_diffCommits_info_127_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_127_vlWen;
        io_diffCommits_info_128_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_128_ldest;
        io_diffCommits_info_128_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_128_pdest;
        io_diffCommits_info_128_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_128_rfWen;
        io_diffCommits_info_128_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_128_fpWen;
        io_diffCommits_info_128_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_128_vecWen;
        io_diffCommits_info_128_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_128_v0Wen;
        io_diffCommits_info_128_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_128_vlWen;
        io_diffCommits_info_129_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_129_ldest;
        io_diffCommits_info_129_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_129_pdest;
        io_diffCommits_info_129_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_129_rfWen;
        io_diffCommits_info_129_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_129_fpWen;
        io_diffCommits_info_129_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_129_vecWen;
        io_diffCommits_info_129_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_129_v0Wen;
        io_diffCommits_info_129_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_129_vlWen;
        io_diffCommits_info_130_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_130_ldest;
        io_diffCommits_info_130_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_130_pdest;
        io_diffCommits_info_130_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_130_rfWen;
        io_diffCommits_info_130_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_130_fpWen;
        io_diffCommits_info_130_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_130_vecWen;
        io_diffCommits_info_130_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_130_v0Wen;
        io_diffCommits_info_130_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_130_vlWen;
        io_diffCommits_info_131_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_131_ldest;
        io_diffCommits_info_131_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_131_pdest;
        io_diffCommits_info_131_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_131_rfWen;
        io_diffCommits_info_131_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_131_fpWen;
        io_diffCommits_info_131_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_131_vecWen;
        io_diffCommits_info_131_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_131_v0Wen;
        io_diffCommits_info_131_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_131_vlWen;
        io_diffCommits_info_132_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_132_ldest;
        io_diffCommits_info_132_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_132_pdest;
        io_diffCommits_info_132_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_132_rfWen;
        io_diffCommits_info_132_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_132_fpWen;
        io_diffCommits_info_132_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_132_vecWen;
        io_diffCommits_info_132_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_132_v0Wen;
        io_diffCommits_info_132_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_132_vlWen;
        io_diffCommits_info_133_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_133_ldest;
        io_diffCommits_info_133_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_133_pdest;
        io_diffCommits_info_133_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_133_rfWen;
        io_diffCommits_info_133_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_133_fpWen;
        io_diffCommits_info_133_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_133_vecWen;
        io_diffCommits_info_133_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_133_v0Wen;
        io_diffCommits_info_133_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_133_vlWen;
        io_diffCommits_info_134_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_134_ldest;
        io_diffCommits_info_134_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_134_pdest;
        io_diffCommits_info_134_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_134_rfWen;
        io_diffCommits_info_134_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_134_fpWen;
        io_diffCommits_info_134_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_134_vecWen;
        io_diffCommits_info_134_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_134_v0Wen;
        io_diffCommits_info_134_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_134_vlWen;
        io_diffCommits_info_135_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_135_ldest;
        io_diffCommits_info_135_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_135_pdest;
        io_diffCommits_info_135_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_135_rfWen;
        io_diffCommits_info_135_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_135_fpWen;
        io_diffCommits_info_135_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_135_vecWen;
        io_diffCommits_info_135_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_135_v0Wen;
        io_diffCommits_info_135_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_135_vlWen;
        io_diffCommits_info_136_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_136_ldest;
        io_diffCommits_info_136_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_136_pdest;
        io_diffCommits_info_136_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_136_rfWen;
        io_diffCommits_info_136_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_136_fpWen;
        io_diffCommits_info_136_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_136_vecWen;
        io_diffCommits_info_136_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_136_v0Wen;
        io_diffCommits_info_136_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_136_vlWen;
        io_diffCommits_info_137_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_137_ldest;
        io_diffCommits_info_137_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_137_pdest;
        io_diffCommits_info_137_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_137_rfWen;
        io_diffCommits_info_137_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_137_fpWen;
        io_diffCommits_info_137_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_137_vecWen;
        io_diffCommits_info_137_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_137_v0Wen;
        io_diffCommits_info_137_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_137_vlWen;
        io_diffCommits_info_138_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_138_ldest;
        io_diffCommits_info_138_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_138_pdest;
        io_diffCommits_info_138_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_138_rfWen;
        io_diffCommits_info_138_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_138_fpWen;
        io_diffCommits_info_138_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_138_vecWen;
        io_diffCommits_info_138_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_138_v0Wen;
        io_diffCommits_info_138_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_138_vlWen;
        io_diffCommits_info_139_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_139_ldest;
        io_diffCommits_info_139_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_139_pdest;
        io_diffCommits_info_139_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_139_rfWen;
        io_diffCommits_info_139_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_139_fpWen;
        io_diffCommits_info_139_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_139_vecWen;
        io_diffCommits_info_139_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_139_v0Wen;
        io_diffCommits_info_139_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_139_vlWen;
        io_diffCommits_info_140_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_140_ldest;
        io_diffCommits_info_140_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_140_pdest;
        io_diffCommits_info_140_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_140_rfWen;
        io_diffCommits_info_140_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_140_fpWen;
        io_diffCommits_info_140_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_140_vecWen;
        io_diffCommits_info_140_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_140_v0Wen;
        io_diffCommits_info_140_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_140_vlWen;
        io_diffCommits_info_141_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_141_ldest;
        io_diffCommits_info_141_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_141_pdest;
        io_diffCommits_info_141_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_141_rfWen;
        io_diffCommits_info_141_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_141_fpWen;
        io_diffCommits_info_141_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_141_vecWen;
        io_diffCommits_info_141_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_141_v0Wen;
        io_diffCommits_info_141_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_141_vlWen;
        io_diffCommits_info_142_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_142_ldest;
        io_diffCommits_info_142_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_142_pdest;
        io_diffCommits_info_142_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_142_rfWen;
        io_diffCommits_info_142_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_142_fpWen;
        io_diffCommits_info_142_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_142_vecWen;
        io_diffCommits_info_142_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_142_v0Wen;
        io_diffCommits_info_142_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_142_vlWen;
        io_diffCommits_info_143_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_143_ldest;
        io_diffCommits_info_143_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_143_pdest;
        io_diffCommits_info_143_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_143_rfWen;
        io_diffCommits_info_143_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_143_fpWen;
        io_diffCommits_info_143_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_143_vecWen;
        io_diffCommits_info_143_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_143_v0Wen;
        io_diffCommits_info_143_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_143_vlWen;
        io_diffCommits_info_144_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_144_ldest;
        io_diffCommits_info_144_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_144_pdest;
        io_diffCommits_info_144_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_144_rfWen;
        io_diffCommits_info_144_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_144_fpWen;
        io_diffCommits_info_144_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_144_vecWen;
        io_diffCommits_info_144_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_144_v0Wen;
        io_diffCommits_info_144_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_144_vlWen;
        io_diffCommits_info_145_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_145_ldest;
        io_diffCommits_info_145_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_145_pdest;
        io_diffCommits_info_145_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_145_rfWen;
        io_diffCommits_info_145_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_145_fpWen;
        io_diffCommits_info_145_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_145_vecWen;
        io_diffCommits_info_145_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_145_v0Wen;
        io_diffCommits_info_145_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_145_vlWen;
        io_diffCommits_info_146_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_146_ldest;
        io_diffCommits_info_146_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_146_pdest;
        io_diffCommits_info_146_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_146_rfWen;
        io_diffCommits_info_146_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_146_fpWen;
        io_diffCommits_info_146_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_146_vecWen;
        io_diffCommits_info_146_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_146_v0Wen;
        io_diffCommits_info_146_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_146_vlWen;
        io_diffCommits_info_147_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_147_ldest;
        io_diffCommits_info_147_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_147_pdest;
        io_diffCommits_info_147_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_147_rfWen;
        io_diffCommits_info_147_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_147_fpWen;
        io_diffCommits_info_147_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_147_vecWen;
        io_diffCommits_info_147_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_147_v0Wen;
        io_diffCommits_info_147_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_147_vlWen;
        io_diffCommits_info_148_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_148_ldest;
        io_diffCommits_info_148_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_148_pdest;
        io_diffCommits_info_148_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_148_rfWen;
        io_diffCommits_info_148_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_148_fpWen;
        io_diffCommits_info_148_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_148_vecWen;
        io_diffCommits_info_148_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_148_v0Wen;
        io_diffCommits_info_148_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_148_vlWen;
        io_diffCommits_info_149_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_149_ldest;
        io_diffCommits_info_149_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_149_pdest;
        io_diffCommits_info_149_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_149_rfWen;
        io_diffCommits_info_149_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_149_fpWen;
        io_diffCommits_info_149_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_149_vecWen;
        io_diffCommits_info_149_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_149_v0Wen;
        io_diffCommits_info_149_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_149_vlWen;
        io_diffCommits_info_150_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_150_ldest;
        io_diffCommits_info_150_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_150_pdest;
        io_diffCommits_info_150_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_150_rfWen;
        io_diffCommits_info_150_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_150_fpWen;
        io_diffCommits_info_150_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_150_vecWen;
        io_diffCommits_info_150_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_150_v0Wen;
        io_diffCommits_info_150_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_150_vlWen;
        io_diffCommits_info_151_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_151_ldest;
        io_diffCommits_info_151_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_151_pdest;
        io_diffCommits_info_151_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_151_rfWen;
        io_diffCommits_info_151_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_151_fpWen;
        io_diffCommits_info_151_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_151_vecWen;
        io_diffCommits_info_151_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_151_v0Wen;
        io_diffCommits_info_151_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_151_vlWen;
        io_diffCommits_info_152_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_152_ldest;
        io_diffCommits_info_152_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_152_pdest;
        io_diffCommits_info_152_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_152_rfWen;
        io_diffCommits_info_152_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_152_fpWen;
        io_diffCommits_info_152_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_152_vecWen;
        io_diffCommits_info_152_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_152_v0Wen;
        io_diffCommits_info_152_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_152_vlWen;
        io_diffCommits_info_153_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_153_ldest;
        io_diffCommits_info_153_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_153_pdest;
        io_diffCommits_info_153_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_153_rfWen;
        io_diffCommits_info_153_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_153_fpWen;
        io_diffCommits_info_153_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_153_vecWen;
        io_diffCommits_info_153_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_153_v0Wen;
        io_diffCommits_info_153_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_153_vlWen;
        io_diffCommits_info_154_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_154_ldest;
        io_diffCommits_info_154_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_154_pdest;
        io_diffCommits_info_154_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_154_rfWen;
        io_diffCommits_info_154_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_154_fpWen;
        io_diffCommits_info_154_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_154_vecWen;
        io_diffCommits_info_154_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_154_v0Wen;
        io_diffCommits_info_154_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_154_vlWen;
        io_diffCommits_info_155_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_155_ldest;
        io_diffCommits_info_155_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_155_pdest;
        io_diffCommits_info_155_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_155_rfWen;
        io_diffCommits_info_155_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_155_fpWen;
        io_diffCommits_info_155_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_155_vecWen;
        io_diffCommits_info_155_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_155_v0Wen;
        io_diffCommits_info_155_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_155_vlWen;
        io_diffCommits_info_156_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_156_ldest;
        io_diffCommits_info_156_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_156_pdest;
        io_diffCommits_info_156_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_156_rfWen;
        io_diffCommits_info_156_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_156_fpWen;
        io_diffCommits_info_156_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_156_vecWen;
        io_diffCommits_info_156_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_156_v0Wen;
        io_diffCommits_info_156_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_156_vlWen;
        io_diffCommits_info_157_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_157_ldest;
        io_diffCommits_info_157_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_157_pdest;
        io_diffCommits_info_157_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_157_rfWen;
        io_diffCommits_info_157_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_157_fpWen;
        io_diffCommits_info_157_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_157_vecWen;
        io_diffCommits_info_157_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_157_v0Wen;
        io_diffCommits_info_157_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_157_vlWen;
        io_diffCommits_info_158_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_158_ldest;
        io_diffCommits_info_158_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_158_pdest;
        io_diffCommits_info_158_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_158_rfWen;
        io_diffCommits_info_158_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_158_fpWen;
        io_diffCommits_info_158_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_158_vecWen;
        io_diffCommits_info_158_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_158_v0Wen;
        io_diffCommits_info_158_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_158_vlWen;
        io_diffCommits_info_159_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_159_ldest;
        io_diffCommits_info_159_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_159_pdest;
        io_diffCommits_info_159_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_159_rfWen;
        io_diffCommits_info_159_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_159_fpWen;
        io_diffCommits_info_159_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_159_vecWen;
        io_diffCommits_info_159_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_159_v0Wen;
        io_diffCommits_info_159_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_159_vlWen;
        io_diffCommits_info_160_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_160_ldest;
        io_diffCommits_info_160_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_160_pdest;
        io_diffCommits_info_160_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_160_rfWen;
        io_diffCommits_info_160_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_160_fpWen;
        io_diffCommits_info_160_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_160_vecWen;
        io_diffCommits_info_160_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_160_v0Wen;
        io_diffCommits_info_160_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_160_vlWen;
        io_diffCommits_info_161_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_161_ldest;
        io_diffCommits_info_161_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_161_pdest;
        io_diffCommits_info_161_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_161_rfWen;
        io_diffCommits_info_161_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_161_fpWen;
        io_diffCommits_info_161_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_161_vecWen;
        io_diffCommits_info_161_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_161_v0Wen;
        io_diffCommits_info_161_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_161_vlWen;
        io_diffCommits_info_162_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_162_ldest;
        io_diffCommits_info_162_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_162_pdest;
        io_diffCommits_info_162_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_162_rfWen;
        io_diffCommits_info_162_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_162_fpWen;
        io_diffCommits_info_162_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_162_vecWen;
        io_diffCommits_info_162_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_162_v0Wen;
        io_diffCommits_info_162_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_162_vlWen;
        io_diffCommits_info_163_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_163_ldest;
        io_diffCommits_info_163_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_163_pdest;
        io_diffCommits_info_163_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_163_rfWen;
        io_diffCommits_info_163_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_163_fpWen;
        io_diffCommits_info_163_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_163_vecWen;
        io_diffCommits_info_163_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_163_v0Wen;
        io_diffCommits_info_163_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_163_vlWen;
        io_diffCommits_info_164_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_164_ldest;
        io_diffCommits_info_164_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_164_pdest;
        io_diffCommits_info_164_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_164_rfWen;
        io_diffCommits_info_164_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_164_fpWen;
        io_diffCommits_info_164_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_164_vecWen;
        io_diffCommits_info_164_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_164_v0Wen;
        io_diffCommits_info_164_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_164_vlWen;
        io_diffCommits_info_165_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_165_ldest;
        io_diffCommits_info_165_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_165_pdest;
        io_diffCommits_info_165_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_165_rfWen;
        io_diffCommits_info_165_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_165_fpWen;
        io_diffCommits_info_165_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_165_vecWen;
        io_diffCommits_info_165_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_165_v0Wen;
        io_diffCommits_info_165_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_165_vlWen;
        io_diffCommits_info_166_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_166_ldest;
        io_diffCommits_info_166_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_166_pdest;
        io_diffCommits_info_166_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_166_rfWen;
        io_diffCommits_info_166_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_166_fpWen;
        io_diffCommits_info_166_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_166_vecWen;
        io_diffCommits_info_166_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_166_v0Wen;
        io_diffCommits_info_166_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_166_vlWen;
        io_diffCommits_info_167_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_167_ldest;
        io_diffCommits_info_167_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_167_pdest;
        io_diffCommits_info_167_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_167_rfWen;
        io_diffCommits_info_167_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_167_fpWen;
        io_diffCommits_info_167_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_167_vecWen;
        io_diffCommits_info_167_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_167_v0Wen;
        io_diffCommits_info_167_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_167_vlWen;
        io_diffCommits_info_168_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_168_ldest;
        io_diffCommits_info_168_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_168_pdest;
        io_diffCommits_info_168_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_168_rfWen;
        io_diffCommits_info_168_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_168_fpWen;
        io_diffCommits_info_168_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_168_vecWen;
        io_diffCommits_info_168_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_168_v0Wen;
        io_diffCommits_info_168_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_168_vlWen;
        io_diffCommits_info_169_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_169_ldest;
        io_diffCommits_info_169_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_169_pdest;
        io_diffCommits_info_169_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_169_rfWen;
        io_diffCommits_info_169_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_169_fpWen;
        io_diffCommits_info_169_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_169_vecWen;
        io_diffCommits_info_169_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_169_v0Wen;
        io_diffCommits_info_169_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_169_vlWen;
        io_diffCommits_info_170_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_170_ldest;
        io_diffCommits_info_170_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_170_pdest;
        io_diffCommits_info_170_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_170_rfWen;
        io_diffCommits_info_170_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_170_fpWen;
        io_diffCommits_info_170_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_170_vecWen;
        io_diffCommits_info_170_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_170_v0Wen;
        io_diffCommits_info_170_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_170_vlWen;
        io_diffCommits_info_171_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_171_ldest;
        io_diffCommits_info_171_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_171_pdest;
        io_diffCommits_info_171_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_171_rfWen;
        io_diffCommits_info_171_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_171_fpWen;
        io_diffCommits_info_171_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_171_vecWen;
        io_diffCommits_info_171_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_171_v0Wen;
        io_diffCommits_info_171_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_171_vlWen;
        io_diffCommits_info_172_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_172_ldest;
        io_diffCommits_info_172_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_172_pdest;
        io_diffCommits_info_172_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_172_rfWen;
        io_diffCommits_info_172_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_172_fpWen;
        io_diffCommits_info_172_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_172_vecWen;
        io_diffCommits_info_172_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_172_v0Wen;
        io_diffCommits_info_172_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_172_vlWen;
        io_diffCommits_info_173_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_173_ldest;
        io_diffCommits_info_173_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_173_pdest;
        io_diffCommits_info_173_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_173_rfWen;
        io_diffCommits_info_173_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_173_fpWen;
        io_diffCommits_info_173_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_173_vecWen;
        io_diffCommits_info_173_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_173_v0Wen;
        io_diffCommits_info_173_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_173_vlWen;
        io_diffCommits_info_174_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_174_ldest;
        io_diffCommits_info_174_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_174_pdest;
        io_diffCommits_info_174_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_174_rfWen;
        io_diffCommits_info_174_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_174_fpWen;
        io_diffCommits_info_174_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_174_vecWen;
        io_diffCommits_info_174_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_174_v0Wen;
        io_diffCommits_info_174_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_174_vlWen;
        io_diffCommits_info_175_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_175_ldest;
        io_diffCommits_info_175_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_175_pdest;
        io_diffCommits_info_175_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_175_rfWen;
        io_diffCommits_info_175_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_175_fpWen;
        io_diffCommits_info_175_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_175_vecWen;
        io_diffCommits_info_175_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_175_v0Wen;
        io_diffCommits_info_175_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_175_vlWen;
        io_diffCommits_info_176_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_176_ldest;
        io_diffCommits_info_176_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_176_pdest;
        io_diffCommits_info_176_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_176_rfWen;
        io_diffCommits_info_176_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_176_fpWen;
        io_diffCommits_info_176_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_176_vecWen;
        io_diffCommits_info_176_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_176_v0Wen;
        io_diffCommits_info_176_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_176_vlWen;
        io_diffCommits_info_177_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_177_ldest;
        io_diffCommits_info_177_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_177_pdest;
        io_diffCommits_info_177_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_177_rfWen;
        io_diffCommits_info_177_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_177_fpWen;
        io_diffCommits_info_177_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_177_vecWen;
        io_diffCommits_info_177_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_177_v0Wen;
        io_diffCommits_info_177_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_177_vlWen;
        io_diffCommits_info_178_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_178_ldest;
        io_diffCommits_info_178_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_178_pdest;
        io_diffCommits_info_178_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_178_rfWen;
        io_diffCommits_info_178_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_178_fpWen;
        io_diffCommits_info_178_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_178_vecWen;
        io_diffCommits_info_178_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_178_v0Wen;
        io_diffCommits_info_178_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_178_vlWen;
        io_diffCommits_info_179_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_179_ldest;
        io_diffCommits_info_179_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_179_pdest;
        io_diffCommits_info_179_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_179_rfWen;
        io_diffCommits_info_179_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_179_fpWen;
        io_diffCommits_info_179_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_179_vecWen;
        io_diffCommits_info_179_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_179_v0Wen;
        io_diffCommits_info_179_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_179_vlWen;
        io_diffCommits_info_180_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_180_ldest;
        io_diffCommits_info_180_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_180_pdest;
        io_diffCommits_info_180_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_180_rfWen;
        io_diffCommits_info_180_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_180_fpWen;
        io_diffCommits_info_180_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_180_vecWen;
        io_diffCommits_info_180_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_180_v0Wen;
        io_diffCommits_info_180_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_180_vlWen;
        io_diffCommits_info_181_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_181_ldest;
        io_diffCommits_info_181_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_181_pdest;
        io_diffCommits_info_181_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_181_rfWen;
        io_diffCommits_info_181_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_181_fpWen;
        io_diffCommits_info_181_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_181_vecWen;
        io_diffCommits_info_181_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_181_v0Wen;
        io_diffCommits_info_181_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_181_vlWen;
        io_diffCommits_info_182_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_182_ldest;
        io_diffCommits_info_182_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_182_pdest;
        io_diffCommits_info_182_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_182_rfWen;
        io_diffCommits_info_182_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_182_fpWen;
        io_diffCommits_info_182_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_182_vecWen;
        io_diffCommits_info_182_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_182_v0Wen;
        io_diffCommits_info_182_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_182_vlWen;
        io_diffCommits_info_183_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_183_ldest;
        io_diffCommits_info_183_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_183_pdest;
        io_diffCommits_info_183_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_183_rfWen;
        io_diffCommits_info_183_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_183_fpWen;
        io_diffCommits_info_183_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_183_vecWen;
        io_diffCommits_info_183_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_183_v0Wen;
        io_diffCommits_info_183_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_183_vlWen;
        io_diffCommits_info_184_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_184_ldest;
        io_diffCommits_info_184_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_184_pdest;
        io_diffCommits_info_184_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_184_rfWen;
        io_diffCommits_info_184_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_184_fpWen;
        io_diffCommits_info_184_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_184_vecWen;
        io_diffCommits_info_184_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_184_v0Wen;
        io_diffCommits_info_184_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_184_vlWen;
        io_diffCommits_info_185_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_185_ldest;
        io_diffCommits_info_185_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_185_pdest;
        io_diffCommits_info_185_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_185_rfWen;
        io_diffCommits_info_185_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_185_fpWen;
        io_diffCommits_info_185_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_185_vecWen;
        io_diffCommits_info_185_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_185_v0Wen;
        io_diffCommits_info_185_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_185_vlWen;
        io_diffCommits_info_186_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_186_ldest;
        io_diffCommits_info_186_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_186_pdest;
        io_diffCommits_info_186_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_186_rfWen;
        io_diffCommits_info_186_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_186_fpWen;
        io_diffCommits_info_186_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_186_vecWen;
        io_diffCommits_info_186_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_186_v0Wen;
        io_diffCommits_info_186_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_186_vlWen;
        io_diffCommits_info_187_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_187_ldest;
        io_diffCommits_info_187_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_187_pdest;
        io_diffCommits_info_187_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_187_rfWen;
        io_diffCommits_info_187_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_187_fpWen;
        io_diffCommits_info_187_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_187_vecWen;
        io_diffCommits_info_187_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_187_v0Wen;
        io_diffCommits_info_187_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_187_vlWen;
        io_diffCommits_info_188_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_188_ldest;
        io_diffCommits_info_188_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_188_pdest;
        io_diffCommits_info_188_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_188_rfWen;
        io_diffCommits_info_188_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_188_fpWen;
        io_diffCommits_info_188_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_188_vecWen;
        io_diffCommits_info_188_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_188_v0Wen;
        io_diffCommits_info_188_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_188_vlWen;
        io_diffCommits_info_189_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_189_ldest;
        io_diffCommits_info_189_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_189_pdest;
        io_diffCommits_info_189_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_189_rfWen;
        io_diffCommits_info_189_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_189_fpWen;
        io_diffCommits_info_189_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_189_vecWen;
        io_diffCommits_info_189_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_189_v0Wen;
        io_diffCommits_info_189_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_189_vlWen;
        io_diffCommits_info_190_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_190_ldest;
        io_diffCommits_info_190_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_190_pdest;
        io_diffCommits_info_190_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_190_rfWen;
        io_diffCommits_info_190_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_190_fpWen;
        io_diffCommits_info_190_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_190_vecWen;
        io_diffCommits_info_190_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_190_v0Wen;
        io_diffCommits_info_190_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_190_vlWen;
        io_diffCommits_info_191_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_191_ldest;
        io_diffCommits_info_191_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_191_pdest;
        io_diffCommits_info_191_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_191_rfWen;
        io_diffCommits_info_191_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_191_fpWen;
        io_diffCommits_info_191_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_191_vecWen;
        io_diffCommits_info_191_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_191_v0Wen;
        io_diffCommits_info_191_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_191_vlWen;
        io_diffCommits_info_192_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_192_ldest;
        io_diffCommits_info_192_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_192_pdest;
        io_diffCommits_info_192_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_192_rfWen;
        io_diffCommits_info_192_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_192_fpWen;
        io_diffCommits_info_192_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_192_vecWen;
        io_diffCommits_info_192_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_192_v0Wen;
        io_diffCommits_info_192_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_192_vlWen;
        io_diffCommits_info_193_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_193_ldest;
        io_diffCommits_info_193_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_193_pdest;
        io_diffCommits_info_193_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_193_rfWen;
        io_diffCommits_info_193_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_193_fpWen;
        io_diffCommits_info_193_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_193_vecWen;
        io_diffCommits_info_193_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_193_v0Wen;
        io_diffCommits_info_193_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_193_vlWen;
        io_diffCommits_info_194_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_194_ldest;
        io_diffCommits_info_194_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_194_pdest;
        io_diffCommits_info_194_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_194_rfWen;
        io_diffCommits_info_194_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_194_fpWen;
        io_diffCommits_info_194_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_194_vecWen;
        io_diffCommits_info_194_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_194_v0Wen;
        io_diffCommits_info_194_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_194_vlWen;
        io_diffCommits_info_195_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_195_ldest;
        io_diffCommits_info_195_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_195_pdest;
        io_diffCommits_info_195_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_195_rfWen;
        io_diffCommits_info_195_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_195_fpWen;
        io_diffCommits_info_195_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_195_vecWen;
        io_diffCommits_info_195_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_195_v0Wen;
        io_diffCommits_info_195_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_195_vlWen;
        io_diffCommits_info_196_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_196_ldest;
        io_diffCommits_info_196_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_196_pdest;
        io_diffCommits_info_196_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_196_rfWen;
        io_diffCommits_info_196_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_196_fpWen;
        io_diffCommits_info_196_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_196_vecWen;
        io_diffCommits_info_196_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_196_v0Wen;
        io_diffCommits_info_196_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_196_vlWen;
        io_diffCommits_info_197_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_197_ldest;
        io_diffCommits_info_197_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_197_pdest;
        io_diffCommits_info_197_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_197_rfWen;
        io_diffCommits_info_197_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_197_fpWen;
        io_diffCommits_info_197_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_197_vecWen;
        io_diffCommits_info_197_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_197_v0Wen;
        io_diffCommits_info_197_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_197_vlWen;
        io_diffCommits_info_198_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_198_ldest;
        io_diffCommits_info_198_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_198_pdest;
        io_diffCommits_info_198_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_198_rfWen;
        io_diffCommits_info_198_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_198_fpWen;
        io_diffCommits_info_198_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_198_vecWen;
        io_diffCommits_info_198_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_198_v0Wen;
        io_diffCommits_info_198_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_198_vlWen;
        io_diffCommits_info_199_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_199_ldest;
        io_diffCommits_info_199_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_199_pdest;
        io_diffCommits_info_199_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_199_rfWen;
        io_diffCommits_info_199_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_199_fpWen;
        io_diffCommits_info_199_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_199_vecWen;
        io_diffCommits_info_199_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_199_v0Wen;
        io_diffCommits_info_199_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_199_vlWen;
        io_diffCommits_info_200_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_200_ldest;
        io_diffCommits_info_200_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_200_pdest;
        io_diffCommits_info_200_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_200_rfWen;
        io_diffCommits_info_200_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_200_fpWen;
        io_diffCommits_info_200_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_200_vecWen;
        io_diffCommits_info_200_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_200_v0Wen;
        io_diffCommits_info_200_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_200_vlWen;
        io_diffCommits_info_201_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_201_ldest;
        io_diffCommits_info_201_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_201_pdest;
        io_diffCommits_info_201_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_201_rfWen;
        io_diffCommits_info_201_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_201_fpWen;
        io_diffCommits_info_201_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_201_vecWen;
        io_diffCommits_info_201_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_201_v0Wen;
        io_diffCommits_info_201_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_201_vlWen;
        io_diffCommits_info_202_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_202_ldest;
        io_diffCommits_info_202_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_202_pdest;
        io_diffCommits_info_202_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_202_rfWen;
        io_diffCommits_info_202_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_202_fpWen;
        io_diffCommits_info_202_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_202_vecWen;
        io_diffCommits_info_202_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_202_v0Wen;
        io_diffCommits_info_202_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_202_vlWen;
        io_diffCommits_info_203_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_203_ldest;
        io_diffCommits_info_203_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_203_pdest;
        io_diffCommits_info_203_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_203_rfWen;
        io_diffCommits_info_203_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_203_fpWen;
        io_diffCommits_info_203_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_203_vecWen;
        io_diffCommits_info_203_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_203_v0Wen;
        io_diffCommits_info_203_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_203_vlWen;
        io_diffCommits_info_204_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_204_ldest;
        io_diffCommits_info_204_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_204_pdest;
        io_diffCommits_info_204_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_204_rfWen;
        io_diffCommits_info_204_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_204_fpWen;
        io_diffCommits_info_204_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_204_vecWen;
        io_diffCommits_info_204_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_204_v0Wen;
        io_diffCommits_info_204_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_204_vlWen;
        io_diffCommits_info_205_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_205_ldest;
        io_diffCommits_info_205_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_205_pdest;
        io_diffCommits_info_205_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_205_rfWen;
        io_diffCommits_info_205_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_205_fpWen;
        io_diffCommits_info_205_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_205_vecWen;
        io_diffCommits_info_205_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_205_v0Wen;
        io_diffCommits_info_205_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_205_vlWen;
        io_diffCommits_info_206_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_206_ldest;
        io_diffCommits_info_206_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_206_pdest;
        io_diffCommits_info_206_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_206_rfWen;
        io_diffCommits_info_206_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_206_fpWen;
        io_diffCommits_info_206_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_206_vecWen;
        io_diffCommits_info_206_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_206_v0Wen;
        io_diffCommits_info_206_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_206_vlWen;
        io_diffCommits_info_207_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_207_ldest;
        io_diffCommits_info_207_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_207_pdest;
        io_diffCommits_info_207_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_207_rfWen;
        io_diffCommits_info_207_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_207_fpWen;
        io_diffCommits_info_207_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_207_vecWen;
        io_diffCommits_info_207_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_207_v0Wen;
        io_diffCommits_info_207_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_207_vlWen;
        io_diffCommits_info_208_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_208_ldest;
        io_diffCommits_info_208_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_208_pdest;
        io_diffCommits_info_208_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_208_rfWen;
        io_diffCommits_info_208_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_208_fpWen;
        io_diffCommits_info_208_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_208_vecWen;
        io_diffCommits_info_208_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_208_v0Wen;
        io_diffCommits_info_208_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_208_vlWen;
        io_diffCommits_info_209_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_209_ldest;
        io_diffCommits_info_209_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_209_pdest;
        io_diffCommits_info_209_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_209_rfWen;
        io_diffCommits_info_209_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_209_fpWen;
        io_diffCommits_info_209_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_209_vecWen;
        io_diffCommits_info_209_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_209_v0Wen;
        io_diffCommits_info_209_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_209_vlWen;
        io_diffCommits_info_210_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_210_ldest;
        io_diffCommits_info_210_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_210_pdest;
        io_diffCommits_info_210_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_210_rfWen;
        io_diffCommits_info_210_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_210_fpWen;
        io_diffCommits_info_210_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_210_vecWen;
        io_diffCommits_info_210_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_210_v0Wen;
        io_diffCommits_info_210_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_210_vlWen;
        io_diffCommits_info_211_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_211_ldest;
        io_diffCommits_info_211_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_211_pdest;
        io_diffCommits_info_211_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_211_rfWen;
        io_diffCommits_info_211_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_211_fpWen;
        io_diffCommits_info_211_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_211_vecWen;
        io_diffCommits_info_211_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_211_v0Wen;
        io_diffCommits_info_211_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_211_vlWen;
        io_diffCommits_info_212_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_212_ldest;
        io_diffCommits_info_212_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_212_pdest;
        io_diffCommits_info_212_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_212_rfWen;
        io_diffCommits_info_212_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_212_fpWen;
        io_diffCommits_info_212_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_212_vecWen;
        io_diffCommits_info_212_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_212_v0Wen;
        io_diffCommits_info_212_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_212_vlWen;
        io_diffCommits_info_213_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_213_ldest;
        io_diffCommits_info_213_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_213_pdest;
        io_diffCommits_info_213_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_213_rfWen;
        io_diffCommits_info_213_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_213_fpWen;
        io_diffCommits_info_213_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_213_vecWen;
        io_diffCommits_info_213_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_213_v0Wen;
        io_diffCommits_info_213_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_213_vlWen;
        io_diffCommits_info_214_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_214_ldest;
        io_diffCommits_info_214_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_214_pdest;
        io_diffCommits_info_214_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_214_rfWen;
        io_diffCommits_info_214_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_214_fpWen;
        io_diffCommits_info_214_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_214_vecWen;
        io_diffCommits_info_214_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_214_v0Wen;
        io_diffCommits_info_214_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_214_vlWen;
        io_diffCommits_info_215_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_215_ldest;
        io_diffCommits_info_215_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_215_pdest;
        io_diffCommits_info_215_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_215_rfWen;
        io_diffCommits_info_215_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_215_fpWen;
        io_diffCommits_info_215_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_215_vecWen;
        io_diffCommits_info_215_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_215_v0Wen;
        io_diffCommits_info_215_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_215_vlWen;
        io_diffCommits_info_216_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_216_ldest;
        io_diffCommits_info_216_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_216_pdest;
        io_diffCommits_info_216_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_216_rfWen;
        io_diffCommits_info_216_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_216_fpWen;
        io_diffCommits_info_216_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_216_vecWen;
        io_diffCommits_info_216_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_216_v0Wen;
        io_diffCommits_info_216_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_216_vlWen;
        io_diffCommits_info_217_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_217_ldest;
        io_diffCommits_info_217_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_217_pdest;
        io_diffCommits_info_217_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_217_rfWen;
        io_diffCommits_info_217_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_217_fpWen;
        io_diffCommits_info_217_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_217_vecWen;
        io_diffCommits_info_217_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_217_v0Wen;
        io_diffCommits_info_217_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_217_vlWen;
        io_diffCommits_info_218_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_218_ldest;
        io_diffCommits_info_218_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_218_pdest;
        io_diffCommits_info_218_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_218_rfWen;
        io_diffCommits_info_218_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_218_fpWen;
        io_diffCommits_info_218_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_218_vecWen;
        io_diffCommits_info_218_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_218_v0Wen;
        io_diffCommits_info_218_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_218_vlWen;
        io_diffCommits_info_219_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_219_ldest;
        io_diffCommits_info_219_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_219_pdest;
        io_diffCommits_info_219_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_219_rfWen;
        io_diffCommits_info_219_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_219_fpWen;
        io_diffCommits_info_219_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_219_vecWen;
        io_diffCommits_info_219_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_219_v0Wen;
        io_diffCommits_info_219_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_219_vlWen;
        io_diffCommits_info_220_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_220_ldest;
        io_diffCommits_info_220_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_220_pdest;
        io_diffCommits_info_220_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_220_rfWen;
        io_diffCommits_info_220_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_220_fpWen;
        io_diffCommits_info_220_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_220_vecWen;
        io_diffCommits_info_220_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_220_v0Wen;
        io_diffCommits_info_220_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_220_vlWen;
        io_diffCommits_info_221_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_221_ldest;
        io_diffCommits_info_221_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_221_pdest;
        io_diffCommits_info_221_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_221_rfWen;
        io_diffCommits_info_221_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_221_fpWen;
        io_diffCommits_info_221_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_221_vecWen;
        io_diffCommits_info_221_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_221_v0Wen;
        io_diffCommits_info_221_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_221_vlWen;
        io_diffCommits_info_222_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_222_ldest;
        io_diffCommits_info_222_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_222_pdest;
        io_diffCommits_info_222_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_222_rfWen;
        io_diffCommits_info_222_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_222_fpWen;
        io_diffCommits_info_222_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_222_vecWen;
        io_diffCommits_info_222_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_222_v0Wen;
        io_diffCommits_info_222_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_222_vlWen;
        io_diffCommits_info_223_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_223_ldest;
        io_diffCommits_info_223_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_223_pdest;
        io_diffCommits_info_223_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_223_rfWen;
        io_diffCommits_info_223_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_223_fpWen;
        io_diffCommits_info_223_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_223_vecWen;
        io_diffCommits_info_223_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_223_v0Wen;
        io_diffCommits_info_223_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_223_vlWen;
        io_diffCommits_info_224_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_224_ldest;
        io_diffCommits_info_224_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_224_pdest;
        io_diffCommits_info_224_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_224_rfWen;
        io_diffCommits_info_224_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_224_fpWen;
        io_diffCommits_info_224_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_224_vecWen;
        io_diffCommits_info_224_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_224_v0Wen;
        io_diffCommits_info_224_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_224_vlWen;
        io_diffCommits_info_225_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_225_ldest;
        io_diffCommits_info_225_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_225_pdest;
        io_diffCommits_info_225_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_225_rfWen;
        io_diffCommits_info_225_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_225_fpWen;
        io_diffCommits_info_225_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_225_vecWen;
        io_diffCommits_info_225_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_225_v0Wen;
        io_diffCommits_info_225_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_225_vlWen;
        io_diffCommits_info_226_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_226_ldest;
        io_diffCommits_info_226_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_226_pdest;
        io_diffCommits_info_226_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_226_rfWen;
        io_diffCommits_info_226_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_226_fpWen;
        io_diffCommits_info_226_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_226_vecWen;
        io_diffCommits_info_226_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_226_v0Wen;
        io_diffCommits_info_226_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_226_vlWen;
        io_diffCommits_info_227_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_227_ldest;
        io_diffCommits_info_227_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_227_pdest;
        io_diffCommits_info_227_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_227_rfWen;
        io_diffCommits_info_227_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_227_fpWen;
        io_diffCommits_info_227_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_227_vecWen;
        io_diffCommits_info_227_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_227_v0Wen;
        io_diffCommits_info_227_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_227_vlWen;
        io_diffCommits_info_228_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_228_ldest;
        io_diffCommits_info_228_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_228_pdest;
        io_diffCommits_info_228_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_228_rfWen;
        io_diffCommits_info_228_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_228_fpWen;
        io_diffCommits_info_228_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_228_vecWen;
        io_diffCommits_info_228_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_228_v0Wen;
        io_diffCommits_info_228_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_228_vlWen;
        io_diffCommits_info_229_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_229_ldest;
        io_diffCommits_info_229_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_229_pdest;
        io_diffCommits_info_229_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_229_rfWen;
        io_diffCommits_info_229_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_229_fpWen;
        io_diffCommits_info_229_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_229_vecWen;
        io_diffCommits_info_229_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_229_v0Wen;
        io_diffCommits_info_229_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_229_vlWen;
        io_diffCommits_info_230_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_230_ldest;
        io_diffCommits_info_230_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_230_pdest;
        io_diffCommits_info_230_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_230_rfWen;
        io_diffCommits_info_230_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_230_fpWen;
        io_diffCommits_info_230_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_230_vecWen;
        io_diffCommits_info_230_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_230_v0Wen;
        io_diffCommits_info_230_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_230_vlWen;
        io_diffCommits_info_231_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_231_ldest;
        io_diffCommits_info_231_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_231_pdest;
        io_diffCommits_info_231_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_231_rfWen;
        io_diffCommits_info_231_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_231_fpWen;
        io_diffCommits_info_231_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_231_vecWen;
        io_diffCommits_info_231_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_231_v0Wen;
        io_diffCommits_info_231_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_231_vlWen;
        io_diffCommits_info_232_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_232_ldest;
        io_diffCommits_info_232_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_232_pdest;
        io_diffCommits_info_232_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_232_rfWen;
        io_diffCommits_info_232_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_232_fpWen;
        io_diffCommits_info_232_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_232_vecWen;
        io_diffCommits_info_232_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_232_v0Wen;
        io_diffCommits_info_232_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_232_vlWen;
        io_diffCommits_info_233_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_233_ldest;
        io_diffCommits_info_233_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_233_pdest;
        io_diffCommits_info_233_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_233_rfWen;
        io_diffCommits_info_233_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_233_fpWen;
        io_diffCommits_info_233_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_233_vecWen;
        io_diffCommits_info_233_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_233_v0Wen;
        io_diffCommits_info_233_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_233_vlWen;
        io_diffCommits_info_234_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_234_ldest;
        io_diffCommits_info_234_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_234_pdest;
        io_diffCommits_info_234_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_234_rfWen;
        io_diffCommits_info_234_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_234_fpWen;
        io_diffCommits_info_234_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_234_vecWen;
        io_diffCommits_info_234_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_234_v0Wen;
        io_diffCommits_info_234_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_234_vlWen;
        io_diffCommits_info_235_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_235_ldest;
        io_diffCommits_info_235_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_235_pdest;
        io_diffCommits_info_235_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_235_rfWen;
        io_diffCommits_info_235_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_235_fpWen;
        io_diffCommits_info_235_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_235_vecWen;
        io_diffCommits_info_235_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_235_v0Wen;
        io_diffCommits_info_235_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_235_vlWen;
        io_diffCommits_info_236_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_236_ldest;
        io_diffCommits_info_236_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_236_pdest;
        io_diffCommits_info_236_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_236_rfWen;
        io_diffCommits_info_236_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_236_fpWen;
        io_diffCommits_info_236_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_236_vecWen;
        io_diffCommits_info_236_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_236_v0Wen;
        io_diffCommits_info_236_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_236_vlWen;
        io_diffCommits_info_237_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_237_ldest;
        io_diffCommits_info_237_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_237_pdest;
        io_diffCommits_info_237_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_237_rfWen;
        io_diffCommits_info_237_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_237_fpWen;
        io_diffCommits_info_237_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_237_vecWen;
        io_diffCommits_info_237_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_237_v0Wen;
        io_diffCommits_info_237_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_237_vlWen;
        io_diffCommits_info_238_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_238_ldest;
        io_diffCommits_info_238_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_238_pdest;
        io_diffCommits_info_238_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_238_rfWen;
        io_diffCommits_info_238_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_238_fpWen;
        io_diffCommits_info_238_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_238_vecWen;
        io_diffCommits_info_238_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_238_v0Wen;
        io_diffCommits_info_238_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_238_vlWen;
        io_diffCommits_info_239_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_239_ldest;
        io_diffCommits_info_239_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_239_pdest;
        io_diffCommits_info_239_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_239_rfWen;
        io_diffCommits_info_239_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_239_fpWen;
        io_diffCommits_info_239_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_239_vecWen;
        io_diffCommits_info_239_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_239_v0Wen;
        io_diffCommits_info_239_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_239_vlWen;
        io_diffCommits_info_240_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_240_ldest;
        io_diffCommits_info_240_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_240_pdest;
        io_diffCommits_info_240_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_240_rfWen;
        io_diffCommits_info_240_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_240_fpWen;
        io_diffCommits_info_240_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_240_vecWen;
        io_diffCommits_info_240_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_240_v0Wen;
        io_diffCommits_info_240_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_240_vlWen;
        io_diffCommits_info_241_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_241_ldest;
        io_diffCommits_info_241_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_241_pdest;
        io_diffCommits_info_241_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_241_rfWen;
        io_diffCommits_info_241_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_241_fpWen;
        io_diffCommits_info_241_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_241_vecWen;
        io_diffCommits_info_241_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_241_v0Wen;
        io_diffCommits_info_241_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_241_vlWen;
        io_diffCommits_info_242_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_242_ldest;
        io_diffCommits_info_242_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_242_pdest;
        io_diffCommits_info_242_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_242_rfWen;
        io_diffCommits_info_242_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_242_fpWen;
        io_diffCommits_info_242_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_242_vecWen;
        io_diffCommits_info_242_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_242_v0Wen;
        io_diffCommits_info_242_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_242_vlWen;
        io_diffCommits_info_243_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_243_ldest;
        io_diffCommits_info_243_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_243_pdest;
        io_diffCommits_info_243_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_243_rfWen;
        io_diffCommits_info_243_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_243_fpWen;
        io_diffCommits_info_243_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_243_vecWen;
        io_diffCommits_info_243_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_243_v0Wen;
        io_diffCommits_info_243_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_243_vlWen;
        io_diffCommits_info_244_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_244_ldest;
        io_diffCommits_info_244_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_244_pdest;
        io_diffCommits_info_244_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_244_rfWen;
        io_diffCommits_info_244_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_244_fpWen;
        io_diffCommits_info_244_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_244_vecWen;
        io_diffCommits_info_244_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_244_v0Wen;
        io_diffCommits_info_244_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_244_vlWen;
        io_diffCommits_info_245_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_245_ldest;
        io_diffCommits_info_245_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_245_pdest;
        io_diffCommits_info_245_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_245_rfWen;
        io_diffCommits_info_245_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_245_fpWen;
        io_diffCommits_info_245_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_245_vecWen;
        io_diffCommits_info_245_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_245_v0Wen;
        io_diffCommits_info_245_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_245_vlWen;
        io_diffCommits_info_246_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_246_ldest;
        io_diffCommits_info_246_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_246_pdest;
        io_diffCommits_info_246_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_246_rfWen;
        io_diffCommits_info_246_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_246_fpWen;
        io_diffCommits_info_246_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_246_vecWen;
        io_diffCommits_info_246_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_246_v0Wen;
        io_diffCommits_info_246_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_246_vlWen;
        io_diffCommits_info_247_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_247_ldest;
        io_diffCommits_info_247_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_247_pdest;
        io_diffCommits_info_247_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_247_rfWen;
        io_diffCommits_info_247_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_247_fpWen;
        io_diffCommits_info_247_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_247_vecWen;
        io_diffCommits_info_247_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_247_v0Wen;
        io_diffCommits_info_247_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_247_vlWen;
        io_diffCommits_info_248_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_248_ldest;
        io_diffCommits_info_248_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_248_pdest;
        io_diffCommits_info_248_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_248_rfWen;
        io_diffCommits_info_248_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_248_fpWen;
        io_diffCommits_info_248_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_248_vecWen;
        io_diffCommits_info_248_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_248_v0Wen;
        io_diffCommits_info_248_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_248_vlWen;
        io_diffCommits_info_249_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_249_ldest;
        io_diffCommits_info_249_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_249_pdest;
        io_diffCommits_info_249_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_249_rfWen;
        io_diffCommits_info_249_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_249_fpWen;
        io_diffCommits_info_249_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_249_vecWen;
        io_diffCommits_info_249_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_249_v0Wen;
        io_diffCommits_info_249_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_249_vlWen;
        io_diffCommits_info_250_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_250_ldest;
        io_diffCommits_info_250_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_250_pdest;
        io_diffCommits_info_250_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_250_rfWen;
        io_diffCommits_info_250_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_250_fpWen;
        io_diffCommits_info_250_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_250_vecWen;
        io_diffCommits_info_250_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_250_v0Wen;
        io_diffCommits_info_250_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_250_vlWen;
        io_diffCommits_info_251_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_251_ldest;
        io_diffCommits_info_251_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_251_pdest;
        io_diffCommits_info_251_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_251_rfWen;
        io_diffCommits_info_251_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_251_fpWen;
        io_diffCommits_info_251_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_251_vecWen;
        io_diffCommits_info_251_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_251_v0Wen;
        io_diffCommits_info_251_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_251_vlWen;
        io_diffCommits_info_252_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_252_ldest;
        io_diffCommits_info_252_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_252_pdest;
        io_diffCommits_info_252_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_252_rfWen;
        io_diffCommits_info_252_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_252_fpWen;
        io_diffCommits_info_252_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_252_vecWen;
        io_diffCommits_info_252_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_252_v0Wen;
        io_diffCommits_info_252_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_252_vlWen;
        io_diffCommits_info_253_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_253_ldest;
        io_diffCommits_info_253_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_253_pdest;
        io_diffCommits_info_253_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_253_rfWen;
        io_diffCommits_info_253_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_253_fpWen;
        io_diffCommits_info_253_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_253_vecWen;
        io_diffCommits_info_253_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_253_v0Wen;
        io_diffCommits_info_253_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_253_vlWen;
        io_diffCommits_info_254_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_254_ldest;
        io_diffCommits_info_254_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_254_pdest;
        io_diffCommits_info_254_rfWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_254_rfWen;
        io_diffCommits_info_254_fpWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_254_fpWen;
        io_diffCommits_info_254_vecWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_254_vecWen;
        io_diffCommits_info_254_v0Wen = this.vif.mon_mp.mon_cb.io_diffCommits_info_254_v0Wen;
        io_diffCommits_info_254_vlWen = this.vif.mon_mp.mon_cb.io_diffCommits_info_254_vlWen;
        io_diffCommits_info_255_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_255_ldest;
        io_diffCommits_info_255_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_255_pdest;
        io_diffCommits_info_256_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_256_ldest;
        io_diffCommits_info_256_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_256_pdest;
        io_diffCommits_info_257_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_257_ldest;
        io_diffCommits_info_257_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_257_pdest;
        io_diffCommits_info_258_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_258_ldest;
        io_diffCommits_info_258_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_258_pdest;
        io_diffCommits_info_259_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_259_ldest;
        io_diffCommits_info_259_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_259_pdest;
        io_diffCommits_info_260_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_260_ldest;
        io_diffCommits_info_260_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_260_pdest;
        io_diffCommits_info_261_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_261_ldest;
        io_diffCommits_info_261_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_261_pdest;
        io_diffCommits_info_262_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_262_ldest;
        io_diffCommits_info_262_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_262_pdest;
        io_diffCommits_info_263_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_263_ldest;
        io_diffCommits_info_263_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_263_pdest;
        io_diffCommits_info_264_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_264_ldest;
        io_diffCommits_info_264_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_264_pdest;
        io_diffCommits_info_265_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_265_ldest;
        io_diffCommits_info_265_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_265_pdest;
        io_diffCommits_info_266_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_266_ldest;
        io_diffCommits_info_266_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_266_pdest;
        io_diffCommits_info_267_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_267_ldest;
        io_diffCommits_info_267_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_267_pdest;
        io_diffCommits_info_268_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_268_ldest;
        io_diffCommits_info_268_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_268_pdest;
        io_diffCommits_info_269_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_269_ldest;
        io_diffCommits_info_269_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_269_pdest;
        io_diffCommits_info_270_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_270_ldest;
        io_diffCommits_info_270_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_270_pdest;
        io_diffCommits_info_271_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_271_ldest;
        io_diffCommits_info_271_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_271_pdest;
        io_diffCommits_info_272_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_272_ldest;
        io_diffCommits_info_272_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_272_pdest;
        io_diffCommits_info_273_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_273_ldest;
        io_diffCommits_info_273_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_273_pdest;
        io_diffCommits_info_274_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_274_ldest;
        io_diffCommits_info_274_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_274_pdest;
        io_diffCommits_info_275_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_275_ldest;
        io_diffCommits_info_275_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_275_pdest;
        io_diffCommits_info_276_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_276_ldest;
        io_diffCommits_info_276_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_276_pdest;
        io_diffCommits_info_277_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_277_ldest;
        io_diffCommits_info_277_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_277_pdest;
        io_diffCommits_info_278_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_278_ldest;
        io_diffCommits_info_278_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_278_pdest;
        io_diffCommits_info_279_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_279_ldest;
        io_diffCommits_info_279_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_279_pdest;
        io_diffCommits_info_280_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_280_ldest;
        io_diffCommits_info_280_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_280_pdest;
        io_diffCommits_info_281_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_281_ldest;
        io_diffCommits_info_281_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_281_pdest;
        io_diffCommits_info_282_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_282_ldest;
        io_diffCommits_info_282_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_282_pdest;
        io_diffCommits_info_283_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_283_ldest;
        io_diffCommits_info_283_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_283_pdest;
        io_diffCommits_info_284_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_284_ldest;
        io_diffCommits_info_284_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_284_pdest;
        io_diffCommits_info_285_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_285_ldest;
        io_diffCommits_info_285_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_285_pdest;
        io_diffCommits_info_286_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_286_ldest;
        io_diffCommits_info_286_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_286_pdest;
        io_diffCommits_info_287_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_287_ldest;
        io_diffCommits_info_287_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_287_pdest;
        io_diffCommits_info_288_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_288_ldest;
        io_diffCommits_info_288_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_288_pdest;
        io_diffCommits_info_289_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_289_ldest;
        io_diffCommits_info_289_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_289_pdest;
        io_diffCommits_info_290_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_290_ldest;
        io_diffCommits_info_290_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_290_pdest;
        io_diffCommits_info_291_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_291_ldest;
        io_diffCommits_info_291_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_291_pdest;
        io_diffCommits_info_292_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_292_ldest;
        io_diffCommits_info_292_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_292_pdest;
        io_diffCommits_info_293_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_293_ldest;
        io_diffCommits_info_293_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_293_pdest;
        io_diffCommits_info_294_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_294_ldest;
        io_diffCommits_info_294_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_294_pdest;
        io_diffCommits_info_295_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_295_ldest;
        io_diffCommits_info_295_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_295_pdest;
        io_diffCommits_info_296_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_296_ldest;
        io_diffCommits_info_296_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_296_pdest;
        io_diffCommits_info_297_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_297_ldest;
        io_diffCommits_info_297_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_297_pdest;
        io_diffCommits_info_298_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_298_ldest;
        io_diffCommits_info_298_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_298_pdest;
        io_diffCommits_info_299_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_299_ldest;
        io_diffCommits_info_299_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_299_pdest;
        io_diffCommits_info_300_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_300_ldest;
        io_diffCommits_info_300_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_300_pdest;
        io_diffCommits_info_301_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_301_ldest;
        io_diffCommits_info_301_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_301_pdest;
        io_diffCommits_info_302_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_302_ldest;
        io_diffCommits_info_302_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_302_pdest;
        io_diffCommits_info_303_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_303_ldest;
        io_diffCommits_info_303_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_303_pdest;
        io_diffCommits_info_304_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_304_ldest;
        io_diffCommits_info_304_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_304_pdest;
        io_diffCommits_info_305_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_305_ldest;
        io_diffCommits_info_305_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_305_pdest;
        io_diffCommits_info_306_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_306_ldest;
        io_diffCommits_info_306_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_306_pdest;
        io_diffCommits_info_307_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_307_ldest;
        io_diffCommits_info_307_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_307_pdest;
        io_diffCommits_info_308_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_308_ldest;
        io_diffCommits_info_308_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_308_pdest;
        io_diffCommits_info_309_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_309_ldest;
        io_diffCommits_info_309_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_309_pdest;
        io_diffCommits_info_310_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_310_ldest;
        io_diffCommits_info_310_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_310_pdest;
        io_diffCommits_info_311_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_311_ldest;
        io_diffCommits_info_311_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_311_pdest;
        io_diffCommits_info_312_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_312_ldest;
        io_diffCommits_info_312_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_312_pdest;
        io_diffCommits_info_313_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_313_ldest;
        io_diffCommits_info_313_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_313_pdest;
        io_diffCommits_info_314_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_314_ldest;
        io_diffCommits_info_314_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_314_pdest;
        io_diffCommits_info_315_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_315_ldest;
        io_diffCommits_info_315_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_315_pdest;
        io_diffCommits_info_316_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_316_ldest;
        io_diffCommits_info_316_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_316_pdest;
        io_diffCommits_info_317_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_317_ldest;
        io_diffCommits_info_317_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_317_pdest;
        io_diffCommits_info_318_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_318_ldest;
        io_diffCommits_info_318_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_318_pdest;
        io_diffCommits_info_319_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_319_ldest;
        io_diffCommits_info_319_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_319_pdest;
        io_diffCommits_info_320_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_320_ldest;
        io_diffCommits_info_320_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_320_pdest;
        io_diffCommits_info_321_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_321_ldest;
        io_diffCommits_info_321_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_321_pdest;
        io_diffCommits_info_322_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_322_ldest;
        io_diffCommits_info_322_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_322_pdest;
        io_diffCommits_info_323_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_323_ldest;
        io_diffCommits_info_323_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_323_pdest;
        io_diffCommits_info_324_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_324_ldest;
        io_diffCommits_info_324_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_324_pdest;
        io_diffCommits_info_325_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_325_ldest;
        io_diffCommits_info_325_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_325_pdest;
        io_diffCommits_info_326_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_326_ldest;
        io_diffCommits_info_326_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_326_pdest;
        io_diffCommits_info_327_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_327_ldest;
        io_diffCommits_info_327_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_327_pdest;
        io_diffCommits_info_328_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_328_ldest;
        io_diffCommits_info_328_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_328_pdest;
        io_diffCommits_info_329_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_329_ldest;
        io_diffCommits_info_329_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_329_pdest;
        io_diffCommits_info_330_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_330_ldest;
        io_diffCommits_info_330_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_330_pdest;
        io_diffCommits_info_331_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_331_ldest;
        io_diffCommits_info_331_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_331_pdest;
        io_diffCommits_info_332_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_332_ldest;
        io_diffCommits_info_332_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_332_pdest;
        io_diffCommits_info_333_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_333_ldest;
        io_diffCommits_info_333_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_333_pdest;
        io_diffCommits_info_334_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_334_ldest;
        io_diffCommits_info_334_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_334_pdest;
        io_diffCommits_info_335_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_335_ldest;
        io_diffCommits_info_335_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_335_pdest;
        io_diffCommits_info_336_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_336_ldest;
        io_diffCommits_info_336_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_336_pdest;
        io_diffCommits_info_337_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_337_ldest;
        io_diffCommits_info_337_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_337_pdest;
        io_diffCommits_info_338_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_338_ldest;
        io_diffCommits_info_338_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_338_pdest;
        io_diffCommits_info_339_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_339_ldest;
        io_diffCommits_info_339_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_339_pdest;
        io_diffCommits_info_340_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_340_ldest;
        io_diffCommits_info_340_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_340_pdest;
        io_diffCommits_info_341_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_341_ldest;
        io_diffCommits_info_341_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_341_pdest;
        io_diffCommits_info_342_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_342_ldest;
        io_diffCommits_info_342_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_342_pdest;
        io_diffCommits_info_343_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_343_ldest;
        io_diffCommits_info_343_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_343_pdest;
        io_diffCommits_info_344_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_344_ldest;
        io_diffCommits_info_344_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_344_pdest;
        io_diffCommits_info_345_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_345_ldest;
        io_diffCommits_info_345_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_345_pdest;
        io_diffCommits_info_346_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_346_ldest;
        io_diffCommits_info_346_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_346_pdest;
        io_diffCommits_info_347_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_347_ldest;
        io_diffCommits_info_347_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_347_pdest;
        io_diffCommits_info_348_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_348_ldest;
        io_diffCommits_info_348_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_348_pdest;
        io_diffCommits_info_349_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_349_ldest;
        io_diffCommits_info_349_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_349_pdest;
        io_diffCommits_info_350_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_350_ldest;
        io_diffCommits_info_350_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_350_pdest;
        io_diffCommits_info_351_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_351_ldest;
        io_diffCommits_info_351_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_351_pdest;
        io_diffCommits_info_352_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_352_ldest;
        io_diffCommits_info_352_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_352_pdest;
        io_diffCommits_info_353_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_353_ldest;
        io_diffCommits_info_353_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_353_pdest;
        io_diffCommits_info_354_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_354_ldest;
        io_diffCommits_info_354_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_354_pdest;
        io_diffCommits_info_355_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_355_ldest;
        io_diffCommits_info_355_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_355_pdest;
        io_diffCommits_info_356_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_356_ldest;
        io_diffCommits_info_356_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_356_pdest;
        io_diffCommits_info_357_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_357_ldest;
        io_diffCommits_info_357_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_357_pdest;
        io_diffCommits_info_358_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_358_ldest;
        io_diffCommits_info_358_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_358_pdest;
        io_diffCommits_info_359_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_359_ldest;
        io_diffCommits_info_359_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_359_pdest;
        io_diffCommits_info_360_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_360_ldest;
        io_diffCommits_info_360_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_360_pdest;
        io_diffCommits_info_361_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_361_ldest;
        io_diffCommits_info_361_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_361_pdest;
        io_diffCommits_info_362_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_362_ldest;
        io_diffCommits_info_362_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_362_pdest;
        io_diffCommits_info_363_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_363_ldest;
        io_diffCommits_info_363_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_363_pdest;
        io_diffCommits_info_364_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_364_ldest;
        io_diffCommits_info_364_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_364_pdest;
        io_diffCommits_info_365_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_365_ldest;
        io_diffCommits_info_365_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_365_pdest;
        io_diffCommits_info_366_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_366_ldest;
        io_diffCommits_info_366_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_366_pdest;
        io_diffCommits_info_367_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_367_ldest;
        io_diffCommits_info_367_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_367_pdest;
        io_diffCommits_info_368_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_368_ldest;
        io_diffCommits_info_368_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_368_pdest;
        io_diffCommits_info_369_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_369_ldest;
        io_diffCommits_info_369_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_369_pdest;
        io_diffCommits_info_370_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_370_ldest;
        io_diffCommits_info_370_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_370_pdest;
        io_diffCommits_info_371_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_371_ldest;
        io_diffCommits_info_371_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_371_pdest;
        io_diffCommits_info_372_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_372_ldest;
        io_diffCommits_info_372_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_372_pdest;
        io_diffCommits_info_373_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_373_ldest;
        io_diffCommits_info_373_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_373_pdest;
        io_diffCommits_info_374_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_374_ldest;
        io_diffCommits_info_374_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_374_pdest;
        io_diffCommits_info_375_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_375_ldest;
        io_diffCommits_info_375_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_375_pdest;
        io_diffCommits_info_376_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_376_ldest;
        io_diffCommits_info_376_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_376_pdest;
        io_diffCommits_info_377_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_377_ldest;
        io_diffCommits_info_377_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_377_pdest;
        io_diffCommits_info_378_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_378_ldest;
        io_diffCommits_info_378_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_378_pdest;
        io_diffCommits_info_379_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_379_ldest;
        io_diffCommits_info_379_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_379_pdest;
        io_diffCommits_info_380_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_380_ldest;
        io_diffCommits_info_380_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_380_pdest;
        io_diffCommits_info_381_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_381_ldest;
        io_diffCommits_info_381_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_381_pdest;
        io_diffCommits_info_382_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_382_ldest;
        io_diffCommits_info_382_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_382_pdest;
        io_diffCommits_info_383_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_383_ldest;
        io_diffCommits_info_383_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_383_pdest;
        io_diffCommits_info_384_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_384_ldest;
        io_diffCommits_info_384_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_384_pdest;
        io_diffCommits_info_385_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_385_ldest;
        io_diffCommits_info_385_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_385_pdest;
        io_diffCommits_info_386_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_386_ldest;
        io_diffCommits_info_386_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_386_pdest;
        io_diffCommits_info_387_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_387_ldest;
        io_diffCommits_info_387_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_387_pdest;
        io_diffCommits_info_388_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_388_ldest;
        io_diffCommits_info_388_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_388_pdest;
        io_diffCommits_info_389_ldest = this.vif.mon_mp.mon_cb.io_diffCommits_info_389_ldest;
        io_diffCommits_info_389_pdest = this.vif.mon_mp.mon_cb.io_diffCommits_info_389_pdest;
        io_lsq_scommit = this.vif.mon_mp.mon_cb.io_lsq_scommit;
        io_lsq_pendingMMIOld = this.vif.mon_mp.mon_cb.io_lsq_pendingMMIOld;
        io_lsq_pendingst = this.vif.mon_mp.mon_cb.io_lsq_pendingst;
        io_lsq_pendingPtr_flag = this.vif.mon_mp.mon_cb.io_lsq_pendingPtr_flag;
        io_lsq_pendingPtr_value = this.vif.mon_mp.mon_cb.io_lsq_pendingPtr_value;
        io_robDeqPtr_flag = this.vif.mon_mp.mon_cb.io_robDeqPtr_flag;
        io_robDeqPtr_value = this.vif.mon_mp.mon_cb.io_robDeqPtr_value;
        io_csr_fflags_valid = this.vif.mon_mp.mon_cb.io_csr_fflags_valid;
        io_csr_fflags_bits = this.vif.mon_mp.mon_cb.io_csr_fflags_bits;
        io_csr_vxsat_valid = this.vif.mon_mp.mon_cb.io_csr_vxsat_valid;
        io_csr_vxsat_bits = this.vif.mon_mp.mon_cb.io_csr_vxsat_bits;
        io_csr_vstart_valid = this.vif.mon_mp.mon_cb.io_csr_vstart_valid;
        io_csr_vstart_bits = this.vif.mon_mp.mon_cb.io_csr_vstart_bits;
        io_csr_dirty_fs = this.vif.mon_mp.mon_cb.io_csr_dirty_fs;
        io_csr_dirty_vs = this.vif.mon_mp.mon_cb.io_csr_dirty_vs;
        io_csr_perfinfo_retiredInstr = this.vif.mon_mp.mon_cb.io_csr_perfinfo_retiredInstr;
        io_cpu_halt = this.vif.mon_mp.mon_cb.io_cpu_halt;
        io_wfi_wfiReq = this.vif.mon_mp.mon_cb.io_wfi_wfiReq;
        io_toDecode_isResumeVType = this.vif.mon_mp.mon_cb.io_toDecode_isResumeVType;
        io_toDecode_walkToArchVType = this.vif.mon_mp.mon_cb.io_toDecode_walkToArchVType;
        io_toDecode_walkVType_valid = this.vif.mon_mp.mon_cb.io_toDecode_walkVType_valid;
        io_toDecode_walkVType_bits_illegal = this.vif.mon_mp.mon_cb.io_toDecode_walkVType_bits_illegal;
        io_toDecode_walkVType_bits_vma = this.vif.mon_mp.mon_cb.io_toDecode_walkVType_bits_vma;
        io_toDecode_walkVType_bits_vta = this.vif.mon_mp.mon_cb.io_toDecode_walkVType_bits_vta;
        io_toDecode_walkVType_bits_vsew = this.vif.mon_mp.mon_cb.io_toDecode_walkVType_bits_vsew;
        io_toDecode_walkVType_bits_vlmul = this.vif.mon_mp.mon_cb.io_toDecode_walkVType_bits_vlmul;
        io_toDecode_commitVType_vtype_valid = this.vif.mon_mp.mon_cb.io_toDecode_commitVType_vtype_valid;
        io_toDecode_commitVType_vtype_bits_illegal = this.vif.mon_mp.mon_cb.io_toDecode_commitVType_vtype_bits_illegal;
        io_toDecode_commitVType_vtype_bits_vma = this.vif.mon_mp.mon_cb.io_toDecode_commitVType_vtype_bits_vma;
        io_toDecode_commitVType_vtype_bits_vta = this.vif.mon_mp.mon_cb.io_toDecode_commitVType_vtype_bits_vta;
        io_toDecode_commitVType_vtype_bits_vsew = this.vif.mon_mp.mon_cb.io_toDecode_commitVType_vtype_bits_vsew;
        io_toDecode_commitVType_vtype_bits_vlmul = this.vif.mon_mp.mon_cb.io_toDecode_commitVType_vtype_bits_vlmul;
        io_toDecode_commitVType_hasVsetvl = this.vif.mon_mp.mon_cb.io_toDecode_commitVType_hasVsetvl;
        io_readGPAMemAddr_valid = this.vif.mon_mp.mon_cb.io_readGPAMemAddr_valid;
        io_readGPAMemAddr_bits_ftqPtr_value = this.vif.mon_mp.mon_cb.io_readGPAMemAddr_bits_ftqPtr_value;
        io_readGPAMemAddr_bits_ftqOffset = this.vif.mon_mp.mon_cb.io_readGPAMemAddr_bits_ftqOffset;
        io_toVecExcpMod_logicPhyRegMap_0_valid = this.vif.mon_mp.mon_cb.io_toVecExcpMod_logicPhyRegMap_0_valid;
        io_toVecExcpMod_logicPhyRegMap_0_bits_lreg = this.vif.mon_mp.mon_cb.io_toVecExcpMod_logicPhyRegMap_0_bits_lreg;
        io_toVecExcpMod_logicPhyRegMap_0_bits_preg = this.vif.mon_mp.mon_cb.io_toVecExcpMod_logicPhyRegMap_0_bits_preg;
        io_toVecExcpMod_logicPhyRegMap_1_valid = this.vif.mon_mp.mon_cb.io_toVecExcpMod_logicPhyRegMap_1_valid;
        io_toVecExcpMod_logicPhyRegMap_1_bits_lreg = this.vif.mon_mp.mon_cb.io_toVecExcpMod_logicPhyRegMap_1_bits_lreg;
        io_toVecExcpMod_logicPhyRegMap_1_bits_preg = this.vif.mon_mp.mon_cb.io_toVecExcpMod_logicPhyRegMap_1_bits_preg;
        io_toVecExcpMod_logicPhyRegMap_2_valid = this.vif.mon_mp.mon_cb.io_toVecExcpMod_logicPhyRegMap_2_valid;
        io_toVecExcpMod_logicPhyRegMap_2_bits_lreg = this.vif.mon_mp.mon_cb.io_toVecExcpMod_logicPhyRegMap_2_bits_lreg;
        io_toVecExcpMod_logicPhyRegMap_2_bits_preg = this.vif.mon_mp.mon_cb.io_toVecExcpMod_logicPhyRegMap_2_bits_preg;
        io_toVecExcpMod_logicPhyRegMap_3_valid = this.vif.mon_mp.mon_cb.io_toVecExcpMod_logicPhyRegMap_3_valid;
        io_toVecExcpMod_logicPhyRegMap_3_bits_lreg = this.vif.mon_mp.mon_cb.io_toVecExcpMod_logicPhyRegMap_3_bits_lreg;
        io_toVecExcpMod_logicPhyRegMap_3_bits_preg = this.vif.mon_mp.mon_cb.io_toVecExcpMod_logicPhyRegMap_3_bits_preg;
        io_toVecExcpMod_logicPhyRegMap_4_valid = this.vif.mon_mp.mon_cb.io_toVecExcpMod_logicPhyRegMap_4_valid;
        io_toVecExcpMod_logicPhyRegMap_4_bits_lreg = this.vif.mon_mp.mon_cb.io_toVecExcpMod_logicPhyRegMap_4_bits_lreg;
        io_toVecExcpMod_logicPhyRegMap_4_bits_preg = this.vif.mon_mp.mon_cb.io_toVecExcpMod_logicPhyRegMap_4_bits_preg;
        io_toVecExcpMod_logicPhyRegMap_5_valid = this.vif.mon_mp.mon_cb.io_toVecExcpMod_logicPhyRegMap_5_valid;
        io_toVecExcpMod_logicPhyRegMap_5_bits_lreg = this.vif.mon_mp.mon_cb.io_toVecExcpMod_logicPhyRegMap_5_bits_lreg;
        io_toVecExcpMod_logicPhyRegMap_5_bits_preg = this.vif.mon_mp.mon_cb.io_toVecExcpMod_logicPhyRegMap_5_bits_preg;
        io_toVecExcpMod_excpInfo_valid = this.vif.mon_mp.mon_cb.io_toVecExcpMod_excpInfo_valid;
        io_toVecExcpMod_excpInfo_bits_vstart = this.vif.mon_mp.mon_cb.io_toVecExcpMod_excpInfo_bits_vstart;
        io_toVecExcpMod_excpInfo_bits_vsew = this.vif.mon_mp.mon_cb.io_toVecExcpMod_excpInfo_bits_vsew;
        io_toVecExcpMod_excpInfo_bits_veew = this.vif.mon_mp.mon_cb.io_toVecExcpMod_excpInfo_bits_veew;
        io_toVecExcpMod_excpInfo_bits_vlmul = this.vif.mon_mp.mon_cb.io_toVecExcpMod_excpInfo_bits_vlmul;
        io_toVecExcpMod_excpInfo_bits_nf = this.vif.mon_mp.mon_cb.io_toVecExcpMod_excpInfo_bits_nf;
        io_toVecExcpMod_excpInfo_bits_isStride = this.vif.mon_mp.mon_cb.io_toVecExcpMod_excpInfo_bits_isStride;
        io_toVecExcpMod_excpInfo_bits_isIndexed = this.vif.mon_mp.mon_cb.io_toVecExcpMod_excpInfo_bits_isIndexed;
        io_toVecExcpMod_excpInfo_bits_isWhole = this.vif.mon_mp.mon_cb.io_toVecExcpMod_excpInfo_bits_isWhole;
        io_toVecExcpMod_excpInfo_bits_isVlm = this.vif.mon_mp.mon_cb.io_toVecExcpMod_excpInfo_bits_isVlm;
        io_storeDebugInfo_1_pc = this.vif.mon_mp.mon_cb.io_storeDebugInfo_1_pc;
        io_perf_0_value = this.vif.mon_mp.mon_cb.io_perf_0_value;
        io_perf_1_value = this.vif.mon_mp.mon_cb.io_perf_1_value;
        io_perf_2_value = this.vif.mon_mp.mon_cb.io_perf_2_value;
        io_perf_3_value = this.vif.mon_mp.mon_cb.io_perf_3_value;
        io_perf_4_value = this.vif.mon_mp.mon_cb.io_perf_4_value;
        io_perf_5_value = this.vif.mon_mp.mon_cb.io_perf_5_value;
        io_perf_6_value = this.vif.mon_mp.mon_cb.io_perf_6_value;
        io_perf_7_value = this.vif.mon_mp.mon_cb.io_perf_7_value;
        io_perf_8_value = this.vif.mon_mp.mon_cb.io_perf_8_value;
        io_perf_9_value = this.vif.mon_mp.mon_cb.io_perf_9_value;
        io_perf_10_value = this.vif.mon_mp.mon_cb.io_perf_10_value;
        io_perf_11_value = this.vif.mon_mp.mon_cb.io_perf_11_value;
        io_perf_12_value = this.vif.mon_mp.mon_cb.io_perf_12_value;
        io_perf_13_value = this.vif.mon_mp.mon_cb.io_perf_13_value;
        io_perf_14_value = this.vif.mon_mp.mon_cb.io_perf_14_value;
        io_perf_15_value = this.vif.mon_mp.mon_cb.io_perf_15_value;
        io_perf_16_value = this.vif.mon_mp.mon_cb.io_perf_16_value;
        io_perf_17_value = this.vif.mon_mp.mon_cb.io_perf_17_value;
        io_error_0 = this.vif.mon_mp.mon_cb.io_error_0;

        // if(this.cfg.xz_sw==tcnt_dec_base::ON & this.vif.rst_n==1'b1) begin
        //     `TCNT_CHECK_SIG_XZ(io_enq_canAccept,io_enq_canAccept,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_canAcceptForDispatch,io_enq_canAcceptForDispatch,1);
        //     `TCNT_CHECK_SIG_XZ(io_enq_isEmpty,io_enq_isEmpty,1);
        //     `TCNT_CHECK_SIG_XZ(io_flushOut_valid,io_flushOut_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_flushOut_bits_isRVC,io_flushOut_bits_isRVC,1);
        //     `TCNT_CHECK_SIG_XZ(io_flushOut_bits_robIdx_flag,io_flushOut_bits_robIdx_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_flushOut_bits_robIdx_value,io_flushOut_bits_robIdx_value,8);
        //     `TCNT_CHECK_SIG_XZ(io_flushOut_bits_ftqIdx_flag,io_flushOut_bits_ftqIdx_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_flushOut_bits_ftqIdx_value,io_flushOut_bits_ftqIdx_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_flushOut_bits_ftqOffset,io_flushOut_bits_ftqOffset,4);
        //     `TCNT_CHECK_SIG_XZ(io_flushOut_bits_level,io_flushOut_bits_level,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_valid,io_exception_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_instr,io_exception_bits_instr,32);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_commitType,io_exception_bits_commitType,3);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_exceptionVec_0,io_exception_bits_exceptionVec_0,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_exceptionVec_1,io_exception_bits_exceptionVec_1,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_exceptionVec_2,io_exception_bits_exceptionVec_2,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_exceptionVec_3,io_exception_bits_exceptionVec_3,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_exceptionVec_4,io_exception_bits_exceptionVec_4,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_exceptionVec_5,io_exception_bits_exceptionVec_5,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_exceptionVec_6,io_exception_bits_exceptionVec_6,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_exceptionVec_7,io_exception_bits_exceptionVec_7,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_exceptionVec_8,io_exception_bits_exceptionVec_8,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_exceptionVec_9,io_exception_bits_exceptionVec_9,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_exceptionVec_10,io_exception_bits_exceptionVec_10,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_exceptionVec_11,io_exception_bits_exceptionVec_11,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_exceptionVec_12,io_exception_bits_exceptionVec_12,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_exceptionVec_13,io_exception_bits_exceptionVec_13,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_exceptionVec_14,io_exception_bits_exceptionVec_14,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_exceptionVec_15,io_exception_bits_exceptionVec_15,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_exceptionVec_16,io_exception_bits_exceptionVec_16,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_exceptionVec_17,io_exception_bits_exceptionVec_17,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_exceptionVec_18,io_exception_bits_exceptionVec_18,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_exceptionVec_19,io_exception_bits_exceptionVec_19,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_exceptionVec_20,io_exception_bits_exceptionVec_20,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_exceptionVec_21,io_exception_bits_exceptionVec_21,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_exceptionVec_22,io_exception_bits_exceptionVec_22,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_exceptionVec_23,io_exception_bits_exceptionVec_23,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_isPcBkpt,io_exception_bits_isPcBkpt,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_isFetchMalAddr,io_exception_bits_isFetchMalAddr,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_gpaddr,io_exception_bits_gpaddr,64);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_singleStep,io_exception_bits_singleStep,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_crossPageIPFFix,io_exception_bits_crossPageIPFFix,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_isInterrupt,io_exception_bits_isInterrupt,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_isHls,io_exception_bits_isHls,1);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_trigger,io_exception_bits_trigger,4);
        //     `TCNT_CHECK_SIG_XZ(io_exception_bits_isForVSnonLeafPTE,io_exception_bits_isForVSnonLeafPTE,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_isCommit,io_commits_isCommit,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_commitValid_0,io_commits_commitValid_0,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_commitValid_1,io_commits_commitValid_1,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_commitValid_2,io_commits_commitValid_2,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_commitValid_3,io_commits_commitValid_3,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_commitValid_4,io_commits_commitValid_4,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_commitValid_5,io_commits_commitValid_5,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_commitValid_6,io_commits_commitValid_6,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_commitValid_7,io_commits_commitValid_7,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_isWalk,io_commits_isWalk,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_walkValid_0,io_commits_walkValid_0,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_walkValid_1,io_commits_walkValid_1,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_walkValid_2,io_commits_walkValid_2,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_walkValid_3,io_commits_walkValid_3,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_walkValid_4,io_commits_walkValid_4,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_walkValid_5,io_commits_walkValid_5,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_walkValid_6,io_commits_walkValid_6,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_walkValid_7,io_commits_walkValid_7,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_walk_v,io_commits_info_0_walk_v,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_commit_v,io_commits_info_0_commit_v,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_commit_w,io_commits_info_0_commit_w,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_realDestSize,io_commits_info_0_realDestSize,7);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_interrupt_safe,io_commits_info_0_interrupt_safe,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_wflags,io_commits_info_0_wflags,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_fflags,io_commits_info_0_fflags,5);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_vxsat,io_commits_info_0_vxsat,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_isRVC,io_commits_info_0_isRVC,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_isVset,io_commits_info_0_isVset,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_isHls,io_commits_info_0_isHls,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_isVls,io_commits_info_0_isVls,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_vls,io_commits_info_0_vls,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_mmio,io_commits_info_0_mmio,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_commitType,io_commits_info_0_commitType,3);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_ftqIdx_flag,io_commits_info_0_ftqIdx_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_ftqIdx_value,io_commits_info_0_ftqIdx_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_ftqOffset,io_commits_info_0_ftqOffset,4);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_instrSize,io_commits_info_0_instrSize,3);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_fpWen,io_commits_info_0_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_rfWen,io_commits_info_0_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_needFlush,io_commits_info_0_needFlush,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_traceBlockInPipe_itype,io_commits_info_0_traceBlockInPipe_itype,4);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_traceBlockInPipe_iretire,io_commits_info_0_traceBlockInPipe_iretire,4);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_traceBlockInPipe_ilastsize,io_commits_info_0_traceBlockInPipe_ilastsize,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_debug_pc,io_commits_info_0_debug_pc,50);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_debug_instr,io_commits_info_0_debug_instr,32);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_debug_ldest,io_commits_info_0_debug_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_debug_pdest,io_commits_info_0_debug_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_debug_otherPdest_0,io_commits_info_0_debug_otherPdest_0,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_debug_otherPdest_1,io_commits_info_0_debug_otherPdest_1,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_debug_otherPdest_2,io_commits_info_0_debug_otherPdest_2,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_debug_otherPdest_3,io_commits_info_0_debug_otherPdest_3,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_debug_otherPdest_4,io_commits_info_0_debug_otherPdest_4,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_debug_otherPdest_5,io_commits_info_0_debug_otherPdest_5,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_debug_otherPdest_6,io_commits_info_0_debug_otherPdest_6,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_debug_fuType,io_commits_info_0_debug_fuType,35);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_dirtyFs,io_commits_info_0_dirtyFs,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_0_dirtyVs,io_commits_info_0_dirtyVs,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_walk_v,io_commits_info_1_walk_v,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_commit_v,io_commits_info_1_commit_v,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_commit_w,io_commits_info_1_commit_w,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_realDestSize,io_commits_info_1_realDestSize,7);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_interrupt_safe,io_commits_info_1_interrupt_safe,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_wflags,io_commits_info_1_wflags,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_fflags,io_commits_info_1_fflags,5);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_vxsat,io_commits_info_1_vxsat,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_isRVC,io_commits_info_1_isRVC,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_isVset,io_commits_info_1_isVset,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_isHls,io_commits_info_1_isHls,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_isVls,io_commits_info_1_isVls,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_vls,io_commits_info_1_vls,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_mmio,io_commits_info_1_mmio,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_commitType,io_commits_info_1_commitType,3);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_ftqIdx_flag,io_commits_info_1_ftqIdx_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_ftqIdx_value,io_commits_info_1_ftqIdx_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_ftqOffset,io_commits_info_1_ftqOffset,4);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_instrSize,io_commits_info_1_instrSize,3);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_fpWen,io_commits_info_1_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_rfWen,io_commits_info_1_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_needFlush,io_commits_info_1_needFlush,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_traceBlockInPipe_itype,io_commits_info_1_traceBlockInPipe_itype,4);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_traceBlockInPipe_iretire,io_commits_info_1_traceBlockInPipe_iretire,4);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_traceBlockInPipe_ilastsize,io_commits_info_1_traceBlockInPipe_ilastsize,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_debug_pc,io_commits_info_1_debug_pc,50);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_debug_instr,io_commits_info_1_debug_instr,32);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_debug_ldest,io_commits_info_1_debug_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_debug_pdest,io_commits_info_1_debug_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_debug_otherPdest_0,io_commits_info_1_debug_otherPdest_0,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_debug_otherPdest_1,io_commits_info_1_debug_otherPdest_1,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_debug_otherPdest_2,io_commits_info_1_debug_otherPdest_2,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_debug_otherPdest_3,io_commits_info_1_debug_otherPdest_3,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_debug_otherPdest_4,io_commits_info_1_debug_otherPdest_4,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_debug_otherPdest_5,io_commits_info_1_debug_otherPdest_5,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_debug_otherPdest_6,io_commits_info_1_debug_otherPdest_6,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_debug_fuType,io_commits_info_1_debug_fuType,35);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_dirtyFs,io_commits_info_1_dirtyFs,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_1_dirtyVs,io_commits_info_1_dirtyVs,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_walk_v,io_commits_info_2_walk_v,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_commit_v,io_commits_info_2_commit_v,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_commit_w,io_commits_info_2_commit_w,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_realDestSize,io_commits_info_2_realDestSize,7);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_interrupt_safe,io_commits_info_2_interrupt_safe,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_wflags,io_commits_info_2_wflags,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_fflags,io_commits_info_2_fflags,5);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_vxsat,io_commits_info_2_vxsat,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_isRVC,io_commits_info_2_isRVC,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_isVset,io_commits_info_2_isVset,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_isHls,io_commits_info_2_isHls,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_isVls,io_commits_info_2_isVls,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_vls,io_commits_info_2_vls,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_mmio,io_commits_info_2_mmio,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_commitType,io_commits_info_2_commitType,3);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_ftqIdx_flag,io_commits_info_2_ftqIdx_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_ftqIdx_value,io_commits_info_2_ftqIdx_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_ftqOffset,io_commits_info_2_ftqOffset,4);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_instrSize,io_commits_info_2_instrSize,3);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_fpWen,io_commits_info_2_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_rfWen,io_commits_info_2_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_needFlush,io_commits_info_2_needFlush,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_traceBlockInPipe_itype,io_commits_info_2_traceBlockInPipe_itype,4);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_traceBlockInPipe_iretire,io_commits_info_2_traceBlockInPipe_iretire,4);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_traceBlockInPipe_ilastsize,io_commits_info_2_traceBlockInPipe_ilastsize,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_debug_pc,io_commits_info_2_debug_pc,50);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_debug_instr,io_commits_info_2_debug_instr,32);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_debug_ldest,io_commits_info_2_debug_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_debug_pdest,io_commits_info_2_debug_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_debug_otherPdest_0,io_commits_info_2_debug_otherPdest_0,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_debug_otherPdest_1,io_commits_info_2_debug_otherPdest_1,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_debug_otherPdest_2,io_commits_info_2_debug_otherPdest_2,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_debug_otherPdest_3,io_commits_info_2_debug_otherPdest_3,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_debug_otherPdest_4,io_commits_info_2_debug_otherPdest_4,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_debug_otherPdest_5,io_commits_info_2_debug_otherPdest_5,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_debug_otherPdest_6,io_commits_info_2_debug_otherPdest_6,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_debug_fuType,io_commits_info_2_debug_fuType,35);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_dirtyFs,io_commits_info_2_dirtyFs,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_2_dirtyVs,io_commits_info_2_dirtyVs,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_walk_v,io_commits_info_3_walk_v,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_commit_v,io_commits_info_3_commit_v,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_commit_w,io_commits_info_3_commit_w,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_realDestSize,io_commits_info_3_realDestSize,7);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_interrupt_safe,io_commits_info_3_interrupt_safe,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_wflags,io_commits_info_3_wflags,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_fflags,io_commits_info_3_fflags,5);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_vxsat,io_commits_info_3_vxsat,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_isRVC,io_commits_info_3_isRVC,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_isVset,io_commits_info_3_isVset,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_isHls,io_commits_info_3_isHls,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_isVls,io_commits_info_3_isVls,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_vls,io_commits_info_3_vls,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_mmio,io_commits_info_3_mmio,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_commitType,io_commits_info_3_commitType,3);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_ftqIdx_flag,io_commits_info_3_ftqIdx_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_ftqIdx_value,io_commits_info_3_ftqIdx_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_ftqOffset,io_commits_info_3_ftqOffset,4);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_instrSize,io_commits_info_3_instrSize,3);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_fpWen,io_commits_info_3_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_rfWen,io_commits_info_3_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_needFlush,io_commits_info_3_needFlush,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_traceBlockInPipe_itype,io_commits_info_3_traceBlockInPipe_itype,4);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_traceBlockInPipe_iretire,io_commits_info_3_traceBlockInPipe_iretire,4);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_traceBlockInPipe_ilastsize,io_commits_info_3_traceBlockInPipe_ilastsize,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_debug_pc,io_commits_info_3_debug_pc,50);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_debug_instr,io_commits_info_3_debug_instr,32);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_debug_ldest,io_commits_info_3_debug_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_debug_pdest,io_commits_info_3_debug_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_debug_otherPdest_0,io_commits_info_3_debug_otherPdest_0,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_debug_otherPdest_1,io_commits_info_3_debug_otherPdest_1,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_debug_otherPdest_2,io_commits_info_3_debug_otherPdest_2,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_debug_otherPdest_3,io_commits_info_3_debug_otherPdest_3,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_debug_otherPdest_4,io_commits_info_3_debug_otherPdest_4,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_debug_otherPdest_5,io_commits_info_3_debug_otherPdest_5,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_debug_otherPdest_6,io_commits_info_3_debug_otherPdest_6,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_debug_fuType,io_commits_info_3_debug_fuType,35);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_dirtyFs,io_commits_info_3_dirtyFs,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_3_dirtyVs,io_commits_info_3_dirtyVs,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_walk_v,io_commits_info_4_walk_v,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_commit_v,io_commits_info_4_commit_v,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_commit_w,io_commits_info_4_commit_w,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_realDestSize,io_commits_info_4_realDestSize,7);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_interrupt_safe,io_commits_info_4_interrupt_safe,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_wflags,io_commits_info_4_wflags,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_fflags,io_commits_info_4_fflags,5);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_vxsat,io_commits_info_4_vxsat,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_isRVC,io_commits_info_4_isRVC,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_isVset,io_commits_info_4_isVset,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_isHls,io_commits_info_4_isHls,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_isVls,io_commits_info_4_isVls,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_vls,io_commits_info_4_vls,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_mmio,io_commits_info_4_mmio,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_commitType,io_commits_info_4_commitType,3);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_ftqIdx_flag,io_commits_info_4_ftqIdx_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_ftqIdx_value,io_commits_info_4_ftqIdx_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_ftqOffset,io_commits_info_4_ftqOffset,4);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_instrSize,io_commits_info_4_instrSize,3);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_fpWen,io_commits_info_4_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_rfWen,io_commits_info_4_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_needFlush,io_commits_info_4_needFlush,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_traceBlockInPipe_itype,io_commits_info_4_traceBlockInPipe_itype,4);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_traceBlockInPipe_iretire,io_commits_info_4_traceBlockInPipe_iretire,4);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_traceBlockInPipe_ilastsize,io_commits_info_4_traceBlockInPipe_ilastsize,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_debug_pc,io_commits_info_4_debug_pc,50);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_debug_instr,io_commits_info_4_debug_instr,32);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_debug_ldest,io_commits_info_4_debug_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_debug_pdest,io_commits_info_4_debug_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_debug_otherPdest_0,io_commits_info_4_debug_otherPdest_0,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_debug_otherPdest_1,io_commits_info_4_debug_otherPdest_1,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_debug_otherPdest_2,io_commits_info_4_debug_otherPdest_2,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_debug_otherPdest_3,io_commits_info_4_debug_otherPdest_3,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_debug_otherPdest_4,io_commits_info_4_debug_otherPdest_4,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_debug_otherPdest_5,io_commits_info_4_debug_otherPdest_5,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_debug_otherPdest_6,io_commits_info_4_debug_otherPdest_6,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_debug_fuType,io_commits_info_4_debug_fuType,35);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_dirtyFs,io_commits_info_4_dirtyFs,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_4_dirtyVs,io_commits_info_4_dirtyVs,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_walk_v,io_commits_info_5_walk_v,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_commit_v,io_commits_info_5_commit_v,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_commit_w,io_commits_info_5_commit_w,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_realDestSize,io_commits_info_5_realDestSize,7);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_interrupt_safe,io_commits_info_5_interrupt_safe,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_wflags,io_commits_info_5_wflags,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_fflags,io_commits_info_5_fflags,5);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_vxsat,io_commits_info_5_vxsat,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_isRVC,io_commits_info_5_isRVC,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_isVset,io_commits_info_5_isVset,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_isHls,io_commits_info_5_isHls,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_isVls,io_commits_info_5_isVls,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_vls,io_commits_info_5_vls,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_mmio,io_commits_info_5_mmio,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_commitType,io_commits_info_5_commitType,3);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_ftqIdx_flag,io_commits_info_5_ftqIdx_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_ftqIdx_value,io_commits_info_5_ftqIdx_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_ftqOffset,io_commits_info_5_ftqOffset,4);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_instrSize,io_commits_info_5_instrSize,3);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_fpWen,io_commits_info_5_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_rfWen,io_commits_info_5_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_needFlush,io_commits_info_5_needFlush,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_traceBlockInPipe_itype,io_commits_info_5_traceBlockInPipe_itype,4);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_traceBlockInPipe_iretire,io_commits_info_5_traceBlockInPipe_iretire,4);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_traceBlockInPipe_ilastsize,io_commits_info_5_traceBlockInPipe_ilastsize,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_debug_pc,io_commits_info_5_debug_pc,50);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_debug_instr,io_commits_info_5_debug_instr,32);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_debug_ldest,io_commits_info_5_debug_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_debug_pdest,io_commits_info_5_debug_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_debug_otherPdest_0,io_commits_info_5_debug_otherPdest_0,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_debug_otherPdest_1,io_commits_info_5_debug_otherPdest_1,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_debug_otherPdest_2,io_commits_info_5_debug_otherPdest_2,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_debug_otherPdest_3,io_commits_info_5_debug_otherPdest_3,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_debug_otherPdest_4,io_commits_info_5_debug_otherPdest_4,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_debug_otherPdest_5,io_commits_info_5_debug_otherPdest_5,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_debug_otherPdest_6,io_commits_info_5_debug_otherPdest_6,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_debug_fuType,io_commits_info_5_debug_fuType,35);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_dirtyFs,io_commits_info_5_dirtyFs,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_5_dirtyVs,io_commits_info_5_dirtyVs,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_walk_v,io_commits_info_6_walk_v,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_commit_v,io_commits_info_6_commit_v,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_commit_w,io_commits_info_6_commit_w,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_realDestSize,io_commits_info_6_realDestSize,7);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_interrupt_safe,io_commits_info_6_interrupt_safe,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_wflags,io_commits_info_6_wflags,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_fflags,io_commits_info_6_fflags,5);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_vxsat,io_commits_info_6_vxsat,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_isRVC,io_commits_info_6_isRVC,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_isVset,io_commits_info_6_isVset,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_isHls,io_commits_info_6_isHls,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_isVls,io_commits_info_6_isVls,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_vls,io_commits_info_6_vls,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_mmio,io_commits_info_6_mmio,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_commitType,io_commits_info_6_commitType,3);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_ftqIdx_flag,io_commits_info_6_ftqIdx_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_ftqIdx_value,io_commits_info_6_ftqIdx_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_ftqOffset,io_commits_info_6_ftqOffset,4);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_instrSize,io_commits_info_6_instrSize,3);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_fpWen,io_commits_info_6_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_rfWen,io_commits_info_6_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_needFlush,io_commits_info_6_needFlush,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_traceBlockInPipe_itype,io_commits_info_6_traceBlockInPipe_itype,4);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_traceBlockInPipe_iretire,io_commits_info_6_traceBlockInPipe_iretire,4);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_traceBlockInPipe_ilastsize,io_commits_info_6_traceBlockInPipe_ilastsize,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_debug_pc,io_commits_info_6_debug_pc,50);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_debug_instr,io_commits_info_6_debug_instr,32);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_debug_ldest,io_commits_info_6_debug_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_debug_pdest,io_commits_info_6_debug_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_debug_otherPdest_0,io_commits_info_6_debug_otherPdest_0,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_debug_otherPdest_1,io_commits_info_6_debug_otherPdest_1,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_debug_otherPdest_2,io_commits_info_6_debug_otherPdest_2,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_debug_otherPdest_3,io_commits_info_6_debug_otherPdest_3,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_debug_otherPdest_4,io_commits_info_6_debug_otherPdest_4,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_debug_otherPdest_5,io_commits_info_6_debug_otherPdest_5,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_debug_otherPdest_6,io_commits_info_6_debug_otherPdest_6,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_debug_fuType,io_commits_info_6_debug_fuType,35);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_dirtyFs,io_commits_info_6_dirtyFs,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_6_dirtyVs,io_commits_info_6_dirtyVs,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_walk_v,io_commits_info_7_walk_v,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_commit_v,io_commits_info_7_commit_v,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_commit_w,io_commits_info_7_commit_w,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_realDestSize,io_commits_info_7_realDestSize,7);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_interrupt_safe,io_commits_info_7_interrupt_safe,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_wflags,io_commits_info_7_wflags,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_fflags,io_commits_info_7_fflags,5);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_vxsat,io_commits_info_7_vxsat,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_isRVC,io_commits_info_7_isRVC,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_isVset,io_commits_info_7_isVset,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_isHls,io_commits_info_7_isHls,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_isVls,io_commits_info_7_isVls,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_vls,io_commits_info_7_vls,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_mmio,io_commits_info_7_mmio,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_commitType,io_commits_info_7_commitType,3);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_ftqIdx_flag,io_commits_info_7_ftqIdx_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_ftqIdx_value,io_commits_info_7_ftqIdx_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_ftqOffset,io_commits_info_7_ftqOffset,4);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_instrSize,io_commits_info_7_instrSize,3);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_fpWen,io_commits_info_7_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_rfWen,io_commits_info_7_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_needFlush,io_commits_info_7_needFlush,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_traceBlockInPipe_itype,io_commits_info_7_traceBlockInPipe_itype,4);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_traceBlockInPipe_iretire,io_commits_info_7_traceBlockInPipe_iretire,4);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_traceBlockInPipe_ilastsize,io_commits_info_7_traceBlockInPipe_ilastsize,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_debug_pc,io_commits_info_7_debug_pc,50);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_debug_instr,io_commits_info_7_debug_instr,32);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_debug_ldest,io_commits_info_7_debug_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_debug_pdest,io_commits_info_7_debug_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_debug_otherPdest_0,io_commits_info_7_debug_otherPdest_0,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_debug_otherPdest_1,io_commits_info_7_debug_otherPdest_1,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_debug_otherPdest_2,io_commits_info_7_debug_otherPdest_2,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_debug_otherPdest_3,io_commits_info_7_debug_otherPdest_3,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_debug_otherPdest_4,io_commits_info_7_debug_otherPdest_4,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_debug_otherPdest_5,io_commits_info_7_debug_otherPdest_5,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_debug_otherPdest_6,io_commits_info_7_debug_otherPdest_6,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_debug_fuType,io_commits_info_7_debug_fuType,35);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_dirtyFs,io_commits_info_7_dirtyFs,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_info_7_dirtyVs,io_commits_info_7_dirtyVs,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_robIdx_0_flag,io_commits_robIdx_0_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_robIdx_0_value,io_commits_robIdx_0_value,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_robIdx_1_flag,io_commits_robIdx_1_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_robIdx_1_value,io_commits_robIdx_1_value,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_robIdx_2_flag,io_commits_robIdx_2_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_robIdx_2_value,io_commits_robIdx_2_value,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_robIdx_3_flag,io_commits_robIdx_3_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_robIdx_3_value,io_commits_robIdx_3_value,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_robIdx_4_flag,io_commits_robIdx_4_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_robIdx_4_value,io_commits_robIdx_4_value,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_robIdx_5_flag,io_commits_robIdx_5_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_robIdx_5_value,io_commits_robIdx_5_value,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_robIdx_6_flag,io_commits_robIdx_6_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_robIdx_6_value,io_commits_robIdx_6_value,8);
        //     `TCNT_CHECK_SIG_XZ(io_commits_robIdx_7_flag,io_commits_robIdx_7_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_commits_robIdx_7_value,io_commits_robIdx_7_value,8);
        //     `TCNT_CHECK_SIG_XZ(io_trace_blockCommit,io_trace_blockCommit,1);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_0_valid,io_trace_traceCommitInfo_blocks_0_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value,io_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_0_bits_ftqOffset,io_trace_traceCommitInfo_blocks_0_bits_ftqOffset,4);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype,io_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype,4);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire,io_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire,4);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize,io_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize,1);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_1_valid,io_trace_traceCommitInfo_blocks_1_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value,io_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_1_bits_ftqOffset,io_trace_traceCommitInfo_blocks_1_bits_ftqOffset,4);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype,io_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype,4);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire,io_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire,4);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize,io_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize,1);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_2_valid,io_trace_traceCommitInfo_blocks_2_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value,io_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_2_bits_ftqOffset,io_trace_traceCommitInfo_blocks_2_bits_ftqOffset,4);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype,io_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype,4);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire,io_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire,4);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize,io_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize,1);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_3_valid,io_trace_traceCommitInfo_blocks_3_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value,io_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_3_bits_ftqOffset,io_trace_traceCommitInfo_blocks_3_bits_ftqOffset,4);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype,io_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype,4);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire,io_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire,4);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize,io_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize,1);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_4_valid,io_trace_traceCommitInfo_blocks_4_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value,io_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_4_bits_ftqOffset,io_trace_traceCommitInfo_blocks_4_bits_ftqOffset,4);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype,io_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype,4);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire,io_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire,4);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize,io_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize,1);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_5_valid,io_trace_traceCommitInfo_blocks_5_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value,io_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_5_bits_ftqOffset,io_trace_traceCommitInfo_blocks_5_bits_ftqOffset,4);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype,io_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype,4);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire,io_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire,4);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize,io_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize,1);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_6_valid,io_trace_traceCommitInfo_blocks_6_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value,io_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_6_bits_ftqOffset,io_trace_traceCommitInfo_blocks_6_bits_ftqOffset,4);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype,io_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype,4);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire,io_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire,4);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize,io_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize,1);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_7_valid,io_trace_traceCommitInfo_blocks_7_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value,io_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_7_bits_ftqOffset,io_trace_traceCommitInfo_blocks_7_bits_ftqOffset,4);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype,io_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype,4);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire,io_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire,4);
        //     `TCNT_CHECK_SIG_XZ(io_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize,io_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_isCommit,io_rabCommits_isCommit,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_commitValid_0,io_rabCommits_commitValid_0,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_commitValid_1,io_rabCommits_commitValid_1,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_commitValid_2,io_rabCommits_commitValid_2,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_commitValid_3,io_rabCommits_commitValid_3,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_commitValid_4,io_rabCommits_commitValid_4,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_commitValid_5,io_rabCommits_commitValid_5,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_isWalk,io_rabCommits_isWalk,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_walkValid_0,io_rabCommits_walkValid_0,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_walkValid_1,io_rabCommits_walkValid_1,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_walkValid_2,io_rabCommits_walkValid_2,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_walkValid_3,io_rabCommits_walkValid_3,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_walkValid_4,io_rabCommits_walkValid_4,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_walkValid_5,io_rabCommits_walkValid_5,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_0_ldest,io_rabCommits_info_0_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_0_pdest,io_rabCommits_info_0_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_0_rfWen,io_rabCommits_info_0_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_0_fpWen,io_rabCommits_info_0_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_0_vecWen,io_rabCommits_info_0_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_0_v0Wen,io_rabCommits_info_0_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_0_vlWen,io_rabCommits_info_0_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_0_isMove,io_rabCommits_info_0_isMove,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_1_ldest,io_rabCommits_info_1_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_1_pdest,io_rabCommits_info_1_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_1_rfWen,io_rabCommits_info_1_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_1_fpWen,io_rabCommits_info_1_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_1_vecWen,io_rabCommits_info_1_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_1_v0Wen,io_rabCommits_info_1_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_1_vlWen,io_rabCommits_info_1_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_1_isMove,io_rabCommits_info_1_isMove,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_2_ldest,io_rabCommits_info_2_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_2_pdest,io_rabCommits_info_2_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_2_rfWen,io_rabCommits_info_2_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_2_fpWen,io_rabCommits_info_2_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_2_vecWen,io_rabCommits_info_2_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_2_v0Wen,io_rabCommits_info_2_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_2_vlWen,io_rabCommits_info_2_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_2_isMove,io_rabCommits_info_2_isMove,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_3_ldest,io_rabCommits_info_3_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_3_pdest,io_rabCommits_info_3_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_3_rfWen,io_rabCommits_info_3_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_3_fpWen,io_rabCommits_info_3_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_3_vecWen,io_rabCommits_info_3_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_3_v0Wen,io_rabCommits_info_3_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_3_vlWen,io_rabCommits_info_3_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_3_isMove,io_rabCommits_info_3_isMove,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_4_ldest,io_rabCommits_info_4_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_4_pdest,io_rabCommits_info_4_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_4_rfWen,io_rabCommits_info_4_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_4_fpWen,io_rabCommits_info_4_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_4_vecWen,io_rabCommits_info_4_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_4_v0Wen,io_rabCommits_info_4_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_4_vlWen,io_rabCommits_info_4_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_4_isMove,io_rabCommits_info_4_isMove,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_5_ldest,io_rabCommits_info_5_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_5_pdest,io_rabCommits_info_5_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_5_rfWen,io_rabCommits_info_5_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_5_fpWen,io_rabCommits_info_5_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_5_vecWen,io_rabCommits_info_5_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_5_v0Wen,io_rabCommits_info_5_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_5_vlWen,io_rabCommits_info_5_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_rabCommits_info_5_isMove,io_rabCommits_info_5_isMove,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_0,io_diffCommits_commitValid_0,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_1,io_diffCommits_commitValid_1,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_2,io_diffCommits_commitValid_2,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_3,io_diffCommits_commitValid_3,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_4,io_diffCommits_commitValid_4,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_5,io_diffCommits_commitValid_5,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_6,io_diffCommits_commitValid_6,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_7,io_diffCommits_commitValid_7,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_8,io_diffCommits_commitValid_8,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_9,io_diffCommits_commitValid_9,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_10,io_diffCommits_commitValid_10,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_11,io_diffCommits_commitValid_11,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_12,io_diffCommits_commitValid_12,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_13,io_diffCommits_commitValid_13,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_14,io_diffCommits_commitValid_14,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_15,io_diffCommits_commitValid_15,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_16,io_diffCommits_commitValid_16,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_17,io_diffCommits_commitValid_17,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_18,io_diffCommits_commitValid_18,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_19,io_diffCommits_commitValid_19,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_20,io_diffCommits_commitValid_20,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_21,io_diffCommits_commitValid_21,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_22,io_diffCommits_commitValid_22,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_23,io_diffCommits_commitValid_23,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_24,io_diffCommits_commitValid_24,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_25,io_diffCommits_commitValid_25,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_26,io_diffCommits_commitValid_26,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_27,io_diffCommits_commitValid_27,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_28,io_diffCommits_commitValid_28,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_29,io_diffCommits_commitValid_29,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_30,io_diffCommits_commitValid_30,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_31,io_diffCommits_commitValid_31,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_32,io_diffCommits_commitValid_32,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_33,io_diffCommits_commitValid_33,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_34,io_diffCommits_commitValid_34,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_35,io_diffCommits_commitValid_35,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_36,io_diffCommits_commitValid_36,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_37,io_diffCommits_commitValid_37,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_38,io_diffCommits_commitValid_38,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_39,io_diffCommits_commitValid_39,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_40,io_diffCommits_commitValid_40,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_41,io_diffCommits_commitValid_41,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_42,io_diffCommits_commitValid_42,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_43,io_diffCommits_commitValid_43,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_44,io_diffCommits_commitValid_44,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_45,io_diffCommits_commitValid_45,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_46,io_diffCommits_commitValid_46,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_47,io_diffCommits_commitValid_47,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_48,io_diffCommits_commitValid_48,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_49,io_diffCommits_commitValid_49,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_50,io_diffCommits_commitValid_50,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_51,io_diffCommits_commitValid_51,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_52,io_diffCommits_commitValid_52,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_53,io_diffCommits_commitValid_53,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_54,io_diffCommits_commitValid_54,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_55,io_diffCommits_commitValid_55,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_56,io_diffCommits_commitValid_56,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_57,io_diffCommits_commitValid_57,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_58,io_diffCommits_commitValid_58,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_59,io_diffCommits_commitValid_59,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_60,io_diffCommits_commitValid_60,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_61,io_diffCommits_commitValid_61,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_62,io_diffCommits_commitValid_62,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_63,io_diffCommits_commitValid_63,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_64,io_diffCommits_commitValid_64,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_65,io_diffCommits_commitValid_65,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_66,io_diffCommits_commitValid_66,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_67,io_diffCommits_commitValid_67,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_68,io_diffCommits_commitValid_68,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_69,io_diffCommits_commitValid_69,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_70,io_diffCommits_commitValid_70,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_71,io_diffCommits_commitValid_71,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_72,io_diffCommits_commitValid_72,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_73,io_diffCommits_commitValid_73,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_74,io_diffCommits_commitValid_74,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_75,io_diffCommits_commitValid_75,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_76,io_diffCommits_commitValid_76,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_77,io_diffCommits_commitValid_77,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_78,io_diffCommits_commitValid_78,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_79,io_diffCommits_commitValid_79,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_80,io_diffCommits_commitValid_80,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_81,io_diffCommits_commitValid_81,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_82,io_diffCommits_commitValid_82,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_83,io_diffCommits_commitValid_83,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_84,io_diffCommits_commitValid_84,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_85,io_diffCommits_commitValid_85,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_86,io_diffCommits_commitValid_86,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_87,io_diffCommits_commitValid_87,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_88,io_diffCommits_commitValid_88,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_89,io_diffCommits_commitValid_89,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_90,io_diffCommits_commitValid_90,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_91,io_diffCommits_commitValid_91,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_92,io_diffCommits_commitValid_92,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_93,io_diffCommits_commitValid_93,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_94,io_diffCommits_commitValid_94,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_95,io_diffCommits_commitValid_95,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_96,io_diffCommits_commitValid_96,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_97,io_diffCommits_commitValid_97,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_98,io_diffCommits_commitValid_98,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_99,io_diffCommits_commitValid_99,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_100,io_diffCommits_commitValid_100,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_101,io_diffCommits_commitValid_101,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_102,io_diffCommits_commitValid_102,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_103,io_diffCommits_commitValid_103,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_104,io_diffCommits_commitValid_104,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_105,io_diffCommits_commitValid_105,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_106,io_diffCommits_commitValid_106,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_107,io_diffCommits_commitValid_107,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_108,io_diffCommits_commitValid_108,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_109,io_diffCommits_commitValid_109,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_110,io_diffCommits_commitValid_110,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_111,io_diffCommits_commitValid_111,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_112,io_diffCommits_commitValid_112,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_113,io_diffCommits_commitValid_113,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_114,io_diffCommits_commitValid_114,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_115,io_diffCommits_commitValid_115,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_116,io_diffCommits_commitValid_116,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_117,io_diffCommits_commitValid_117,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_118,io_diffCommits_commitValid_118,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_119,io_diffCommits_commitValid_119,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_120,io_diffCommits_commitValid_120,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_121,io_diffCommits_commitValid_121,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_122,io_diffCommits_commitValid_122,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_123,io_diffCommits_commitValid_123,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_124,io_diffCommits_commitValid_124,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_125,io_diffCommits_commitValid_125,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_126,io_diffCommits_commitValid_126,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_127,io_diffCommits_commitValid_127,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_128,io_diffCommits_commitValid_128,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_129,io_diffCommits_commitValid_129,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_130,io_diffCommits_commitValid_130,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_131,io_diffCommits_commitValid_131,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_132,io_diffCommits_commitValid_132,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_133,io_diffCommits_commitValid_133,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_134,io_diffCommits_commitValid_134,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_135,io_diffCommits_commitValid_135,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_136,io_diffCommits_commitValid_136,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_137,io_diffCommits_commitValid_137,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_138,io_diffCommits_commitValid_138,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_139,io_diffCommits_commitValid_139,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_140,io_diffCommits_commitValid_140,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_141,io_diffCommits_commitValid_141,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_142,io_diffCommits_commitValid_142,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_143,io_diffCommits_commitValid_143,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_144,io_diffCommits_commitValid_144,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_145,io_diffCommits_commitValid_145,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_146,io_diffCommits_commitValid_146,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_147,io_diffCommits_commitValid_147,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_148,io_diffCommits_commitValid_148,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_149,io_diffCommits_commitValid_149,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_150,io_diffCommits_commitValid_150,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_151,io_diffCommits_commitValid_151,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_152,io_diffCommits_commitValid_152,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_153,io_diffCommits_commitValid_153,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_154,io_diffCommits_commitValid_154,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_155,io_diffCommits_commitValid_155,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_156,io_diffCommits_commitValid_156,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_157,io_diffCommits_commitValid_157,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_158,io_diffCommits_commitValid_158,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_159,io_diffCommits_commitValid_159,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_160,io_diffCommits_commitValid_160,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_161,io_diffCommits_commitValid_161,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_162,io_diffCommits_commitValid_162,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_163,io_diffCommits_commitValid_163,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_164,io_diffCommits_commitValid_164,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_165,io_diffCommits_commitValid_165,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_166,io_diffCommits_commitValid_166,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_167,io_diffCommits_commitValid_167,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_168,io_diffCommits_commitValid_168,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_169,io_diffCommits_commitValid_169,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_170,io_diffCommits_commitValid_170,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_171,io_diffCommits_commitValid_171,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_172,io_diffCommits_commitValid_172,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_173,io_diffCommits_commitValid_173,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_174,io_diffCommits_commitValid_174,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_175,io_diffCommits_commitValid_175,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_176,io_diffCommits_commitValid_176,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_177,io_diffCommits_commitValid_177,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_178,io_diffCommits_commitValid_178,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_179,io_diffCommits_commitValid_179,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_180,io_diffCommits_commitValid_180,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_181,io_diffCommits_commitValid_181,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_182,io_diffCommits_commitValid_182,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_183,io_diffCommits_commitValid_183,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_184,io_diffCommits_commitValid_184,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_185,io_diffCommits_commitValid_185,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_186,io_diffCommits_commitValid_186,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_187,io_diffCommits_commitValid_187,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_188,io_diffCommits_commitValid_188,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_189,io_diffCommits_commitValid_189,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_190,io_diffCommits_commitValid_190,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_191,io_diffCommits_commitValid_191,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_192,io_diffCommits_commitValid_192,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_193,io_diffCommits_commitValid_193,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_194,io_diffCommits_commitValid_194,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_195,io_diffCommits_commitValid_195,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_196,io_diffCommits_commitValid_196,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_197,io_diffCommits_commitValid_197,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_198,io_diffCommits_commitValid_198,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_199,io_diffCommits_commitValid_199,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_200,io_diffCommits_commitValid_200,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_201,io_diffCommits_commitValid_201,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_202,io_diffCommits_commitValid_202,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_203,io_diffCommits_commitValid_203,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_204,io_diffCommits_commitValid_204,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_205,io_diffCommits_commitValid_205,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_206,io_diffCommits_commitValid_206,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_207,io_diffCommits_commitValid_207,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_208,io_diffCommits_commitValid_208,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_209,io_diffCommits_commitValid_209,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_210,io_diffCommits_commitValid_210,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_211,io_diffCommits_commitValid_211,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_212,io_diffCommits_commitValid_212,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_213,io_diffCommits_commitValid_213,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_214,io_diffCommits_commitValid_214,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_215,io_diffCommits_commitValid_215,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_216,io_diffCommits_commitValid_216,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_217,io_diffCommits_commitValid_217,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_218,io_diffCommits_commitValid_218,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_219,io_diffCommits_commitValid_219,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_220,io_diffCommits_commitValid_220,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_221,io_diffCommits_commitValid_221,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_222,io_diffCommits_commitValid_222,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_223,io_diffCommits_commitValid_223,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_224,io_diffCommits_commitValid_224,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_225,io_diffCommits_commitValid_225,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_226,io_diffCommits_commitValid_226,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_227,io_diffCommits_commitValid_227,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_228,io_diffCommits_commitValid_228,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_229,io_diffCommits_commitValid_229,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_230,io_diffCommits_commitValid_230,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_231,io_diffCommits_commitValid_231,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_232,io_diffCommits_commitValid_232,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_233,io_diffCommits_commitValid_233,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_234,io_diffCommits_commitValid_234,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_235,io_diffCommits_commitValid_235,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_236,io_diffCommits_commitValid_236,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_237,io_diffCommits_commitValid_237,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_238,io_diffCommits_commitValid_238,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_239,io_diffCommits_commitValid_239,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_240,io_diffCommits_commitValid_240,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_241,io_diffCommits_commitValid_241,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_242,io_diffCommits_commitValid_242,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_243,io_diffCommits_commitValid_243,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_244,io_diffCommits_commitValid_244,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_245,io_diffCommits_commitValid_245,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_246,io_diffCommits_commitValid_246,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_247,io_diffCommits_commitValid_247,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_248,io_diffCommits_commitValid_248,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_249,io_diffCommits_commitValid_249,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_250,io_diffCommits_commitValid_250,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_251,io_diffCommits_commitValid_251,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_252,io_diffCommits_commitValid_252,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_253,io_diffCommits_commitValid_253,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_commitValid_254,io_diffCommits_commitValid_254,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_0_ldest,io_diffCommits_info_0_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_0_pdest,io_diffCommits_info_0_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_0_rfWen,io_diffCommits_info_0_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_0_fpWen,io_diffCommits_info_0_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_0_vecWen,io_diffCommits_info_0_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_0_v0Wen,io_diffCommits_info_0_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_0_vlWen,io_diffCommits_info_0_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_1_ldest,io_diffCommits_info_1_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_1_pdest,io_diffCommits_info_1_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_1_rfWen,io_diffCommits_info_1_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_1_fpWen,io_diffCommits_info_1_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_1_vecWen,io_diffCommits_info_1_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_1_v0Wen,io_diffCommits_info_1_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_1_vlWen,io_diffCommits_info_1_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_2_ldest,io_diffCommits_info_2_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_2_pdest,io_diffCommits_info_2_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_2_rfWen,io_diffCommits_info_2_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_2_fpWen,io_diffCommits_info_2_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_2_vecWen,io_diffCommits_info_2_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_2_v0Wen,io_diffCommits_info_2_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_2_vlWen,io_diffCommits_info_2_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_3_ldest,io_diffCommits_info_3_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_3_pdest,io_diffCommits_info_3_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_3_rfWen,io_diffCommits_info_3_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_3_fpWen,io_diffCommits_info_3_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_3_vecWen,io_diffCommits_info_3_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_3_v0Wen,io_diffCommits_info_3_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_3_vlWen,io_diffCommits_info_3_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_4_ldest,io_diffCommits_info_4_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_4_pdest,io_diffCommits_info_4_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_4_rfWen,io_diffCommits_info_4_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_4_fpWen,io_diffCommits_info_4_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_4_vecWen,io_diffCommits_info_4_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_4_v0Wen,io_diffCommits_info_4_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_4_vlWen,io_diffCommits_info_4_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_5_ldest,io_diffCommits_info_5_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_5_pdest,io_diffCommits_info_5_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_5_rfWen,io_diffCommits_info_5_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_5_fpWen,io_diffCommits_info_5_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_5_vecWen,io_diffCommits_info_5_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_5_v0Wen,io_diffCommits_info_5_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_5_vlWen,io_diffCommits_info_5_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_6_ldest,io_diffCommits_info_6_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_6_pdest,io_diffCommits_info_6_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_6_rfWen,io_diffCommits_info_6_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_6_fpWen,io_diffCommits_info_6_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_6_vecWen,io_diffCommits_info_6_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_6_v0Wen,io_diffCommits_info_6_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_6_vlWen,io_diffCommits_info_6_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_7_ldest,io_diffCommits_info_7_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_7_pdest,io_diffCommits_info_7_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_7_rfWen,io_diffCommits_info_7_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_7_fpWen,io_diffCommits_info_7_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_7_vecWen,io_diffCommits_info_7_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_7_v0Wen,io_diffCommits_info_7_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_7_vlWen,io_diffCommits_info_7_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_8_ldest,io_diffCommits_info_8_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_8_pdest,io_diffCommits_info_8_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_8_rfWen,io_diffCommits_info_8_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_8_fpWen,io_diffCommits_info_8_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_8_vecWen,io_diffCommits_info_8_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_8_v0Wen,io_diffCommits_info_8_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_8_vlWen,io_diffCommits_info_8_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_9_ldest,io_diffCommits_info_9_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_9_pdest,io_diffCommits_info_9_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_9_rfWen,io_diffCommits_info_9_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_9_fpWen,io_diffCommits_info_9_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_9_vecWen,io_diffCommits_info_9_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_9_v0Wen,io_diffCommits_info_9_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_9_vlWen,io_diffCommits_info_9_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_10_ldest,io_diffCommits_info_10_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_10_pdest,io_diffCommits_info_10_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_10_rfWen,io_diffCommits_info_10_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_10_fpWen,io_diffCommits_info_10_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_10_vecWen,io_diffCommits_info_10_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_10_v0Wen,io_diffCommits_info_10_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_10_vlWen,io_diffCommits_info_10_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_11_ldest,io_diffCommits_info_11_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_11_pdest,io_diffCommits_info_11_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_11_rfWen,io_diffCommits_info_11_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_11_fpWen,io_diffCommits_info_11_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_11_vecWen,io_diffCommits_info_11_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_11_v0Wen,io_diffCommits_info_11_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_11_vlWen,io_diffCommits_info_11_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_12_ldest,io_diffCommits_info_12_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_12_pdest,io_diffCommits_info_12_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_12_rfWen,io_diffCommits_info_12_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_12_fpWen,io_diffCommits_info_12_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_12_vecWen,io_diffCommits_info_12_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_12_v0Wen,io_diffCommits_info_12_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_12_vlWen,io_diffCommits_info_12_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_13_ldest,io_diffCommits_info_13_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_13_pdest,io_diffCommits_info_13_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_13_rfWen,io_diffCommits_info_13_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_13_fpWen,io_diffCommits_info_13_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_13_vecWen,io_diffCommits_info_13_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_13_v0Wen,io_diffCommits_info_13_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_13_vlWen,io_diffCommits_info_13_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_14_ldest,io_diffCommits_info_14_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_14_pdest,io_diffCommits_info_14_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_14_rfWen,io_diffCommits_info_14_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_14_fpWen,io_diffCommits_info_14_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_14_vecWen,io_diffCommits_info_14_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_14_v0Wen,io_diffCommits_info_14_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_14_vlWen,io_diffCommits_info_14_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_15_ldest,io_diffCommits_info_15_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_15_pdest,io_diffCommits_info_15_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_15_rfWen,io_diffCommits_info_15_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_15_fpWen,io_diffCommits_info_15_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_15_vecWen,io_diffCommits_info_15_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_15_v0Wen,io_diffCommits_info_15_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_15_vlWen,io_diffCommits_info_15_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_16_ldest,io_diffCommits_info_16_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_16_pdest,io_diffCommits_info_16_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_16_rfWen,io_diffCommits_info_16_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_16_fpWen,io_diffCommits_info_16_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_16_vecWen,io_diffCommits_info_16_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_16_v0Wen,io_diffCommits_info_16_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_16_vlWen,io_diffCommits_info_16_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_17_ldest,io_diffCommits_info_17_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_17_pdest,io_diffCommits_info_17_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_17_rfWen,io_diffCommits_info_17_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_17_fpWen,io_diffCommits_info_17_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_17_vecWen,io_diffCommits_info_17_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_17_v0Wen,io_diffCommits_info_17_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_17_vlWen,io_diffCommits_info_17_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_18_ldest,io_diffCommits_info_18_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_18_pdest,io_diffCommits_info_18_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_18_rfWen,io_diffCommits_info_18_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_18_fpWen,io_diffCommits_info_18_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_18_vecWen,io_diffCommits_info_18_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_18_v0Wen,io_diffCommits_info_18_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_18_vlWen,io_diffCommits_info_18_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_19_ldest,io_diffCommits_info_19_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_19_pdest,io_diffCommits_info_19_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_19_rfWen,io_diffCommits_info_19_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_19_fpWen,io_diffCommits_info_19_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_19_vecWen,io_diffCommits_info_19_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_19_v0Wen,io_diffCommits_info_19_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_19_vlWen,io_diffCommits_info_19_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_20_ldest,io_diffCommits_info_20_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_20_pdest,io_diffCommits_info_20_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_20_rfWen,io_diffCommits_info_20_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_20_fpWen,io_diffCommits_info_20_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_20_vecWen,io_diffCommits_info_20_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_20_v0Wen,io_diffCommits_info_20_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_20_vlWen,io_diffCommits_info_20_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_21_ldest,io_diffCommits_info_21_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_21_pdest,io_diffCommits_info_21_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_21_rfWen,io_diffCommits_info_21_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_21_fpWen,io_diffCommits_info_21_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_21_vecWen,io_diffCommits_info_21_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_21_v0Wen,io_diffCommits_info_21_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_21_vlWen,io_diffCommits_info_21_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_22_ldest,io_diffCommits_info_22_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_22_pdest,io_diffCommits_info_22_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_22_rfWen,io_diffCommits_info_22_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_22_fpWen,io_diffCommits_info_22_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_22_vecWen,io_diffCommits_info_22_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_22_v0Wen,io_diffCommits_info_22_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_22_vlWen,io_diffCommits_info_22_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_23_ldest,io_diffCommits_info_23_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_23_pdest,io_diffCommits_info_23_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_23_rfWen,io_diffCommits_info_23_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_23_fpWen,io_diffCommits_info_23_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_23_vecWen,io_diffCommits_info_23_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_23_v0Wen,io_diffCommits_info_23_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_23_vlWen,io_diffCommits_info_23_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_24_ldest,io_diffCommits_info_24_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_24_pdest,io_diffCommits_info_24_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_24_rfWen,io_diffCommits_info_24_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_24_fpWen,io_diffCommits_info_24_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_24_vecWen,io_diffCommits_info_24_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_24_v0Wen,io_diffCommits_info_24_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_24_vlWen,io_diffCommits_info_24_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_25_ldest,io_diffCommits_info_25_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_25_pdest,io_diffCommits_info_25_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_25_rfWen,io_diffCommits_info_25_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_25_fpWen,io_diffCommits_info_25_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_25_vecWen,io_diffCommits_info_25_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_25_v0Wen,io_diffCommits_info_25_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_25_vlWen,io_diffCommits_info_25_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_26_ldest,io_diffCommits_info_26_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_26_pdest,io_diffCommits_info_26_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_26_rfWen,io_diffCommits_info_26_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_26_fpWen,io_diffCommits_info_26_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_26_vecWen,io_diffCommits_info_26_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_26_v0Wen,io_diffCommits_info_26_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_26_vlWen,io_diffCommits_info_26_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_27_ldest,io_diffCommits_info_27_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_27_pdest,io_diffCommits_info_27_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_27_rfWen,io_diffCommits_info_27_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_27_fpWen,io_diffCommits_info_27_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_27_vecWen,io_diffCommits_info_27_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_27_v0Wen,io_diffCommits_info_27_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_27_vlWen,io_diffCommits_info_27_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_28_ldest,io_diffCommits_info_28_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_28_pdest,io_diffCommits_info_28_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_28_rfWen,io_diffCommits_info_28_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_28_fpWen,io_diffCommits_info_28_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_28_vecWen,io_diffCommits_info_28_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_28_v0Wen,io_diffCommits_info_28_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_28_vlWen,io_diffCommits_info_28_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_29_ldest,io_diffCommits_info_29_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_29_pdest,io_diffCommits_info_29_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_29_rfWen,io_diffCommits_info_29_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_29_fpWen,io_diffCommits_info_29_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_29_vecWen,io_diffCommits_info_29_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_29_v0Wen,io_diffCommits_info_29_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_29_vlWen,io_diffCommits_info_29_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_30_ldest,io_diffCommits_info_30_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_30_pdest,io_diffCommits_info_30_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_30_rfWen,io_diffCommits_info_30_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_30_fpWen,io_diffCommits_info_30_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_30_vecWen,io_diffCommits_info_30_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_30_v0Wen,io_diffCommits_info_30_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_30_vlWen,io_diffCommits_info_30_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_31_ldest,io_diffCommits_info_31_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_31_pdest,io_diffCommits_info_31_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_31_rfWen,io_diffCommits_info_31_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_31_fpWen,io_diffCommits_info_31_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_31_vecWen,io_diffCommits_info_31_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_31_v0Wen,io_diffCommits_info_31_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_31_vlWen,io_diffCommits_info_31_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_32_ldest,io_diffCommits_info_32_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_32_pdest,io_diffCommits_info_32_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_32_rfWen,io_diffCommits_info_32_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_32_fpWen,io_diffCommits_info_32_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_32_vecWen,io_diffCommits_info_32_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_32_v0Wen,io_diffCommits_info_32_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_32_vlWen,io_diffCommits_info_32_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_33_ldest,io_diffCommits_info_33_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_33_pdest,io_diffCommits_info_33_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_33_rfWen,io_diffCommits_info_33_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_33_fpWen,io_diffCommits_info_33_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_33_vecWen,io_diffCommits_info_33_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_33_v0Wen,io_diffCommits_info_33_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_33_vlWen,io_diffCommits_info_33_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_34_ldest,io_diffCommits_info_34_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_34_pdest,io_diffCommits_info_34_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_34_rfWen,io_diffCommits_info_34_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_34_fpWen,io_diffCommits_info_34_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_34_vecWen,io_diffCommits_info_34_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_34_v0Wen,io_diffCommits_info_34_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_34_vlWen,io_diffCommits_info_34_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_35_ldest,io_diffCommits_info_35_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_35_pdest,io_diffCommits_info_35_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_35_rfWen,io_diffCommits_info_35_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_35_fpWen,io_diffCommits_info_35_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_35_vecWen,io_diffCommits_info_35_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_35_v0Wen,io_diffCommits_info_35_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_35_vlWen,io_diffCommits_info_35_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_36_ldest,io_diffCommits_info_36_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_36_pdest,io_diffCommits_info_36_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_36_rfWen,io_diffCommits_info_36_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_36_fpWen,io_diffCommits_info_36_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_36_vecWen,io_diffCommits_info_36_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_36_v0Wen,io_diffCommits_info_36_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_36_vlWen,io_diffCommits_info_36_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_37_ldest,io_diffCommits_info_37_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_37_pdest,io_diffCommits_info_37_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_37_rfWen,io_diffCommits_info_37_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_37_fpWen,io_diffCommits_info_37_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_37_vecWen,io_diffCommits_info_37_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_37_v0Wen,io_diffCommits_info_37_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_37_vlWen,io_diffCommits_info_37_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_38_ldest,io_diffCommits_info_38_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_38_pdest,io_diffCommits_info_38_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_38_rfWen,io_diffCommits_info_38_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_38_fpWen,io_diffCommits_info_38_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_38_vecWen,io_diffCommits_info_38_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_38_v0Wen,io_diffCommits_info_38_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_38_vlWen,io_diffCommits_info_38_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_39_ldest,io_diffCommits_info_39_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_39_pdest,io_diffCommits_info_39_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_39_rfWen,io_diffCommits_info_39_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_39_fpWen,io_diffCommits_info_39_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_39_vecWen,io_diffCommits_info_39_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_39_v0Wen,io_diffCommits_info_39_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_39_vlWen,io_diffCommits_info_39_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_40_ldest,io_diffCommits_info_40_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_40_pdest,io_diffCommits_info_40_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_40_rfWen,io_diffCommits_info_40_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_40_fpWen,io_diffCommits_info_40_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_40_vecWen,io_diffCommits_info_40_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_40_v0Wen,io_diffCommits_info_40_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_40_vlWen,io_diffCommits_info_40_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_41_ldest,io_diffCommits_info_41_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_41_pdest,io_diffCommits_info_41_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_41_rfWen,io_diffCommits_info_41_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_41_fpWen,io_diffCommits_info_41_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_41_vecWen,io_diffCommits_info_41_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_41_v0Wen,io_diffCommits_info_41_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_41_vlWen,io_diffCommits_info_41_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_42_ldest,io_diffCommits_info_42_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_42_pdest,io_diffCommits_info_42_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_42_rfWen,io_diffCommits_info_42_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_42_fpWen,io_diffCommits_info_42_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_42_vecWen,io_diffCommits_info_42_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_42_v0Wen,io_diffCommits_info_42_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_42_vlWen,io_diffCommits_info_42_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_43_ldest,io_diffCommits_info_43_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_43_pdest,io_diffCommits_info_43_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_43_rfWen,io_diffCommits_info_43_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_43_fpWen,io_diffCommits_info_43_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_43_vecWen,io_diffCommits_info_43_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_43_v0Wen,io_diffCommits_info_43_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_43_vlWen,io_diffCommits_info_43_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_44_ldest,io_diffCommits_info_44_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_44_pdest,io_diffCommits_info_44_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_44_rfWen,io_diffCommits_info_44_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_44_fpWen,io_diffCommits_info_44_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_44_vecWen,io_diffCommits_info_44_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_44_v0Wen,io_diffCommits_info_44_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_44_vlWen,io_diffCommits_info_44_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_45_ldest,io_diffCommits_info_45_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_45_pdest,io_diffCommits_info_45_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_45_rfWen,io_diffCommits_info_45_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_45_fpWen,io_diffCommits_info_45_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_45_vecWen,io_diffCommits_info_45_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_45_v0Wen,io_diffCommits_info_45_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_45_vlWen,io_diffCommits_info_45_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_46_ldest,io_diffCommits_info_46_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_46_pdest,io_diffCommits_info_46_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_46_rfWen,io_diffCommits_info_46_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_46_fpWen,io_diffCommits_info_46_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_46_vecWen,io_diffCommits_info_46_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_46_v0Wen,io_diffCommits_info_46_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_46_vlWen,io_diffCommits_info_46_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_47_ldest,io_diffCommits_info_47_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_47_pdest,io_diffCommits_info_47_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_47_rfWen,io_diffCommits_info_47_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_47_fpWen,io_diffCommits_info_47_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_47_vecWen,io_diffCommits_info_47_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_47_v0Wen,io_diffCommits_info_47_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_47_vlWen,io_diffCommits_info_47_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_48_ldest,io_diffCommits_info_48_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_48_pdest,io_diffCommits_info_48_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_48_rfWen,io_diffCommits_info_48_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_48_fpWen,io_diffCommits_info_48_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_48_vecWen,io_diffCommits_info_48_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_48_v0Wen,io_diffCommits_info_48_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_48_vlWen,io_diffCommits_info_48_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_49_ldest,io_diffCommits_info_49_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_49_pdest,io_diffCommits_info_49_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_49_rfWen,io_diffCommits_info_49_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_49_fpWen,io_diffCommits_info_49_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_49_vecWen,io_diffCommits_info_49_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_49_v0Wen,io_diffCommits_info_49_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_49_vlWen,io_diffCommits_info_49_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_50_ldest,io_diffCommits_info_50_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_50_pdest,io_diffCommits_info_50_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_50_rfWen,io_diffCommits_info_50_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_50_fpWen,io_diffCommits_info_50_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_50_vecWen,io_diffCommits_info_50_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_50_v0Wen,io_diffCommits_info_50_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_50_vlWen,io_diffCommits_info_50_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_51_ldest,io_diffCommits_info_51_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_51_pdest,io_diffCommits_info_51_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_51_rfWen,io_diffCommits_info_51_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_51_fpWen,io_diffCommits_info_51_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_51_vecWen,io_diffCommits_info_51_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_51_v0Wen,io_diffCommits_info_51_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_51_vlWen,io_diffCommits_info_51_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_52_ldest,io_diffCommits_info_52_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_52_pdest,io_diffCommits_info_52_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_52_rfWen,io_diffCommits_info_52_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_52_fpWen,io_diffCommits_info_52_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_52_vecWen,io_diffCommits_info_52_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_52_v0Wen,io_diffCommits_info_52_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_52_vlWen,io_diffCommits_info_52_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_53_ldest,io_diffCommits_info_53_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_53_pdest,io_diffCommits_info_53_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_53_rfWen,io_diffCommits_info_53_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_53_fpWen,io_diffCommits_info_53_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_53_vecWen,io_diffCommits_info_53_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_53_v0Wen,io_diffCommits_info_53_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_53_vlWen,io_diffCommits_info_53_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_54_ldest,io_diffCommits_info_54_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_54_pdest,io_diffCommits_info_54_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_54_rfWen,io_diffCommits_info_54_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_54_fpWen,io_diffCommits_info_54_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_54_vecWen,io_diffCommits_info_54_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_54_v0Wen,io_diffCommits_info_54_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_54_vlWen,io_diffCommits_info_54_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_55_ldest,io_diffCommits_info_55_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_55_pdest,io_diffCommits_info_55_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_55_rfWen,io_diffCommits_info_55_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_55_fpWen,io_diffCommits_info_55_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_55_vecWen,io_diffCommits_info_55_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_55_v0Wen,io_diffCommits_info_55_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_55_vlWen,io_diffCommits_info_55_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_56_ldest,io_diffCommits_info_56_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_56_pdest,io_diffCommits_info_56_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_56_rfWen,io_diffCommits_info_56_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_56_fpWen,io_diffCommits_info_56_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_56_vecWen,io_diffCommits_info_56_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_56_v0Wen,io_diffCommits_info_56_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_56_vlWen,io_diffCommits_info_56_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_57_ldest,io_diffCommits_info_57_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_57_pdest,io_diffCommits_info_57_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_57_rfWen,io_diffCommits_info_57_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_57_fpWen,io_diffCommits_info_57_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_57_vecWen,io_diffCommits_info_57_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_57_v0Wen,io_diffCommits_info_57_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_57_vlWen,io_diffCommits_info_57_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_58_ldest,io_diffCommits_info_58_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_58_pdest,io_diffCommits_info_58_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_58_rfWen,io_diffCommits_info_58_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_58_fpWen,io_diffCommits_info_58_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_58_vecWen,io_diffCommits_info_58_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_58_v0Wen,io_diffCommits_info_58_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_58_vlWen,io_diffCommits_info_58_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_59_ldest,io_diffCommits_info_59_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_59_pdest,io_diffCommits_info_59_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_59_rfWen,io_diffCommits_info_59_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_59_fpWen,io_diffCommits_info_59_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_59_vecWen,io_diffCommits_info_59_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_59_v0Wen,io_diffCommits_info_59_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_59_vlWen,io_diffCommits_info_59_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_60_ldest,io_diffCommits_info_60_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_60_pdest,io_diffCommits_info_60_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_60_rfWen,io_diffCommits_info_60_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_60_fpWen,io_diffCommits_info_60_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_60_vecWen,io_diffCommits_info_60_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_60_v0Wen,io_diffCommits_info_60_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_60_vlWen,io_diffCommits_info_60_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_61_ldest,io_diffCommits_info_61_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_61_pdest,io_diffCommits_info_61_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_61_rfWen,io_diffCommits_info_61_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_61_fpWen,io_diffCommits_info_61_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_61_vecWen,io_diffCommits_info_61_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_61_v0Wen,io_diffCommits_info_61_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_61_vlWen,io_diffCommits_info_61_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_62_ldest,io_diffCommits_info_62_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_62_pdest,io_diffCommits_info_62_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_62_rfWen,io_diffCommits_info_62_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_62_fpWen,io_diffCommits_info_62_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_62_vecWen,io_diffCommits_info_62_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_62_v0Wen,io_diffCommits_info_62_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_62_vlWen,io_diffCommits_info_62_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_63_ldest,io_diffCommits_info_63_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_63_pdest,io_diffCommits_info_63_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_63_rfWen,io_diffCommits_info_63_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_63_fpWen,io_diffCommits_info_63_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_63_vecWen,io_diffCommits_info_63_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_63_v0Wen,io_diffCommits_info_63_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_63_vlWen,io_diffCommits_info_63_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_64_ldest,io_diffCommits_info_64_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_64_pdest,io_diffCommits_info_64_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_64_rfWen,io_diffCommits_info_64_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_64_fpWen,io_diffCommits_info_64_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_64_vecWen,io_diffCommits_info_64_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_64_v0Wen,io_diffCommits_info_64_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_64_vlWen,io_diffCommits_info_64_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_65_ldest,io_diffCommits_info_65_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_65_pdest,io_diffCommits_info_65_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_65_rfWen,io_diffCommits_info_65_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_65_fpWen,io_diffCommits_info_65_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_65_vecWen,io_diffCommits_info_65_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_65_v0Wen,io_diffCommits_info_65_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_65_vlWen,io_diffCommits_info_65_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_66_ldest,io_diffCommits_info_66_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_66_pdest,io_diffCommits_info_66_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_66_rfWen,io_diffCommits_info_66_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_66_fpWen,io_diffCommits_info_66_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_66_vecWen,io_diffCommits_info_66_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_66_v0Wen,io_diffCommits_info_66_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_66_vlWen,io_diffCommits_info_66_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_67_ldest,io_diffCommits_info_67_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_67_pdest,io_diffCommits_info_67_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_67_rfWen,io_diffCommits_info_67_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_67_fpWen,io_diffCommits_info_67_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_67_vecWen,io_diffCommits_info_67_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_67_v0Wen,io_diffCommits_info_67_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_67_vlWen,io_diffCommits_info_67_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_68_ldest,io_diffCommits_info_68_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_68_pdest,io_diffCommits_info_68_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_68_rfWen,io_diffCommits_info_68_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_68_fpWen,io_diffCommits_info_68_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_68_vecWen,io_diffCommits_info_68_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_68_v0Wen,io_diffCommits_info_68_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_68_vlWen,io_diffCommits_info_68_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_69_ldest,io_diffCommits_info_69_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_69_pdest,io_diffCommits_info_69_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_69_rfWen,io_diffCommits_info_69_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_69_fpWen,io_diffCommits_info_69_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_69_vecWen,io_diffCommits_info_69_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_69_v0Wen,io_diffCommits_info_69_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_69_vlWen,io_diffCommits_info_69_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_70_ldest,io_diffCommits_info_70_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_70_pdest,io_diffCommits_info_70_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_70_rfWen,io_diffCommits_info_70_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_70_fpWen,io_diffCommits_info_70_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_70_vecWen,io_diffCommits_info_70_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_70_v0Wen,io_diffCommits_info_70_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_70_vlWen,io_diffCommits_info_70_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_71_ldest,io_diffCommits_info_71_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_71_pdest,io_diffCommits_info_71_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_71_rfWen,io_diffCommits_info_71_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_71_fpWen,io_diffCommits_info_71_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_71_vecWen,io_diffCommits_info_71_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_71_v0Wen,io_diffCommits_info_71_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_71_vlWen,io_diffCommits_info_71_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_72_ldest,io_diffCommits_info_72_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_72_pdest,io_diffCommits_info_72_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_72_rfWen,io_diffCommits_info_72_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_72_fpWen,io_diffCommits_info_72_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_72_vecWen,io_diffCommits_info_72_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_72_v0Wen,io_diffCommits_info_72_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_72_vlWen,io_diffCommits_info_72_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_73_ldest,io_diffCommits_info_73_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_73_pdest,io_diffCommits_info_73_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_73_rfWen,io_diffCommits_info_73_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_73_fpWen,io_diffCommits_info_73_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_73_vecWen,io_diffCommits_info_73_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_73_v0Wen,io_diffCommits_info_73_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_73_vlWen,io_diffCommits_info_73_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_74_ldest,io_diffCommits_info_74_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_74_pdest,io_diffCommits_info_74_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_74_rfWen,io_diffCommits_info_74_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_74_fpWen,io_diffCommits_info_74_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_74_vecWen,io_diffCommits_info_74_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_74_v0Wen,io_diffCommits_info_74_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_74_vlWen,io_diffCommits_info_74_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_75_ldest,io_diffCommits_info_75_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_75_pdest,io_diffCommits_info_75_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_75_rfWen,io_diffCommits_info_75_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_75_fpWen,io_diffCommits_info_75_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_75_vecWen,io_diffCommits_info_75_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_75_v0Wen,io_diffCommits_info_75_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_75_vlWen,io_diffCommits_info_75_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_76_ldest,io_diffCommits_info_76_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_76_pdest,io_diffCommits_info_76_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_76_rfWen,io_diffCommits_info_76_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_76_fpWen,io_diffCommits_info_76_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_76_vecWen,io_diffCommits_info_76_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_76_v0Wen,io_diffCommits_info_76_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_76_vlWen,io_diffCommits_info_76_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_77_ldest,io_diffCommits_info_77_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_77_pdest,io_diffCommits_info_77_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_77_rfWen,io_diffCommits_info_77_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_77_fpWen,io_diffCommits_info_77_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_77_vecWen,io_diffCommits_info_77_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_77_v0Wen,io_diffCommits_info_77_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_77_vlWen,io_diffCommits_info_77_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_78_ldest,io_diffCommits_info_78_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_78_pdest,io_diffCommits_info_78_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_78_rfWen,io_diffCommits_info_78_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_78_fpWen,io_diffCommits_info_78_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_78_vecWen,io_diffCommits_info_78_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_78_v0Wen,io_diffCommits_info_78_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_78_vlWen,io_diffCommits_info_78_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_79_ldest,io_diffCommits_info_79_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_79_pdest,io_diffCommits_info_79_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_79_rfWen,io_diffCommits_info_79_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_79_fpWen,io_diffCommits_info_79_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_79_vecWen,io_diffCommits_info_79_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_79_v0Wen,io_diffCommits_info_79_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_79_vlWen,io_diffCommits_info_79_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_80_ldest,io_diffCommits_info_80_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_80_pdest,io_diffCommits_info_80_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_80_rfWen,io_diffCommits_info_80_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_80_fpWen,io_diffCommits_info_80_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_80_vecWen,io_diffCommits_info_80_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_80_v0Wen,io_diffCommits_info_80_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_80_vlWen,io_diffCommits_info_80_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_81_ldest,io_diffCommits_info_81_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_81_pdest,io_diffCommits_info_81_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_81_rfWen,io_diffCommits_info_81_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_81_fpWen,io_diffCommits_info_81_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_81_vecWen,io_diffCommits_info_81_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_81_v0Wen,io_diffCommits_info_81_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_81_vlWen,io_diffCommits_info_81_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_82_ldest,io_diffCommits_info_82_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_82_pdest,io_diffCommits_info_82_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_82_rfWen,io_diffCommits_info_82_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_82_fpWen,io_diffCommits_info_82_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_82_vecWen,io_diffCommits_info_82_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_82_v0Wen,io_diffCommits_info_82_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_82_vlWen,io_diffCommits_info_82_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_83_ldest,io_diffCommits_info_83_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_83_pdest,io_diffCommits_info_83_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_83_rfWen,io_diffCommits_info_83_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_83_fpWen,io_diffCommits_info_83_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_83_vecWen,io_diffCommits_info_83_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_83_v0Wen,io_diffCommits_info_83_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_83_vlWen,io_diffCommits_info_83_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_84_ldest,io_diffCommits_info_84_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_84_pdest,io_diffCommits_info_84_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_84_rfWen,io_diffCommits_info_84_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_84_fpWen,io_diffCommits_info_84_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_84_vecWen,io_diffCommits_info_84_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_84_v0Wen,io_diffCommits_info_84_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_84_vlWen,io_diffCommits_info_84_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_85_ldest,io_diffCommits_info_85_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_85_pdest,io_diffCommits_info_85_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_85_rfWen,io_diffCommits_info_85_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_85_fpWen,io_diffCommits_info_85_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_85_vecWen,io_diffCommits_info_85_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_85_v0Wen,io_diffCommits_info_85_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_85_vlWen,io_diffCommits_info_85_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_86_ldest,io_diffCommits_info_86_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_86_pdest,io_diffCommits_info_86_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_86_rfWen,io_diffCommits_info_86_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_86_fpWen,io_diffCommits_info_86_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_86_vecWen,io_diffCommits_info_86_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_86_v0Wen,io_diffCommits_info_86_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_86_vlWen,io_diffCommits_info_86_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_87_ldest,io_diffCommits_info_87_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_87_pdest,io_diffCommits_info_87_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_87_rfWen,io_diffCommits_info_87_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_87_fpWen,io_diffCommits_info_87_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_87_vecWen,io_diffCommits_info_87_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_87_v0Wen,io_diffCommits_info_87_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_87_vlWen,io_diffCommits_info_87_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_88_ldest,io_diffCommits_info_88_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_88_pdest,io_diffCommits_info_88_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_88_rfWen,io_diffCommits_info_88_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_88_fpWen,io_diffCommits_info_88_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_88_vecWen,io_diffCommits_info_88_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_88_v0Wen,io_diffCommits_info_88_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_88_vlWen,io_diffCommits_info_88_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_89_ldest,io_diffCommits_info_89_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_89_pdest,io_diffCommits_info_89_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_89_rfWen,io_diffCommits_info_89_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_89_fpWen,io_diffCommits_info_89_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_89_vecWen,io_diffCommits_info_89_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_89_v0Wen,io_diffCommits_info_89_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_89_vlWen,io_diffCommits_info_89_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_90_ldest,io_diffCommits_info_90_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_90_pdest,io_diffCommits_info_90_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_90_rfWen,io_diffCommits_info_90_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_90_fpWen,io_diffCommits_info_90_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_90_vecWen,io_diffCommits_info_90_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_90_v0Wen,io_diffCommits_info_90_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_90_vlWen,io_diffCommits_info_90_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_91_ldest,io_diffCommits_info_91_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_91_pdest,io_diffCommits_info_91_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_91_rfWen,io_diffCommits_info_91_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_91_fpWen,io_diffCommits_info_91_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_91_vecWen,io_diffCommits_info_91_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_91_v0Wen,io_diffCommits_info_91_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_91_vlWen,io_diffCommits_info_91_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_92_ldest,io_diffCommits_info_92_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_92_pdest,io_diffCommits_info_92_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_92_rfWen,io_diffCommits_info_92_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_92_fpWen,io_diffCommits_info_92_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_92_vecWen,io_diffCommits_info_92_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_92_v0Wen,io_diffCommits_info_92_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_92_vlWen,io_diffCommits_info_92_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_93_ldest,io_diffCommits_info_93_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_93_pdest,io_diffCommits_info_93_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_93_rfWen,io_diffCommits_info_93_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_93_fpWen,io_diffCommits_info_93_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_93_vecWen,io_diffCommits_info_93_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_93_v0Wen,io_diffCommits_info_93_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_93_vlWen,io_diffCommits_info_93_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_94_ldest,io_diffCommits_info_94_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_94_pdest,io_diffCommits_info_94_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_94_rfWen,io_diffCommits_info_94_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_94_fpWen,io_diffCommits_info_94_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_94_vecWen,io_diffCommits_info_94_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_94_v0Wen,io_diffCommits_info_94_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_94_vlWen,io_diffCommits_info_94_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_95_ldest,io_diffCommits_info_95_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_95_pdest,io_diffCommits_info_95_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_95_rfWen,io_diffCommits_info_95_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_95_fpWen,io_diffCommits_info_95_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_95_vecWen,io_diffCommits_info_95_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_95_v0Wen,io_diffCommits_info_95_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_95_vlWen,io_diffCommits_info_95_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_96_ldest,io_diffCommits_info_96_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_96_pdest,io_diffCommits_info_96_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_96_rfWen,io_diffCommits_info_96_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_96_fpWen,io_diffCommits_info_96_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_96_vecWen,io_diffCommits_info_96_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_96_v0Wen,io_diffCommits_info_96_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_96_vlWen,io_diffCommits_info_96_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_97_ldest,io_diffCommits_info_97_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_97_pdest,io_diffCommits_info_97_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_97_rfWen,io_diffCommits_info_97_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_97_fpWen,io_diffCommits_info_97_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_97_vecWen,io_diffCommits_info_97_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_97_v0Wen,io_diffCommits_info_97_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_97_vlWen,io_diffCommits_info_97_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_98_ldest,io_diffCommits_info_98_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_98_pdest,io_diffCommits_info_98_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_98_rfWen,io_diffCommits_info_98_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_98_fpWen,io_diffCommits_info_98_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_98_vecWen,io_diffCommits_info_98_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_98_v0Wen,io_diffCommits_info_98_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_98_vlWen,io_diffCommits_info_98_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_99_ldest,io_diffCommits_info_99_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_99_pdest,io_diffCommits_info_99_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_99_rfWen,io_diffCommits_info_99_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_99_fpWen,io_diffCommits_info_99_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_99_vecWen,io_diffCommits_info_99_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_99_v0Wen,io_diffCommits_info_99_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_99_vlWen,io_diffCommits_info_99_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_100_ldest,io_diffCommits_info_100_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_100_pdest,io_diffCommits_info_100_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_100_rfWen,io_diffCommits_info_100_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_100_fpWen,io_diffCommits_info_100_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_100_vecWen,io_diffCommits_info_100_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_100_v0Wen,io_diffCommits_info_100_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_100_vlWen,io_diffCommits_info_100_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_101_ldest,io_diffCommits_info_101_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_101_pdest,io_diffCommits_info_101_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_101_rfWen,io_diffCommits_info_101_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_101_fpWen,io_diffCommits_info_101_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_101_vecWen,io_diffCommits_info_101_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_101_v0Wen,io_diffCommits_info_101_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_101_vlWen,io_diffCommits_info_101_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_102_ldest,io_diffCommits_info_102_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_102_pdest,io_diffCommits_info_102_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_102_rfWen,io_diffCommits_info_102_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_102_fpWen,io_diffCommits_info_102_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_102_vecWen,io_diffCommits_info_102_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_102_v0Wen,io_diffCommits_info_102_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_102_vlWen,io_diffCommits_info_102_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_103_ldest,io_diffCommits_info_103_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_103_pdest,io_diffCommits_info_103_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_103_rfWen,io_diffCommits_info_103_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_103_fpWen,io_diffCommits_info_103_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_103_vecWen,io_diffCommits_info_103_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_103_v0Wen,io_diffCommits_info_103_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_103_vlWen,io_diffCommits_info_103_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_104_ldest,io_diffCommits_info_104_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_104_pdest,io_diffCommits_info_104_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_104_rfWen,io_diffCommits_info_104_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_104_fpWen,io_diffCommits_info_104_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_104_vecWen,io_diffCommits_info_104_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_104_v0Wen,io_diffCommits_info_104_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_104_vlWen,io_diffCommits_info_104_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_105_ldest,io_diffCommits_info_105_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_105_pdest,io_diffCommits_info_105_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_105_rfWen,io_diffCommits_info_105_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_105_fpWen,io_diffCommits_info_105_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_105_vecWen,io_diffCommits_info_105_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_105_v0Wen,io_diffCommits_info_105_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_105_vlWen,io_diffCommits_info_105_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_106_ldest,io_diffCommits_info_106_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_106_pdest,io_diffCommits_info_106_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_106_rfWen,io_diffCommits_info_106_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_106_fpWen,io_diffCommits_info_106_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_106_vecWen,io_diffCommits_info_106_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_106_v0Wen,io_diffCommits_info_106_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_106_vlWen,io_diffCommits_info_106_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_107_ldest,io_diffCommits_info_107_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_107_pdest,io_diffCommits_info_107_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_107_rfWen,io_diffCommits_info_107_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_107_fpWen,io_diffCommits_info_107_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_107_vecWen,io_diffCommits_info_107_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_107_v0Wen,io_diffCommits_info_107_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_107_vlWen,io_diffCommits_info_107_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_108_ldest,io_diffCommits_info_108_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_108_pdest,io_diffCommits_info_108_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_108_rfWen,io_diffCommits_info_108_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_108_fpWen,io_diffCommits_info_108_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_108_vecWen,io_diffCommits_info_108_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_108_v0Wen,io_diffCommits_info_108_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_108_vlWen,io_diffCommits_info_108_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_109_ldest,io_diffCommits_info_109_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_109_pdest,io_diffCommits_info_109_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_109_rfWen,io_diffCommits_info_109_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_109_fpWen,io_diffCommits_info_109_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_109_vecWen,io_diffCommits_info_109_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_109_v0Wen,io_diffCommits_info_109_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_109_vlWen,io_diffCommits_info_109_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_110_ldest,io_diffCommits_info_110_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_110_pdest,io_diffCommits_info_110_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_110_rfWen,io_diffCommits_info_110_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_110_fpWen,io_diffCommits_info_110_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_110_vecWen,io_diffCommits_info_110_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_110_v0Wen,io_diffCommits_info_110_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_110_vlWen,io_diffCommits_info_110_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_111_ldest,io_diffCommits_info_111_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_111_pdest,io_diffCommits_info_111_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_111_rfWen,io_diffCommits_info_111_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_111_fpWen,io_diffCommits_info_111_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_111_vecWen,io_diffCommits_info_111_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_111_v0Wen,io_diffCommits_info_111_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_111_vlWen,io_diffCommits_info_111_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_112_ldest,io_diffCommits_info_112_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_112_pdest,io_diffCommits_info_112_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_112_rfWen,io_diffCommits_info_112_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_112_fpWen,io_diffCommits_info_112_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_112_vecWen,io_diffCommits_info_112_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_112_v0Wen,io_diffCommits_info_112_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_112_vlWen,io_diffCommits_info_112_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_113_ldest,io_diffCommits_info_113_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_113_pdest,io_diffCommits_info_113_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_113_rfWen,io_diffCommits_info_113_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_113_fpWen,io_diffCommits_info_113_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_113_vecWen,io_diffCommits_info_113_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_113_v0Wen,io_diffCommits_info_113_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_113_vlWen,io_diffCommits_info_113_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_114_ldest,io_diffCommits_info_114_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_114_pdest,io_diffCommits_info_114_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_114_rfWen,io_diffCommits_info_114_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_114_fpWen,io_diffCommits_info_114_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_114_vecWen,io_diffCommits_info_114_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_114_v0Wen,io_diffCommits_info_114_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_114_vlWen,io_diffCommits_info_114_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_115_ldest,io_diffCommits_info_115_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_115_pdest,io_diffCommits_info_115_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_115_rfWen,io_diffCommits_info_115_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_115_fpWen,io_diffCommits_info_115_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_115_vecWen,io_diffCommits_info_115_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_115_v0Wen,io_diffCommits_info_115_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_115_vlWen,io_diffCommits_info_115_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_116_ldest,io_diffCommits_info_116_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_116_pdest,io_diffCommits_info_116_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_116_rfWen,io_diffCommits_info_116_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_116_fpWen,io_diffCommits_info_116_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_116_vecWen,io_diffCommits_info_116_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_116_v0Wen,io_diffCommits_info_116_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_116_vlWen,io_diffCommits_info_116_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_117_ldest,io_diffCommits_info_117_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_117_pdest,io_diffCommits_info_117_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_117_rfWen,io_diffCommits_info_117_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_117_fpWen,io_diffCommits_info_117_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_117_vecWen,io_diffCommits_info_117_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_117_v0Wen,io_diffCommits_info_117_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_117_vlWen,io_diffCommits_info_117_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_118_ldest,io_diffCommits_info_118_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_118_pdest,io_diffCommits_info_118_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_118_rfWen,io_diffCommits_info_118_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_118_fpWen,io_diffCommits_info_118_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_118_vecWen,io_diffCommits_info_118_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_118_v0Wen,io_diffCommits_info_118_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_118_vlWen,io_diffCommits_info_118_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_119_ldest,io_diffCommits_info_119_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_119_pdest,io_diffCommits_info_119_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_119_rfWen,io_diffCommits_info_119_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_119_fpWen,io_diffCommits_info_119_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_119_vecWen,io_diffCommits_info_119_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_119_v0Wen,io_diffCommits_info_119_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_119_vlWen,io_diffCommits_info_119_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_120_ldest,io_diffCommits_info_120_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_120_pdest,io_diffCommits_info_120_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_120_rfWen,io_diffCommits_info_120_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_120_fpWen,io_diffCommits_info_120_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_120_vecWen,io_diffCommits_info_120_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_120_v0Wen,io_diffCommits_info_120_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_120_vlWen,io_diffCommits_info_120_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_121_ldest,io_diffCommits_info_121_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_121_pdest,io_diffCommits_info_121_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_121_rfWen,io_diffCommits_info_121_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_121_fpWen,io_diffCommits_info_121_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_121_vecWen,io_diffCommits_info_121_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_121_v0Wen,io_diffCommits_info_121_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_121_vlWen,io_diffCommits_info_121_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_122_ldest,io_diffCommits_info_122_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_122_pdest,io_diffCommits_info_122_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_122_rfWen,io_diffCommits_info_122_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_122_fpWen,io_diffCommits_info_122_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_122_vecWen,io_diffCommits_info_122_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_122_v0Wen,io_diffCommits_info_122_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_122_vlWen,io_diffCommits_info_122_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_123_ldest,io_diffCommits_info_123_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_123_pdest,io_diffCommits_info_123_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_123_rfWen,io_diffCommits_info_123_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_123_fpWen,io_diffCommits_info_123_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_123_vecWen,io_diffCommits_info_123_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_123_v0Wen,io_diffCommits_info_123_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_123_vlWen,io_diffCommits_info_123_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_124_ldest,io_diffCommits_info_124_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_124_pdest,io_diffCommits_info_124_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_124_rfWen,io_diffCommits_info_124_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_124_fpWen,io_diffCommits_info_124_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_124_vecWen,io_diffCommits_info_124_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_124_v0Wen,io_diffCommits_info_124_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_124_vlWen,io_diffCommits_info_124_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_125_ldest,io_diffCommits_info_125_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_125_pdest,io_diffCommits_info_125_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_125_rfWen,io_diffCommits_info_125_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_125_fpWen,io_diffCommits_info_125_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_125_vecWen,io_diffCommits_info_125_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_125_v0Wen,io_diffCommits_info_125_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_125_vlWen,io_diffCommits_info_125_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_126_ldest,io_diffCommits_info_126_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_126_pdest,io_diffCommits_info_126_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_126_rfWen,io_diffCommits_info_126_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_126_fpWen,io_diffCommits_info_126_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_126_vecWen,io_diffCommits_info_126_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_126_v0Wen,io_diffCommits_info_126_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_126_vlWen,io_diffCommits_info_126_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_127_ldest,io_diffCommits_info_127_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_127_pdest,io_diffCommits_info_127_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_127_rfWen,io_diffCommits_info_127_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_127_fpWen,io_diffCommits_info_127_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_127_vecWen,io_diffCommits_info_127_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_127_v0Wen,io_diffCommits_info_127_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_127_vlWen,io_diffCommits_info_127_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_128_ldest,io_diffCommits_info_128_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_128_pdest,io_diffCommits_info_128_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_128_rfWen,io_diffCommits_info_128_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_128_fpWen,io_diffCommits_info_128_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_128_vecWen,io_diffCommits_info_128_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_128_v0Wen,io_diffCommits_info_128_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_128_vlWen,io_diffCommits_info_128_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_129_ldest,io_diffCommits_info_129_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_129_pdest,io_diffCommits_info_129_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_129_rfWen,io_diffCommits_info_129_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_129_fpWen,io_diffCommits_info_129_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_129_vecWen,io_diffCommits_info_129_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_129_v0Wen,io_diffCommits_info_129_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_129_vlWen,io_diffCommits_info_129_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_130_ldest,io_diffCommits_info_130_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_130_pdest,io_diffCommits_info_130_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_130_rfWen,io_diffCommits_info_130_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_130_fpWen,io_diffCommits_info_130_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_130_vecWen,io_diffCommits_info_130_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_130_v0Wen,io_diffCommits_info_130_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_130_vlWen,io_diffCommits_info_130_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_131_ldest,io_diffCommits_info_131_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_131_pdest,io_diffCommits_info_131_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_131_rfWen,io_diffCommits_info_131_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_131_fpWen,io_diffCommits_info_131_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_131_vecWen,io_diffCommits_info_131_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_131_v0Wen,io_diffCommits_info_131_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_131_vlWen,io_diffCommits_info_131_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_132_ldest,io_diffCommits_info_132_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_132_pdest,io_diffCommits_info_132_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_132_rfWen,io_diffCommits_info_132_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_132_fpWen,io_diffCommits_info_132_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_132_vecWen,io_diffCommits_info_132_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_132_v0Wen,io_diffCommits_info_132_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_132_vlWen,io_diffCommits_info_132_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_133_ldest,io_diffCommits_info_133_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_133_pdest,io_diffCommits_info_133_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_133_rfWen,io_diffCommits_info_133_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_133_fpWen,io_diffCommits_info_133_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_133_vecWen,io_diffCommits_info_133_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_133_v0Wen,io_diffCommits_info_133_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_133_vlWen,io_diffCommits_info_133_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_134_ldest,io_diffCommits_info_134_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_134_pdest,io_diffCommits_info_134_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_134_rfWen,io_diffCommits_info_134_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_134_fpWen,io_diffCommits_info_134_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_134_vecWen,io_diffCommits_info_134_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_134_v0Wen,io_diffCommits_info_134_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_134_vlWen,io_diffCommits_info_134_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_135_ldest,io_diffCommits_info_135_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_135_pdest,io_diffCommits_info_135_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_135_rfWen,io_diffCommits_info_135_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_135_fpWen,io_diffCommits_info_135_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_135_vecWen,io_diffCommits_info_135_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_135_v0Wen,io_diffCommits_info_135_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_135_vlWen,io_diffCommits_info_135_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_136_ldest,io_diffCommits_info_136_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_136_pdest,io_diffCommits_info_136_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_136_rfWen,io_diffCommits_info_136_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_136_fpWen,io_diffCommits_info_136_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_136_vecWen,io_diffCommits_info_136_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_136_v0Wen,io_diffCommits_info_136_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_136_vlWen,io_diffCommits_info_136_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_137_ldest,io_diffCommits_info_137_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_137_pdest,io_diffCommits_info_137_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_137_rfWen,io_diffCommits_info_137_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_137_fpWen,io_diffCommits_info_137_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_137_vecWen,io_diffCommits_info_137_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_137_v0Wen,io_diffCommits_info_137_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_137_vlWen,io_diffCommits_info_137_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_138_ldest,io_diffCommits_info_138_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_138_pdest,io_diffCommits_info_138_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_138_rfWen,io_diffCommits_info_138_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_138_fpWen,io_diffCommits_info_138_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_138_vecWen,io_diffCommits_info_138_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_138_v0Wen,io_diffCommits_info_138_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_138_vlWen,io_diffCommits_info_138_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_139_ldest,io_diffCommits_info_139_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_139_pdest,io_diffCommits_info_139_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_139_rfWen,io_diffCommits_info_139_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_139_fpWen,io_diffCommits_info_139_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_139_vecWen,io_diffCommits_info_139_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_139_v0Wen,io_diffCommits_info_139_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_139_vlWen,io_diffCommits_info_139_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_140_ldest,io_diffCommits_info_140_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_140_pdest,io_diffCommits_info_140_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_140_rfWen,io_diffCommits_info_140_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_140_fpWen,io_diffCommits_info_140_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_140_vecWen,io_diffCommits_info_140_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_140_v0Wen,io_diffCommits_info_140_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_140_vlWen,io_diffCommits_info_140_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_141_ldest,io_diffCommits_info_141_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_141_pdest,io_diffCommits_info_141_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_141_rfWen,io_diffCommits_info_141_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_141_fpWen,io_diffCommits_info_141_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_141_vecWen,io_diffCommits_info_141_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_141_v0Wen,io_diffCommits_info_141_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_141_vlWen,io_diffCommits_info_141_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_142_ldest,io_diffCommits_info_142_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_142_pdest,io_diffCommits_info_142_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_142_rfWen,io_diffCommits_info_142_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_142_fpWen,io_diffCommits_info_142_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_142_vecWen,io_diffCommits_info_142_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_142_v0Wen,io_diffCommits_info_142_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_142_vlWen,io_diffCommits_info_142_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_143_ldest,io_diffCommits_info_143_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_143_pdest,io_diffCommits_info_143_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_143_rfWen,io_diffCommits_info_143_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_143_fpWen,io_diffCommits_info_143_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_143_vecWen,io_diffCommits_info_143_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_143_v0Wen,io_diffCommits_info_143_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_143_vlWen,io_diffCommits_info_143_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_144_ldest,io_diffCommits_info_144_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_144_pdest,io_diffCommits_info_144_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_144_rfWen,io_diffCommits_info_144_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_144_fpWen,io_diffCommits_info_144_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_144_vecWen,io_diffCommits_info_144_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_144_v0Wen,io_diffCommits_info_144_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_144_vlWen,io_diffCommits_info_144_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_145_ldest,io_diffCommits_info_145_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_145_pdest,io_diffCommits_info_145_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_145_rfWen,io_diffCommits_info_145_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_145_fpWen,io_diffCommits_info_145_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_145_vecWen,io_diffCommits_info_145_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_145_v0Wen,io_diffCommits_info_145_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_145_vlWen,io_diffCommits_info_145_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_146_ldest,io_diffCommits_info_146_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_146_pdest,io_diffCommits_info_146_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_146_rfWen,io_diffCommits_info_146_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_146_fpWen,io_diffCommits_info_146_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_146_vecWen,io_diffCommits_info_146_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_146_v0Wen,io_diffCommits_info_146_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_146_vlWen,io_diffCommits_info_146_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_147_ldest,io_diffCommits_info_147_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_147_pdest,io_diffCommits_info_147_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_147_rfWen,io_diffCommits_info_147_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_147_fpWen,io_diffCommits_info_147_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_147_vecWen,io_diffCommits_info_147_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_147_v0Wen,io_diffCommits_info_147_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_147_vlWen,io_diffCommits_info_147_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_148_ldest,io_diffCommits_info_148_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_148_pdest,io_diffCommits_info_148_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_148_rfWen,io_diffCommits_info_148_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_148_fpWen,io_diffCommits_info_148_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_148_vecWen,io_diffCommits_info_148_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_148_v0Wen,io_diffCommits_info_148_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_148_vlWen,io_diffCommits_info_148_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_149_ldest,io_diffCommits_info_149_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_149_pdest,io_diffCommits_info_149_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_149_rfWen,io_diffCommits_info_149_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_149_fpWen,io_diffCommits_info_149_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_149_vecWen,io_diffCommits_info_149_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_149_v0Wen,io_diffCommits_info_149_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_149_vlWen,io_diffCommits_info_149_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_150_ldest,io_diffCommits_info_150_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_150_pdest,io_diffCommits_info_150_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_150_rfWen,io_diffCommits_info_150_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_150_fpWen,io_diffCommits_info_150_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_150_vecWen,io_diffCommits_info_150_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_150_v0Wen,io_diffCommits_info_150_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_150_vlWen,io_diffCommits_info_150_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_151_ldest,io_diffCommits_info_151_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_151_pdest,io_diffCommits_info_151_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_151_rfWen,io_diffCommits_info_151_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_151_fpWen,io_diffCommits_info_151_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_151_vecWen,io_diffCommits_info_151_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_151_v0Wen,io_diffCommits_info_151_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_151_vlWen,io_diffCommits_info_151_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_152_ldest,io_diffCommits_info_152_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_152_pdest,io_diffCommits_info_152_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_152_rfWen,io_diffCommits_info_152_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_152_fpWen,io_diffCommits_info_152_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_152_vecWen,io_diffCommits_info_152_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_152_v0Wen,io_diffCommits_info_152_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_152_vlWen,io_diffCommits_info_152_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_153_ldest,io_diffCommits_info_153_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_153_pdest,io_diffCommits_info_153_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_153_rfWen,io_diffCommits_info_153_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_153_fpWen,io_diffCommits_info_153_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_153_vecWen,io_diffCommits_info_153_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_153_v0Wen,io_diffCommits_info_153_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_153_vlWen,io_diffCommits_info_153_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_154_ldest,io_diffCommits_info_154_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_154_pdest,io_diffCommits_info_154_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_154_rfWen,io_diffCommits_info_154_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_154_fpWen,io_diffCommits_info_154_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_154_vecWen,io_diffCommits_info_154_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_154_v0Wen,io_diffCommits_info_154_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_154_vlWen,io_diffCommits_info_154_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_155_ldest,io_diffCommits_info_155_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_155_pdest,io_diffCommits_info_155_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_155_rfWen,io_diffCommits_info_155_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_155_fpWen,io_diffCommits_info_155_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_155_vecWen,io_diffCommits_info_155_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_155_v0Wen,io_diffCommits_info_155_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_155_vlWen,io_diffCommits_info_155_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_156_ldest,io_diffCommits_info_156_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_156_pdest,io_diffCommits_info_156_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_156_rfWen,io_diffCommits_info_156_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_156_fpWen,io_diffCommits_info_156_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_156_vecWen,io_diffCommits_info_156_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_156_v0Wen,io_diffCommits_info_156_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_156_vlWen,io_diffCommits_info_156_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_157_ldest,io_diffCommits_info_157_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_157_pdest,io_diffCommits_info_157_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_157_rfWen,io_diffCommits_info_157_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_157_fpWen,io_diffCommits_info_157_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_157_vecWen,io_diffCommits_info_157_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_157_v0Wen,io_diffCommits_info_157_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_157_vlWen,io_diffCommits_info_157_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_158_ldest,io_diffCommits_info_158_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_158_pdest,io_diffCommits_info_158_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_158_rfWen,io_diffCommits_info_158_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_158_fpWen,io_diffCommits_info_158_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_158_vecWen,io_diffCommits_info_158_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_158_v0Wen,io_diffCommits_info_158_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_158_vlWen,io_diffCommits_info_158_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_159_ldest,io_diffCommits_info_159_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_159_pdest,io_diffCommits_info_159_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_159_rfWen,io_diffCommits_info_159_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_159_fpWen,io_diffCommits_info_159_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_159_vecWen,io_diffCommits_info_159_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_159_v0Wen,io_diffCommits_info_159_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_159_vlWen,io_diffCommits_info_159_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_160_ldest,io_diffCommits_info_160_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_160_pdest,io_diffCommits_info_160_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_160_rfWen,io_diffCommits_info_160_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_160_fpWen,io_diffCommits_info_160_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_160_vecWen,io_diffCommits_info_160_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_160_v0Wen,io_diffCommits_info_160_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_160_vlWen,io_diffCommits_info_160_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_161_ldest,io_diffCommits_info_161_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_161_pdest,io_diffCommits_info_161_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_161_rfWen,io_diffCommits_info_161_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_161_fpWen,io_diffCommits_info_161_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_161_vecWen,io_diffCommits_info_161_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_161_v0Wen,io_diffCommits_info_161_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_161_vlWen,io_diffCommits_info_161_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_162_ldest,io_diffCommits_info_162_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_162_pdest,io_diffCommits_info_162_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_162_rfWen,io_diffCommits_info_162_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_162_fpWen,io_diffCommits_info_162_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_162_vecWen,io_diffCommits_info_162_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_162_v0Wen,io_diffCommits_info_162_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_162_vlWen,io_diffCommits_info_162_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_163_ldest,io_diffCommits_info_163_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_163_pdest,io_diffCommits_info_163_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_163_rfWen,io_diffCommits_info_163_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_163_fpWen,io_diffCommits_info_163_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_163_vecWen,io_diffCommits_info_163_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_163_v0Wen,io_diffCommits_info_163_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_163_vlWen,io_diffCommits_info_163_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_164_ldest,io_diffCommits_info_164_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_164_pdest,io_diffCommits_info_164_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_164_rfWen,io_diffCommits_info_164_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_164_fpWen,io_diffCommits_info_164_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_164_vecWen,io_diffCommits_info_164_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_164_v0Wen,io_diffCommits_info_164_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_164_vlWen,io_diffCommits_info_164_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_165_ldest,io_diffCommits_info_165_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_165_pdest,io_diffCommits_info_165_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_165_rfWen,io_diffCommits_info_165_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_165_fpWen,io_diffCommits_info_165_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_165_vecWen,io_diffCommits_info_165_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_165_v0Wen,io_diffCommits_info_165_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_165_vlWen,io_diffCommits_info_165_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_166_ldest,io_diffCommits_info_166_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_166_pdest,io_diffCommits_info_166_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_166_rfWen,io_diffCommits_info_166_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_166_fpWen,io_diffCommits_info_166_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_166_vecWen,io_diffCommits_info_166_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_166_v0Wen,io_diffCommits_info_166_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_166_vlWen,io_diffCommits_info_166_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_167_ldest,io_diffCommits_info_167_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_167_pdest,io_diffCommits_info_167_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_167_rfWen,io_diffCommits_info_167_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_167_fpWen,io_diffCommits_info_167_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_167_vecWen,io_diffCommits_info_167_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_167_v0Wen,io_diffCommits_info_167_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_167_vlWen,io_diffCommits_info_167_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_168_ldest,io_diffCommits_info_168_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_168_pdest,io_diffCommits_info_168_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_168_rfWen,io_diffCommits_info_168_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_168_fpWen,io_diffCommits_info_168_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_168_vecWen,io_diffCommits_info_168_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_168_v0Wen,io_diffCommits_info_168_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_168_vlWen,io_diffCommits_info_168_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_169_ldest,io_diffCommits_info_169_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_169_pdest,io_diffCommits_info_169_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_169_rfWen,io_diffCommits_info_169_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_169_fpWen,io_diffCommits_info_169_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_169_vecWen,io_diffCommits_info_169_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_169_v0Wen,io_diffCommits_info_169_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_169_vlWen,io_diffCommits_info_169_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_170_ldest,io_diffCommits_info_170_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_170_pdest,io_diffCommits_info_170_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_170_rfWen,io_diffCommits_info_170_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_170_fpWen,io_diffCommits_info_170_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_170_vecWen,io_diffCommits_info_170_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_170_v0Wen,io_diffCommits_info_170_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_170_vlWen,io_diffCommits_info_170_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_171_ldest,io_diffCommits_info_171_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_171_pdest,io_diffCommits_info_171_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_171_rfWen,io_diffCommits_info_171_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_171_fpWen,io_diffCommits_info_171_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_171_vecWen,io_diffCommits_info_171_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_171_v0Wen,io_diffCommits_info_171_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_171_vlWen,io_diffCommits_info_171_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_172_ldest,io_diffCommits_info_172_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_172_pdest,io_diffCommits_info_172_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_172_rfWen,io_diffCommits_info_172_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_172_fpWen,io_diffCommits_info_172_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_172_vecWen,io_diffCommits_info_172_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_172_v0Wen,io_diffCommits_info_172_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_172_vlWen,io_diffCommits_info_172_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_173_ldest,io_diffCommits_info_173_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_173_pdest,io_diffCommits_info_173_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_173_rfWen,io_diffCommits_info_173_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_173_fpWen,io_diffCommits_info_173_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_173_vecWen,io_diffCommits_info_173_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_173_v0Wen,io_diffCommits_info_173_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_173_vlWen,io_diffCommits_info_173_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_174_ldest,io_diffCommits_info_174_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_174_pdest,io_diffCommits_info_174_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_174_rfWen,io_diffCommits_info_174_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_174_fpWen,io_diffCommits_info_174_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_174_vecWen,io_diffCommits_info_174_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_174_v0Wen,io_diffCommits_info_174_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_174_vlWen,io_diffCommits_info_174_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_175_ldest,io_diffCommits_info_175_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_175_pdest,io_diffCommits_info_175_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_175_rfWen,io_diffCommits_info_175_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_175_fpWen,io_diffCommits_info_175_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_175_vecWen,io_diffCommits_info_175_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_175_v0Wen,io_diffCommits_info_175_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_175_vlWen,io_diffCommits_info_175_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_176_ldest,io_diffCommits_info_176_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_176_pdest,io_diffCommits_info_176_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_176_rfWen,io_diffCommits_info_176_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_176_fpWen,io_diffCommits_info_176_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_176_vecWen,io_diffCommits_info_176_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_176_v0Wen,io_diffCommits_info_176_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_176_vlWen,io_diffCommits_info_176_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_177_ldest,io_diffCommits_info_177_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_177_pdest,io_diffCommits_info_177_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_177_rfWen,io_diffCommits_info_177_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_177_fpWen,io_diffCommits_info_177_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_177_vecWen,io_diffCommits_info_177_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_177_v0Wen,io_diffCommits_info_177_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_177_vlWen,io_diffCommits_info_177_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_178_ldest,io_diffCommits_info_178_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_178_pdest,io_diffCommits_info_178_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_178_rfWen,io_diffCommits_info_178_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_178_fpWen,io_diffCommits_info_178_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_178_vecWen,io_diffCommits_info_178_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_178_v0Wen,io_diffCommits_info_178_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_178_vlWen,io_diffCommits_info_178_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_179_ldest,io_diffCommits_info_179_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_179_pdest,io_diffCommits_info_179_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_179_rfWen,io_diffCommits_info_179_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_179_fpWen,io_diffCommits_info_179_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_179_vecWen,io_diffCommits_info_179_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_179_v0Wen,io_diffCommits_info_179_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_179_vlWen,io_diffCommits_info_179_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_180_ldest,io_diffCommits_info_180_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_180_pdest,io_diffCommits_info_180_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_180_rfWen,io_diffCommits_info_180_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_180_fpWen,io_diffCommits_info_180_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_180_vecWen,io_diffCommits_info_180_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_180_v0Wen,io_diffCommits_info_180_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_180_vlWen,io_diffCommits_info_180_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_181_ldest,io_diffCommits_info_181_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_181_pdest,io_diffCommits_info_181_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_181_rfWen,io_diffCommits_info_181_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_181_fpWen,io_diffCommits_info_181_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_181_vecWen,io_diffCommits_info_181_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_181_v0Wen,io_diffCommits_info_181_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_181_vlWen,io_diffCommits_info_181_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_182_ldest,io_diffCommits_info_182_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_182_pdest,io_diffCommits_info_182_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_182_rfWen,io_diffCommits_info_182_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_182_fpWen,io_diffCommits_info_182_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_182_vecWen,io_diffCommits_info_182_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_182_v0Wen,io_diffCommits_info_182_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_182_vlWen,io_diffCommits_info_182_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_183_ldest,io_diffCommits_info_183_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_183_pdest,io_diffCommits_info_183_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_183_rfWen,io_diffCommits_info_183_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_183_fpWen,io_diffCommits_info_183_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_183_vecWen,io_diffCommits_info_183_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_183_v0Wen,io_diffCommits_info_183_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_183_vlWen,io_diffCommits_info_183_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_184_ldest,io_diffCommits_info_184_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_184_pdest,io_diffCommits_info_184_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_184_rfWen,io_diffCommits_info_184_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_184_fpWen,io_diffCommits_info_184_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_184_vecWen,io_diffCommits_info_184_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_184_v0Wen,io_diffCommits_info_184_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_184_vlWen,io_diffCommits_info_184_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_185_ldest,io_diffCommits_info_185_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_185_pdest,io_diffCommits_info_185_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_185_rfWen,io_diffCommits_info_185_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_185_fpWen,io_diffCommits_info_185_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_185_vecWen,io_diffCommits_info_185_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_185_v0Wen,io_diffCommits_info_185_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_185_vlWen,io_diffCommits_info_185_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_186_ldest,io_diffCommits_info_186_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_186_pdest,io_diffCommits_info_186_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_186_rfWen,io_diffCommits_info_186_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_186_fpWen,io_diffCommits_info_186_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_186_vecWen,io_diffCommits_info_186_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_186_v0Wen,io_diffCommits_info_186_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_186_vlWen,io_diffCommits_info_186_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_187_ldest,io_diffCommits_info_187_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_187_pdest,io_diffCommits_info_187_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_187_rfWen,io_diffCommits_info_187_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_187_fpWen,io_diffCommits_info_187_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_187_vecWen,io_diffCommits_info_187_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_187_v0Wen,io_diffCommits_info_187_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_187_vlWen,io_diffCommits_info_187_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_188_ldest,io_diffCommits_info_188_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_188_pdest,io_diffCommits_info_188_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_188_rfWen,io_diffCommits_info_188_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_188_fpWen,io_diffCommits_info_188_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_188_vecWen,io_diffCommits_info_188_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_188_v0Wen,io_diffCommits_info_188_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_188_vlWen,io_diffCommits_info_188_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_189_ldest,io_diffCommits_info_189_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_189_pdest,io_diffCommits_info_189_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_189_rfWen,io_diffCommits_info_189_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_189_fpWen,io_diffCommits_info_189_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_189_vecWen,io_diffCommits_info_189_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_189_v0Wen,io_diffCommits_info_189_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_189_vlWen,io_diffCommits_info_189_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_190_ldest,io_diffCommits_info_190_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_190_pdest,io_diffCommits_info_190_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_190_rfWen,io_diffCommits_info_190_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_190_fpWen,io_diffCommits_info_190_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_190_vecWen,io_diffCommits_info_190_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_190_v0Wen,io_diffCommits_info_190_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_190_vlWen,io_diffCommits_info_190_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_191_ldest,io_diffCommits_info_191_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_191_pdest,io_diffCommits_info_191_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_191_rfWen,io_diffCommits_info_191_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_191_fpWen,io_diffCommits_info_191_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_191_vecWen,io_diffCommits_info_191_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_191_v0Wen,io_diffCommits_info_191_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_191_vlWen,io_diffCommits_info_191_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_192_ldest,io_diffCommits_info_192_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_192_pdest,io_diffCommits_info_192_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_192_rfWen,io_diffCommits_info_192_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_192_fpWen,io_diffCommits_info_192_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_192_vecWen,io_diffCommits_info_192_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_192_v0Wen,io_diffCommits_info_192_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_192_vlWen,io_diffCommits_info_192_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_193_ldest,io_diffCommits_info_193_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_193_pdest,io_diffCommits_info_193_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_193_rfWen,io_diffCommits_info_193_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_193_fpWen,io_diffCommits_info_193_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_193_vecWen,io_diffCommits_info_193_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_193_v0Wen,io_diffCommits_info_193_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_193_vlWen,io_diffCommits_info_193_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_194_ldest,io_diffCommits_info_194_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_194_pdest,io_diffCommits_info_194_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_194_rfWen,io_diffCommits_info_194_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_194_fpWen,io_diffCommits_info_194_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_194_vecWen,io_diffCommits_info_194_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_194_v0Wen,io_diffCommits_info_194_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_194_vlWen,io_diffCommits_info_194_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_195_ldest,io_diffCommits_info_195_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_195_pdest,io_diffCommits_info_195_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_195_rfWen,io_diffCommits_info_195_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_195_fpWen,io_diffCommits_info_195_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_195_vecWen,io_diffCommits_info_195_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_195_v0Wen,io_diffCommits_info_195_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_195_vlWen,io_diffCommits_info_195_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_196_ldest,io_diffCommits_info_196_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_196_pdest,io_diffCommits_info_196_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_196_rfWen,io_diffCommits_info_196_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_196_fpWen,io_diffCommits_info_196_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_196_vecWen,io_diffCommits_info_196_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_196_v0Wen,io_diffCommits_info_196_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_196_vlWen,io_diffCommits_info_196_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_197_ldest,io_diffCommits_info_197_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_197_pdest,io_diffCommits_info_197_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_197_rfWen,io_diffCommits_info_197_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_197_fpWen,io_diffCommits_info_197_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_197_vecWen,io_diffCommits_info_197_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_197_v0Wen,io_diffCommits_info_197_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_197_vlWen,io_diffCommits_info_197_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_198_ldest,io_diffCommits_info_198_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_198_pdest,io_diffCommits_info_198_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_198_rfWen,io_diffCommits_info_198_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_198_fpWen,io_diffCommits_info_198_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_198_vecWen,io_diffCommits_info_198_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_198_v0Wen,io_diffCommits_info_198_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_198_vlWen,io_diffCommits_info_198_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_199_ldest,io_diffCommits_info_199_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_199_pdest,io_diffCommits_info_199_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_199_rfWen,io_diffCommits_info_199_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_199_fpWen,io_diffCommits_info_199_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_199_vecWen,io_diffCommits_info_199_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_199_v0Wen,io_diffCommits_info_199_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_199_vlWen,io_diffCommits_info_199_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_200_ldest,io_diffCommits_info_200_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_200_pdest,io_diffCommits_info_200_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_200_rfWen,io_diffCommits_info_200_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_200_fpWen,io_diffCommits_info_200_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_200_vecWen,io_diffCommits_info_200_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_200_v0Wen,io_diffCommits_info_200_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_200_vlWen,io_diffCommits_info_200_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_201_ldest,io_diffCommits_info_201_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_201_pdest,io_diffCommits_info_201_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_201_rfWen,io_diffCommits_info_201_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_201_fpWen,io_diffCommits_info_201_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_201_vecWen,io_diffCommits_info_201_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_201_v0Wen,io_diffCommits_info_201_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_201_vlWen,io_diffCommits_info_201_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_202_ldest,io_diffCommits_info_202_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_202_pdest,io_diffCommits_info_202_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_202_rfWen,io_diffCommits_info_202_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_202_fpWen,io_diffCommits_info_202_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_202_vecWen,io_diffCommits_info_202_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_202_v0Wen,io_diffCommits_info_202_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_202_vlWen,io_diffCommits_info_202_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_203_ldest,io_diffCommits_info_203_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_203_pdest,io_diffCommits_info_203_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_203_rfWen,io_diffCommits_info_203_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_203_fpWen,io_diffCommits_info_203_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_203_vecWen,io_diffCommits_info_203_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_203_v0Wen,io_diffCommits_info_203_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_203_vlWen,io_diffCommits_info_203_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_204_ldest,io_diffCommits_info_204_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_204_pdest,io_diffCommits_info_204_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_204_rfWen,io_diffCommits_info_204_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_204_fpWen,io_diffCommits_info_204_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_204_vecWen,io_diffCommits_info_204_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_204_v0Wen,io_diffCommits_info_204_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_204_vlWen,io_diffCommits_info_204_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_205_ldest,io_diffCommits_info_205_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_205_pdest,io_diffCommits_info_205_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_205_rfWen,io_diffCommits_info_205_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_205_fpWen,io_diffCommits_info_205_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_205_vecWen,io_diffCommits_info_205_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_205_v0Wen,io_diffCommits_info_205_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_205_vlWen,io_diffCommits_info_205_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_206_ldest,io_diffCommits_info_206_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_206_pdest,io_diffCommits_info_206_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_206_rfWen,io_diffCommits_info_206_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_206_fpWen,io_diffCommits_info_206_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_206_vecWen,io_diffCommits_info_206_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_206_v0Wen,io_diffCommits_info_206_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_206_vlWen,io_diffCommits_info_206_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_207_ldest,io_diffCommits_info_207_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_207_pdest,io_diffCommits_info_207_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_207_rfWen,io_diffCommits_info_207_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_207_fpWen,io_diffCommits_info_207_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_207_vecWen,io_diffCommits_info_207_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_207_v0Wen,io_diffCommits_info_207_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_207_vlWen,io_diffCommits_info_207_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_208_ldest,io_diffCommits_info_208_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_208_pdest,io_diffCommits_info_208_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_208_rfWen,io_diffCommits_info_208_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_208_fpWen,io_diffCommits_info_208_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_208_vecWen,io_diffCommits_info_208_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_208_v0Wen,io_diffCommits_info_208_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_208_vlWen,io_diffCommits_info_208_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_209_ldest,io_diffCommits_info_209_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_209_pdest,io_diffCommits_info_209_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_209_rfWen,io_diffCommits_info_209_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_209_fpWen,io_diffCommits_info_209_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_209_vecWen,io_diffCommits_info_209_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_209_v0Wen,io_diffCommits_info_209_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_209_vlWen,io_diffCommits_info_209_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_210_ldest,io_diffCommits_info_210_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_210_pdest,io_diffCommits_info_210_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_210_rfWen,io_diffCommits_info_210_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_210_fpWen,io_diffCommits_info_210_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_210_vecWen,io_diffCommits_info_210_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_210_v0Wen,io_diffCommits_info_210_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_210_vlWen,io_diffCommits_info_210_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_211_ldest,io_diffCommits_info_211_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_211_pdest,io_diffCommits_info_211_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_211_rfWen,io_diffCommits_info_211_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_211_fpWen,io_diffCommits_info_211_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_211_vecWen,io_diffCommits_info_211_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_211_v0Wen,io_diffCommits_info_211_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_211_vlWen,io_diffCommits_info_211_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_212_ldest,io_diffCommits_info_212_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_212_pdest,io_diffCommits_info_212_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_212_rfWen,io_diffCommits_info_212_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_212_fpWen,io_diffCommits_info_212_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_212_vecWen,io_diffCommits_info_212_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_212_v0Wen,io_diffCommits_info_212_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_212_vlWen,io_diffCommits_info_212_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_213_ldest,io_diffCommits_info_213_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_213_pdest,io_diffCommits_info_213_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_213_rfWen,io_diffCommits_info_213_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_213_fpWen,io_diffCommits_info_213_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_213_vecWen,io_diffCommits_info_213_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_213_v0Wen,io_diffCommits_info_213_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_213_vlWen,io_diffCommits_info_213_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_214_ldest,io_diffCommits_info_214_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_214_pdest,io_diffCommits_info_214_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_214_rfWen,io_diffCommits_info_214_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_214_fpWen,io_diffCommits_info_214_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_214_vecWen,io_diffCommits_info_214_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_214_v0Wen,io_diffCommits_info_214_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_214_vlWen,io_diffCommits_info_214_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_215_ldest,io_diffCommits_info_215_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_215_pdest,io_diffCommits_info_215_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_215_rfWen,io_diffCommits_info_215_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_215_fpWen,io_diffCommits_info_215_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_215_vecWen,io_diffCommits_info_215_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_215_v0Wen,io_diffCommits_info_215_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_215_vlWen,io_diffCommits_info_215_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_216_ldest,io_diffCommits_info_216_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_216_pdest,io_diffCommits_info_216_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_216_rfWen,io_diffCommits_info_216_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_216_fpWen,io_diffCommits_info_216_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_216_vecWen,io_diffCommits_info_216_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_216_v0Wen,io_diffCommits_info_216_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_216_vlWen,io_diffCommits_info_216_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_217_ldest,io_diffCommits_info_217_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_217_pdest,io_diffCommits_info_217_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_217_rfWen,io_diffCommits_info_217_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_217_fpWen,io_diffCommits_info_217_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_217_vecWen,io_diffCommits_info_217_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_217_v0Wen,io_diffCommits_info_217_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_217_vlWen,io_diffCommits_info_217_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_218_ldest,io_diffCommits_info_218_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_218_pdest,io_diffCommits_info_218_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_218_rfWen,io_diffCommits_info_218_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_218_fpWen,io_diffCommits_info_218_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_218_vecWen,io_diffCommits_info_218_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_218_v0Wen,io_diffCommits_info_218_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_218_vlWen,io_diffCommits_info_218_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_219_ldest,io_diffCommits_info_219_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_219_pdest,io_diffCommits_info_219_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_219_rfWen,io_diffCommits_info_219_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_219_fpWen,io_diffCommits_info_219_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_219_vecWen,io_diffCommits_info_219_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_219_v0Wen,io_diffCommits_info_219_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_219_vlWen,io_diffCommits_info_219_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_220_ldest,io_diffCommits_info_220_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_220_pdest,io_diffCommits_info_220_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_220_rfWen,io_diffCommits_info_220_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_220_fpWen,io_diffCommits_info_220_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_220_vecWen,io_diffCommits_info_220_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_220_v0Wen,io_diffCommits_info_220_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_220_vlWen,io_diffCommits_info_220_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_221_ldest,io_diffCommits_info_221_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_221_pdest,io_diffCommits_info_221_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_221_rfWen,io_diffCommits_info_221_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_221_fpWen,io_diffCommits_info_221_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_221_vecWen,io_diffCommits_info_221_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_221_v0Wen,io_diffCommits_info_221_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_221_vlWen,io_diffCommits_info_221_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_222_ldest,io_diffCommits_info_222_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_222_pdest,io_diffCommits_info_222_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_222_rfWen,io_diffCommits_info_222_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_222_fpWen,io_diffCommits_info_222_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_222_vecWen,io_diffCommits_info_222_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_222_v0Wen,io_diffCommits_info_222_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_222_vlWen,io_diffCommits_info_222_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_223_ldest,io_diffCommits_info_223_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_223_pdest,io_diffCommits_info_223_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_223_rfWen,io_diffCommits_info_223_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_223_fpWen,io_diffCommits_info_223_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_223_vecWen,io_diffCommits_info_223_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_223_v0Wen,io_diffCommits_info_223_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_223_vlWen,io_diffCommits_info_223_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_224_ldest,io_diffCommits_info_224_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_224_pdest,io_diffCommits_info_224_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_224_rfWen,io_diffCommits_info_224_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_224_fpWen,io_diffCommits_info_224_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_224_vecWen,io_diffCommits_info_224_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_224_v0Wen,io_diffCommits_info_224_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_224_vlWen,io_diffCommits_info_224_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_225_ldest,io_diffCommits_info_225_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_225_pdest,io_diffCommits_info_225_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_225_rfWen,io_diffCommits_info_225_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_225_fpWen,io_diffCommits_info_225_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_225_vecWen,io_diffCommits_info_225_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_225_v0Wen,io_diffCommits_info_225_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_225_vlWen,io_diffCommits_info_225_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_226_ldest,io_diffCommits_info_226_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_226_pdest,io_diffCommits_info_226_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_226_rfWen,io_diffCommits_info_226_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_226_fpWen,io_diffCommits_info_226_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_226_vecWen,io_diffCommits_info_226_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_226_v0Wen,io_diffCommits_info_226_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_226_vlWen,io_diffCommits_info_226_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_227_ldest,io_diffCommits_info_227_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_227_pdest,io_diffCommits_info_227_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_227_rfWen,io_diffCommits_info_227_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_227_fpWen,io_diffCommits_info_227_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_227_vecWen,io_diffCommits_info_227_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_227_v0Wen,io_diffCommits_info_227_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_227_vlWen,io_diffCommits_info_227_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_228_ldest,io_diffCommits_info_228_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_228_pdest,io_diffCommits_info_228_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_228_rfWen,io_diffCommits_info_228_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_228_fpWen,io_diffCommits_info_228_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_228_vecWen,io_diffCommits_info_228_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_228_v0Wen,io_diffCommits_info_228_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_228_vlWen,io_diffCommits_info_228_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_229_ldest,io_diffCommits_info_229_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_229_pdest,io_diffCommits_info_229_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_229_rfWen,io_diffCommits_info_229_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_229_fpWen,io_diffCommits_info_229_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_229_vecWen,io_diffCommits_info_229_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_229_v0Wen,io_diffCommits_info_229_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_229_vlWen,io_diffCommits_info_229_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_230_ldest,io_diffCommits_info_230_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_230_pdest,io_diffCommits_info_230_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_230_rfWen,io_diffCommits_info_230_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_230_fpWen,io_diffCommits_info_230_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_230_vecWen,io_diffCommits_info_230_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_230_v0Wen,io_diffCommits_info_230_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_230_vlWen,io_diffCommits_info_230_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_231_ldest,io_diffCommits_info_231_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_231_pdest,io_diffCommits_info_231_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_231_rfWen,io_diffCommits_info_231_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_231_fpWen,io_diffCommits_info_231_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_231_vecWen,io_diffCommits_info_231_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_231_v0Wen,io_diffCommits_info_231_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_231_vlWen,io_diffCommits_info_231_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_232_ldest,io_diffCommits_info_232_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_232_pdest,io_diffCommits_info_232_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_232_rfWen,io_diffCommits_info_232_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_232_fpWen,io_diffCommits_info_232_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_232_vecWen,io_diffCommits_info_232_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_232_v0Wen,io_diffCommits_info_232_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_232_vlWen,io_diffCommits_info_232_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_233_ldest,io_diffCommits_info_233_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_233_pdest,io_diffCommits_info_233_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_233_rfWen,io_diffCommits_info_233_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_233_fpWen,io_diffCommits_info_233_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_233_vecWen,io_diffCommits_info_233_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_233_v0Wen,io_diffCommits_info_233_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_233_vlWen,io_diffCommits_info_233_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_234_ldest,io_diffCommits_info_234_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_234_pdest,io_diffCommits_info_234_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_234_rfWen,io_diffCommits_info_234_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_234_fpWen,io_diffCommits_info_234_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_234_vecWen,io_diffCommits_info_234_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_234_v0Wen,io_diffCommits_info_234_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_234_vlWen,io_diffCommits_info_234_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_235_ldest,io_diffCommits_info_235_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_235_pdest,io_diffCommits_info_235_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_235_rfWen,io_diffCommits_info_235_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_235_fpWen,io_diffCommits_info_235_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_235_vecWen,io_diffCommits_info_235_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_235_v0Wen,io_diffCommits_info_235_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_235_vlWen,io_diffCommits_info_235_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_236_ldest,io_diffCommits_info_236_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_236_pdest,io_diffCommits_info_236_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_236_rfWen,io_diffCommits_info_236_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_236_fpWen,io_diffCommits_info_236_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_236_vecWen,io_diffCommits_info_236_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_236_v0Wen,io_diffCommits_info_236_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_236_vlWen,io_diffCommits_info_236_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_237_ldest,io_diffCommits_info_237_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_237_pdest,io_diffCommits_info_237_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_237_rfWen,io_diffCommits_info_237_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_237_fpWen,io_diffCommits_info_237_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_237_vecWen,io_diffCommits_info_237_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_237_v0Wen,io_diffCommits_info_237_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_237_vlWen,io_diffCommits_info_237_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_238_ldest,io_diffCommits_info_238_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_238_pdest,io_diffCommits_info_238_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_238_rfWen,io_diffCommits_info_238_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_238_fpWen,io_diffCommits_info_238_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_238_vecWen,io_diffCommits_info_238_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_238_v0Wen,io_diffCommits_info_238_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_238_vlWen,io_diffCommits_info_238_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_239_ldest,io_diffCommits_info_239_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_239_pdest,io_diffCommits_info_239_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_239_rfWen,io_diffCommits_info_239_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_239_fpWen,io_diffCommits_info_239_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_239_vecWen,io_diffCommits_info_239_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_239_v0Wen,io_diffCommits_info_239_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_239_vlWen,io_diffCommits_info_239_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_240_ldest,io_diffCommits_info_240_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_240_pdest,io_diffCommits_info_240_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_240_rfWen,io_diffCommits_info_240_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_240_fpWen,io_diffCommits_info_240_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_240_vecWen,io_diffCommits_info_240_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_240_v0Wen,io_diffCommits_info_240_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_240_vlWen,io_diffCommits_info_240_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_241_ldest,io_diffCommits_info_241_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_241_pdest,io_diffCommits_info_241_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_241_rfWen,io_diffCommits_info_241_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_241_fpWen,io_diffCommits_info_241_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_241_vecWen,io_diffCommits_info_241_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_241_v0Wen,io_diffCommits_info_241_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_241_vlWen,io_diffCommits_info_241_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_242_ldest,io_diffCommits_info_242_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_242_pdest,io_diffCommits_info_242_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_242_rfWen,io_diffCommits_info_242_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_242_fpWen,io_diffCommits_info_242_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_242_vecWen,io_diffCommits_info_242_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_242_v0Wen,io_diffCommits_info_242_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_242_vlWen,io_diffCommits_info_242_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_243_ldest,io_diffCommits_info_243_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_243_pdest,io_diffCommits_info_243_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_243_rfWen,io_diffCommits_info_243_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_243_fpWen,io_diffCommits_info_243_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_243_vecWen,io_diffCommits_info_243_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_243_v0Wen,io_diffCommits_info_243_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_243_vlWen,io_diffCommits_info_243_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_244_ldest,io_diffCommits_info_244_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_244_pdest,io_diffCommits_info_244_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_244_rfWen,io_diffCommits_info_244_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_244_fpWen,io_diffCommits_info_244_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_244_vecWen,io_diffCommits_info_244_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_244_v0Wen,io_diffCommits_info_244_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_244_vlWen,io_diffCommits_info_244_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_245_ldest,io_diffCommits_info_245_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_245_pdest,io_diffCommits_info_245_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_245_rfWen,io_diffCommits_info_245_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_245_fpWen,io_diffCommits_info_245_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_245_vecWen,io_diffCommits_info_245_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_245_v0Wen,io_diffCommits_info_245_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_245_vlWen,io_diffCommits_info_245_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_246_ldest,io_diffCommits_info_246_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_246_pdest,io_diffCommits_info_246_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_246_rfWen,io_diffCommits_info_246_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_246_fpWen,io_diffCommits_info_246_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_246_vecWen,io_diffCommits_info_246_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_246_v0Wen,io_diffCommits_info_246_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_246_vlWen,io_diffCommits_info_246_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_247_ldest,io_diffCommits_info_247_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_247_pdest,io_diffCommits_info_247_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_247_rfWen,io_diffCommits_info_247_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_247_fpWen,io_diffCommits_info_247_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_247_vecWen,io_diffCommits_info_247_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_247_v0Wen,io_diffCommits_info_247_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_247_vlWen,io_diffCommits_info_247_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_248_ldest,io_diffCommits_info_248_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_248_pdest,io_diffCommits_info_248_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_248_rfWen,io_diffCommits_info_248_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_248_fpWen,io_diffCommits_info_248_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_248_vecWen,io_diffCommits_info_248_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_248_v0Wen,io_diffCommits_info_248_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_248_vlWen,io_diffCommits_info_248_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_249_ldest,io_diffCommits_info_249_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_249_pdest,io_diffCommits_info_249_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_249_rfWen,io_diffCommits_info_249_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_249_fpWen,io_diffCommits_info_249_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_249_vecWen,io_diffCommits_info_249_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_249_v0Wen,io_diffCommits_info_249_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_249_vlWen,io_diffCommits_info_249_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_250_ldest,io_diffCommits_info_250_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_250_pdest,io_diffCommits_info_250_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_250_rfWen,io_diffCommits_info_250_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_250_fpWen,io_diffCommits_info_250_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_250_vecWen,io_diffCommits_info_250_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_250_v0Wen,io_diffCommits_info_250_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_250_vlWen,io_diffCommits_info_250_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_251_ldest,io_diffCommits_info_251_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_251_pdest,io_diffCommits_info_251_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_251_rfWen,io_diffCommits_info_251_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_251_fpWen,io_diffCommits_info_251_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_251_vecWen,io_diffCommits_info_251_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_251_v0Wen,io_diffCommits_info_251_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_251_vlWen,io_diffCommits_info_251_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_252_ldest,io_diffCommits_info_252_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_252_pdest,io_diffCommits_info_252_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_252_rfWen,io_diffCommits_info_252_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_252_fpWen,io_diffCommits_info_252_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_252_vecWen,io_diffCommits_info_252_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_252_v0Wen,io_diffCommits_info_252_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_252_vlWen,io_diffCommits_info_252_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_253_ldest,io_diffCommits_info_253_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_253_pdest,io_diffCommits_info_253_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_253_rfWen,io_diffCommits_info_253_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_253_fpWen,io_diffCommits_info_253_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_253_vecWen,io_diffCommits_info_253_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_253_v0Wen,io_diffCommits_info_253_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_253_vlWen,io_diffCommits_info_253_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_254_ldest,io_diffCommits_info_254_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_254_pdest,io_diffCommits_info_254_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_254_rfWen,io_diffCommits_info_254_rfWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_254_fpWen,io_diffCommits_info_254_fpWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_254_vecWen,io_diffCommits_info_254_vecWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_254_v0Wen,io_diffCommits_info_254_v0Wen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_254_vlWen,io_diffCommits_info_254_vlWen,1);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_255_ldest,io_diffCommits_info_255_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_255_pdest,io_diffCommits_info_255_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_256_ldest,io_diffCommits_info_256_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_256_pdest,io_diffCommits_info_256_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_257_ldest,io_diffCommits_info_257_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_257_pdest,io_diffCommits_info_257_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_258_ldest,io_diffCommits_info_258_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_258_pdest,io_diffCommits_info_258_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_259_ldest,io_diffCommits_info_259_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_259_pdest,io_diffCommits_info_259_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_260_ldest,io_diffCommits_info_260_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_260_pdest,io_diffCommits_info_260_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_261_ldest,io_diffCommits_info_261_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_261_pdest,io_diffCommits_info_261_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_262_ldest,io_diffCommits_info_262_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_262_pdest,io_diffCommits_info_262_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_263_ldest,io_diffCommits_info_263_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_263_pdest,io_diffCommits_info_263_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_264_ldest,io_diffCommits_info_264_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_264_pdest,io_diffCommits_info_264_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_265_ldest,io_diffCommits_info_265_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_265_pdest,io_diffCommits_info_265_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_266_ldest,io_diffCommits_info_266_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_266_pdest,io_diffCommits_info_266_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_267_ldest,io_diffCommits_info_267_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_267_pdest,io_diffCommits_info_267_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_268_ldest,io_diffCommits_info_268_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_268_pdest,io_diffCommits_info_268_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_269_ldest,io_diffCommits_info_269_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_269_pdest,io_diffCommits_info_269_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_270_ldest,io_diffCommits_info_270_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_270_pdest,io_diffCommits_info_270_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_271_ldest,io_diffCommits_info_271_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_271_pdest,io_diffCommits_info_271_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_272_ldest,io_diffCommits_info_272_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_272_pdest,io_diffCommits_info_272_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_273_ldest,io_diffCommits_info_273_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_273_pdest,io_diffCommits_info_273_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_274_ldest,io_diffCommits_info_274_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_274_pdest,io_diffCommits_info_274_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_275_ldest,io_diffCommits_info_275_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_275_pdest,io_diffCommits_info_275_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_276_ldest,io_diffCommits_info_276_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_276_pdest,io_diffCommits_info_276_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_277_ldest,io_diffCommits_info_277_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_277_pdest,io_diffCommits_info_277_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_278_ldest,io_diffCommits_info_278_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_278_pdest,io_diffCommits_info_278_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_279_ldest,io_diffCommits_info_279_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_279_pdest,io_diffCommits_info_279_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_280_ldest,io_diffCommits_info_280_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_280_pdest,io_diffCommits_info_280_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_281_ldest,io_diffCommits_info_281_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_281_pdest,io_diffCommits_info_281_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_282_ldest,io_diffCommits_info_282_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_282_pdest,io_diffCommits_info_282_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_283_ldest,io_diffCommits_info_283_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_283_pdest,io_diffCommits_info_283_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_284_ldest,io_diffCommits_info_284_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_284_pdest,io_diffCommits_info_284_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_285_ldest,io_diffCommits_info_285_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_285_pdest,io_diffCommits_info_285_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_286_ldest,io_diffCommits_info_286_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_286_pdest,io_diffCommits_info_286_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_287_ldest,io_diffCommits_info_287_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_287_pdest,io_diffCommits_info_287_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_288_ldest,io_diffCommits_info_288_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_288_pdest,io_diffCommits_info_288_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_289_ldest,io_diffCommits_info_289_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_289_pdest,io_diffCommits_info_289_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_290_ldest,io_diffCommits_info_290_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_290_pdest,io_diffCommits_info_290_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_291_ldest,io_diffCommits_info_291_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_291_pdest,io_diffCommits_info_291_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_292_ldest,io_diffCommits_info_292_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_292_pdest,io_diffCommits_info_292_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_293_ldest,io_diffCommits_info_293_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_293_pdest,io_diffCommits_info_293_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_294_ldest,io_diffCommits_info_294_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_294_pdest,io_diffCommits_info_294_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_295_ldest,io_diffCommits_info_295_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_295_pdest,io_diffCommits_info_295_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_296_ldest,io_diffCommits_info_296_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_296_pdest,io_diffCommits_info_296_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_297_ldest,io_diffCommits_info_297_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_297_pdest,io_diffCommits_info_297_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_298_ldest,io_diffCommits_info_298_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_298_pdest,io_diffCommits_info_298_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_299_ldest,io_diffCommits_info_299_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_299_pdest,io_diffCommits_info_299_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_300_ldest,io_diffCommits_info_300_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_300_pdest,io_diffCommits_info_300_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_301_ldest,io_diffCommits_info_301_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_301_pdest,io_diffCommits_info_301_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_302_ldest,io_diffCommits_info_302_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_302_pdest,io_diffCommits_info_302_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_303_ldest,io_diffCommits_info_303_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_303_pdest,io_diffCommits_info_303_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_304_ldest,io_diffCommits_info_304_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_304_pdest,io_diffCommits_info_304_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_305_ldest,io_diffCommits_info_305_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_305_pdest,io_diffCommits_info_305_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_306_ldest,io_diffCommits_info_306_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_306_pdest,io_diffCommits_info_306_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_307_ldest,io_diffCommits_info_307_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_307_pdest,io_diffCommits_info_307_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_308_ldest,io_diffCommits_info_308_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_308_pdest,io_diffCommits_info_308_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_309_ldest,io_diffCommits_info_309_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_309_pdest,io_diffCommits_info_309_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_310_ldest,io_diffCommits_info_310_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_310_pdest,io_diffCommits_info_310_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_311_ldest,io_diffCommits_info_311_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_311_pdest,io_diffCommits_info_311_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_312_ldest,io_diffCommits_info_312_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_312_pdest,io_diffCommits_info_312_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_313_ldest,io_diffCommits_info_313_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_313_pdest,io_diffCommits_info_313_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_314_ldest,io_diffCommits_info_314_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_314_pdest,io_diffCommits_info_314_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_315_ldest,io_diffCommits_info_315_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_315_pdest,io_diffCommits_info_315_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_316_ldest,io_diffCommits_info_316_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_316_pdest,io_diffCommits_info_316_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_317_ldest,io_diffCommits_info_317_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_317_pdest,io_diffCommits_info_317_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_318_ldest,io_diffCommits_info_318_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_318_pdest,io_diffCommits_info_318_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_319_ldest,io_diffCommits_info_319_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_319_pdest,io_diffCommits_info_319_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_320_ldest,io_diffCommits_info_320_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_320_pdest,io_diffCommits_info_320_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_321_ldest,io_diffCommits_info_321_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_321_pdest,io_diffCommits_info_321_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_322_ldest,io_diffCommits_info_322_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_322_pdest,io_diffCommits_info_322_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_323_ldest,io_diffCommits_info_323_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_323_pdest,io_diffCommits_info_323_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_324_ldest,io_diffCommits_info_324_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_324_pdest,io_diffCommits_info_324_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_325_ldest,io_diffCommits_info_325_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_325_pdest,io_diffCommits_info_325_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_326_ldest,io_diffCommits_info_326_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_326_pdest,io_diffCommits_info_326_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_327_ldest,io_diffCommits_info_327_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_327_pdest,io_diffCommits_info_327_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_328_ldest,io_diffCommits_info_328_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_328_pdest,io_diffCommits_info_328_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_329_ldest,io_diffCommits_info_329_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_329_pdest,io_diffCommits_info_329_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_330_ldest,io_diffCommits_info_330_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_330_pdest,io_diffCommits_info_330_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_331_ldest,io_diffCommits_info_331_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_331_pdest,io_diffCommits_info_331_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_332_ldest,io_diffCommits_info_332_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_332_pdest,io_diffCommits_info_332_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_333_ldest,io_diffCommits_info_333_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_333_pdest,io_diffCommits_info_333_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_334_ldest,io_diffCommits_info_334_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_334_pdest,io_diffCommits_info_334_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_335_ldest,io_diffCommits_info_335_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_335_pdest,io_diffCommits_info_335_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_336_ldest,io_diffCommits_info_336_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_336_pdest,io_diffCommits_info_336_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_337_ldest,io_diffCommits_info_337_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_337_pdest,io_diffCommits_info_337_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_338_ldest,io_diffCommits_info_338_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_338_pdest,io_diffCommits_info_338_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_339_ldest,io_diffCommits_info_339_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_339_pdest,io_diffCommits_info_339_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_340_ldest,io_diffCommits_info_340_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_340_pdest,io_diffCommits_info_340_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_341_ldest,io_diffCommits_info_341_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_341_pdest,io_diffCommits_info_341_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_342_ldest,io_diffCommits_info_342_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_342_pdest,io_diffCommits_info_342_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_343_ldest,io_diffCommits_info_343_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_343_pdest,io_diffCommits_info_343_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_344_ldest,io_diffCommits_info_344_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_344_pdest,io_diffCommits_info_344_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_345_ldest,io_diffCommits_info_345_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_345_pdest,io_diffCommits_info_345_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_346_ldest,io_diffCommits_info_346_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_346_pdest,io_diffCommits_info_346_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_347_ldest,io_diffCommits_info_347_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_347_pdest,io_diffCommits_info_347_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_348_ldest,io_diffCommits_info_348_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_348_pdest,io_diffCommits_info_348_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_349_ldest,io_diffCommits_info_349_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_349_pdest,io_diffCommits_info_349_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_350_ldest,io_diffCommits_info_350_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_350_pdest,io_diffCommits_info_350_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_351_ldest,io_diffCommits_info_351_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_351_pdest,io_diffCommits_info_351_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_352_ldest,io_diffCommits_info_352_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_352_pdest,io_diffCommits_info_352_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_353_ldest,io_diffCommits_info_353_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_353_pdest,io_diffCommits_info_353_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_354_ldest,io_diffCommits_info_354_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_354_pdest,io_diffCommits_info_354_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_355_ldest,io_diffCommits_info_355_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_355_pdest,io_diffCommits_info_355_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_356_ldest,io_diffCommits_info_356_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_356_pdest,io_diffCommits_info_356_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_357_ldest,io_diffCommits_info_357_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_357_pdest,io_diffCommits_info_357_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_358_ldest,io_diffCommits_info_358_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_358_pdest,io_diffCommits_info_358_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_359_ldest,io_diffCommits_info_359_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_359_pdest,io_diffCommits_info_359_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_360_ldest,io_diffCommits_info_360_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_360_pdest,io_diffCommits_info_360_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_361_ldest,io_diffCommits_info_361_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_361_pdest,io_diffCommits_info_361_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_362_ldest,io_diffCommits_info_362_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_362_pdest,io_diffCommits_info_362_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_363_ldest,io_diffCommits_info_363_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_363_pdest,io_diffCommits_info_363_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_364_ldest,io_diffCommits_info_364_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_364_pdest,io_diffCommits_info_364_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_365_ldest,io_diffCommits_info_365_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_365_pdest,io_diffCommits_info_365_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_366_ldest,io_diffCommits_info_366_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_366_pdest,io_diffCommits_info_366_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_367_ldest,io_diffCommits_info_367_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_367_pdest,io_diffCommits_info_367_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_368_ldest,io_diffCommits_info_368_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_368_pdest,io_diffCommits_info_368_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_369_ldest,io_diffCommits_info_369_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_369_pdest,io_diffCommits_info_369_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_370_ldest,io_diffCommits_info_370_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_370_pdest,io_diffCommits_info_370_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_371_ldest,io_diffCommits_info_371_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_371_pdest,io_diffCommits_info_371_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_372_ldest,io_diffCommits_info_372_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_372_pdest,io_diffCommits_info_372_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_373_ldest,io_diffCommits_info_373_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_373_pdest,io_diffCommits_info_373_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_374_ldest,io_diffCommits_info_374_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_374_pdest,io_diffCommits_info_374_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_375_ldest,io_diffCommits_info_375_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_375_pdest,io_diffCommits_info_375_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_376_ldest,io_diffCommits_info_376_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_376_pdest,io_diffCommits_info_376_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_377_ldest,io_diffCommits_info_377_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_377_pdest,io_diffCommits_info_377_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_378_ldest,io_diffCommits_info_378_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_378_pdest,io_diffCommits_info_378_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_379_ldest,io_diffCommits_info_379_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_379_pdest,io_diffCommits_info_379_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_380_ldest,io_diffCommits_info_380_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_380_pdest,io_diffCommits_info_380_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_381_ldest,io_diffCommits_info_381_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_381_pdest,io_diffCommits_info_381_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_382_ldest,io_diffCommits_info_382_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_382_pdest,io_diffCommits_info_382_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_383_ldest,io_diffCommits_info_383_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_383_pdest,io_diffCommits_info_383_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_384_ldest,io_diffCommits_info_384_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_384_pdest,io_diffCommits_info_384_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_385_ldest,io_diffCommits_info_385_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_385_pdest,io_diffCommits_info_385_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_386_ldest,io_diffCommits_info_386_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_386_pdest,io_diffCommits_info_386_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_387_ldest,io_diffCommits_info_387_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_387_pdest,io_diffCommits_info_387_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_388_ldest,io_diffCommits_info_388_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_388_pdest,io_diffCommits_info_388_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_389_ldest,io_diffCommits_info_389_ldest,6);
        //     `TCNT_CHECK_SIG_XZ(io_diffCommits_info_389_pdest,io_diffCommits_info_389_pdest,8);
        //     `TCNT_CHECK_SIG_XZ(io_lsq_scommit,io_lsq_scommit,4);
        //     `TCNT_CHECK_SIG_XZ(io_lsq_pendingMMIOld,io_lsq_pendingMMIOld,1);
        //     `TCNT_CHECK_SIG_XZ(io_lsq_pendingst,io_lsq_pendingst,1);
        //     `TCNT_CHECK_SIG_XZ(io_lsq_pendingPtr_flag,io_lsq_pendingPtr_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_lsq_pendingPtr_value,io_lsq_pendingPtr_value,8);
        //     `TCNT_CHECK_SIG_XZ(io_robDeqPtr_flag,io_robDeqPtr_flag,1);
        //     `TCNT_CHECK_SIG_XZ(io_robDeqPtr_value,io_robDeqPtr_value,8);
        //     `TCNT_CHECK_SIG_XZ(io_csr_fflags_valid,io_csr_fflags_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_csr_fflags_bits,io_csr_fflags_bits,5);
        //     `TCNT_CHECK_SIG_XZ(io_csr_vxsat_valid,io_csr_vxsat_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_csr_vxsat_bits,io_csr_vxsat_bits,1);
        //     `TCNT_CHECK_SIG_XZ(io_csr_vstart_valid,io_csr_vstart_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_csr_vstart_bits,io_csr_vstart_bits,64);
        //     `TCNT_CHECK_SIG_XZ(io_csr_dirty_fs,io_csr_dirty_fs,1);
        //     `TCNT_CHECK_SIG_XZ(io_csr_dirty_vs,io_csr_dirty_vs,1);
        //     `TCNT_CHECK_SIG_XZ(io_csr_perfinfo_retiredInstr,io_csr_perfinfo_retiredInstr,7);
        //     `TCNT_CHECK_SIG_XZ(io_cpu_halt,io_cpu_halt,1);
        //     `TCNT_CHECK_SIG_XZ(io_wfi_wfiReq,io_wfi_wfiReq,1);
        //     `TCNT_CHECK_SIG_XZ(io_toDecode_isResumeVType,io_toDecode_isResumeVType,1);
        //     `TCNT_CHECK_SIG_XZ(io_toDecode_walkToArchVType,io_toDecode_walkToArchVType,1);
        //     `TCNT_CHECK_SIG_XZ(io_toDecode_walkVType_valid,io_toDecode_walkVType_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_toDecode_walkVType_bits_illegal,io_toDecode_walkVType_bits_illegal,1);
        //     `TCNT_CHECK_SIG_XZ(io_toDecode_walkVType_bits_vma,io_toDecode_walkVType_bits_vma,1);
        //     `TCNT_CHECK_SIG_XZ(io_toDecode_walkVType_bits_vta,io_toDecode_walkVType_bits_vta,1);
        //     `TCNT_CHECK_SIG_XZ(io_toDecode_walkVType_bits_vsew,io_toDecode_walkVType_bits_vsew,2);
        //     `TCNT_CHECK_SIG_XZ(io_toDecode_walkVType_bits_vlmul,io_toDecode_walkVType_bits_vlmul,3);
        //     `TCNT_CHECK_SIG_XZ(io_toDecode_commitVType_vtype_valid,io_toDecode_commitVType_vtype_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_toDecode_commitVType_vtype_bits_illegal,io_toDecode_commitVType_vtype_bits_illegal,1);
        //     `TCNT_CHECK_SIG_XZ(io_toDecode_commitVType_vtype_bits_vma,io_toDecode_commitVType_vtype_bits_vma,1);
        //     `TCNT_CHECK_SIG_XZ(io_toDecode_commitVType_vtype_bits_vta,io_toDecode_commitVType_vtype_bits_vta,1);
        //     `TCNT_CHECK_SIG_XZ(io_toDecode_commitVType_vtype_bits_vsew,io_toDecode_commitVType_vtype_bits_vsew,2);
        //     `TCNT_CHECK_SIG_XZ(io_toDecode_commitVType_vtype_bits_vlmul,io_toDecode_commitVType_vtype_bits_vlmul,3);
        //     `TCNT_CHECK_SIG_XZ(io_toDecode_commitVType_hasVsetvl,io_toDecode_commitVType_hasVsetvl,1);
        //     `TCNT_CHECK_SIG_XZ(io_readGPAMemAddr_valid,io_readGPAMemAddr_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_readGPAMemAddr_bits_ftqPtr_value,io_readGPAMemAddr_bits_ftqPtr_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_readGPAMemAddr_bits_ftqOffset,io_readGPAMemAddr_bits_ftqOffset,4);
        //     `TCNT_CHECK_SIG_XZ(io_toVecExcpMod_logicPhyRegMap_0_valid,io_toVecExcpMod_logicPhyRegMap_0_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_toVecExcpMod_logicPhyRegMap_0_bits_lreg,io_toVecExcpMod_logicPhyRegMap_0_bits_lreg,6);
        //     `TCNT_CHECK_SIG_XZ(io_toVecExcpMod_logicPhyRegMap_0_bits_preg,io_toVecExcpMod_logicPhyRegMap_0_bits_preg,7);
        //     `TCNT_CHECK_SIG_XZ(io_toVecExcpMod_logicPhyRegMap_1_valid,io_toVecExcpMod_logicPhyRegMap_1_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_toVecExcpMod_logicPhyRegMap_1_bits_lreg,io_toVecExcpMod_logicPhyRegMap_1_bits_lreg,6);
        //     `TCNT_CHECK_SIG_XZ(io_toVecExcpMod_logicPhyRegMap_1_bits_preg,io_toVecExcpMod_logicPhyRegMap_1_bits_preg,7);
        //     `TCNT_CHECK_SIG_XZ(io_toVecExcpMod_logicPhyRegMap_2_valid,io_toVecExcpMod_logicPhyRegMap_2_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_toVecExcpMod_logicPhyRegMap_2_bits_lreg,io_toVecExcpMod_logicPhyRegMap_2_bits_lreg,6);
        //     `TCNT_CHECK_SIG_XZ(io_toVecExcpMod_logicPhyRegMap_2_bits_preg,io_toVecExcpMod_logicPhyRegMap_2_bits_preg,7);
        //     `TCNT_CHECK_SIG_XZ(io_toVecExcpMod_logicPhyRegMap_3_valid,io_toVecExcpMod_logicPhyRegMap_3_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_toVecExcpMod_logicPhyRegMap_3_bits_lreg,io_toVecExcpMod_logicPhyRegMap_3_bits_lreg,6);
        //     `TCNT_CHECK_SIG_XZ(io_toVecExcpMod_logicPhyRegMap_3_bits_preg,io_toVecExcpMod_logicPhyRegMap_3_bits_preg,7);
        //     `TCNT_CHECK_SIG_XZ(io_toVecExcpMod_logicPhyRegMap_4_valid,io_toVecExcpMod_logicPhyRegMap_4_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_toVecExcpMod_logicPhyRegMap_4_bits_lreg,io_toVecExcpMod_logicPhyRegMap_4_bits_lreg,6);
        //     `TCNT_CHECK_SIG_XZ(io_toVecExcpMod_logicPhyRegMap_4_bits_preg,io_toVecExcpMod_logicPhyRegMap_4_bits_preg,7);
        //     `TCNT_CHECK_SIG_XZ(io_toVecExcpMod_logicPhyRegMap_5_valid,io_toVecExcpMod_logicPhyRegMap_5_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_toVecExcpMod_logicPhyRegMap_5_bits_lreg,io_toVecExcpMod_logicPhyRegMap_5_bits_lreg,6);
        //     `TCNT_CHECK_SIG_XZ(io_toVecExcpMod_logicPhyRegMap_5_bits_preg,io_toVecExcpMod_logicPhyRegMap_5_bits_preg,7);
        //     `TCNT_CHECK_SIG_XZ(io_toVecExcpMod_excpInfo_valid,io_toVecExcpMod_excpInfo_valid,1);
        //     `TCNT_CHECK_SIG_XZ(io_toVecExcpMod_excpInfo_bits_vstart,io_toVecExcpMod_excpInfo_bits_vstart,7);
        //     `TCNT_CHECK_SIG_XZ(io_toVecExcpMod_excpInfo_bits_vsew,io_toVecExcpMod_excpInfo_bits_vsew,2);
        //     `TCNT_CHECK_SIG_XZ(io_toVecExcpMod_excpInfo_bits_veew,io_toVecExcpMod_excpInfo_bits_veew,2);
        //     `TCNT_CHECK_SIG_XZ(io_toVecExcpMod_excpInfo_bits_vlmul,io_toVecExcpMod_excpInfo_bits_vlmul,3);
        //     `TCNT_CHECK_SIG_XZ(io_toVecExcpMod_excpInfo_bits_nf,io_toVecExcpMod_excpInfo_bits_nf,3);
        //     `TCNT_CHECK_SIG_XZ(io_toVecExcpMod_excpInfo_bits_isStride,io_toVecExcpMod_excpInfo_bits_isStride,1);
        //     `TCNT_CHECK_SIG_XZ(io_toVecExcpMod_excpInfo_bits_isIndexed,io_toVecExcpMod_excpInfo_bits_isIndexed,1);
        //     `TCNT_CHECK_SIG_XZ(io_toVecExcpMod_excpInfo_bits_isWhole,io_toVecExcpMod_excpInfo_bits_isWhole,1);
        //     `TCNT_CHECK_SIG_XZ(io_toVecExcpMod_excpInfo_bits_isVlm,io_toVecExcpMod_excpInfo_bits_isVlm,1);
        //     `TCNT_CHECK_SIG_XZ(io_storeDebugInfo_1_pc,io_storeDebugInfo_1_pc,50);
        //     `TCNT_CHECK_SIG_XZ(io_perf_0_value,io_perf_0_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_perf_1_value,io_perf_1_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_perf_2_value,io_perf_2_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_perf_3_value,io_perf_3_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_perf_4_value,io_perf_4_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_perf_5_value,io_perf_5_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_perf_6_value,io_perf_6_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_perf_7_value,io_perf_7_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_perf_8_value,io_perf_8_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_perf_9_value,io_perf_9_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_perf_10_value,io_perf_10_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_perf_11_value,io_perf_11_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_perf_12_value,io_perf_12_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_perf_13_value,io_perf_13_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_perf_14_value,io_perf_14_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_perf_15_value,io_perf_15_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_perf_16_value,io_perf_16_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_perf_17_value,io_perf_17_value,6);
        //     `TCNT_CHECK_SIG_XZ(io_error_0,io_error_0,1);

        // end
        //if(xxxTODOxxx==1'b1) begin
        //    mon_tr = Rob_output_agent_xaction::type_id::create("mon_tr");
        //    mon_tr.io_enq_canAccept = io_enq_canAccept;
        //    mon_tr.io_enq_canAcceptForDispatch = io_enq_canAcceptForDispatch;
        //    mon_tr.io_enq_isEmpty = io_enq_isEmpty;
        //    mon_tr.io_flushOut_valid = io_flushOut_valid;
        //    mon_tr.io_flushOut_bits_isRVC = io_flushOut_bits_isRVC;
        //    mon_tr.io_flushOut_bits_robIdx_flag = io_flushOut_bits_robIdx_flag;
        //    mon_tr.io_flushOut_bits_robIdx_value = io_flushOut_bits_robIdx_value;
        //    mon_tr.io_flushOut_bits_ftqIdx_flag = io_flushOut_bits_ftqIdx_flag;
        //    mon_tr.io_flushOut_bits_ftqIdx_value = io_flushOut_bits_ftqIdx_value;
        //    mon_tr.io_flushOut_bits_ftqOffset = io_flushOut_bits_ftqOffset;
        //    mon_tr.io_flushOut_bits_level = io_flushOut_bits_level;
        //    mon_tr.io_exception_valid = io_exception_valid;
        //    mon_tr.io_exception_bits_instr = io_exception_bits_instr;
        //    mon_tr.io_exception_bits_commitType = io_exception_bits_commitType;
        //    mon_tr.io_exception_bits_exceptionVec_0 = io_exception_bits_exceptionVec_0;
        //    mon_tr.io_exception_bits_exceptionVec_1 = io_exception_bits_exceptionVec_1;
        //    mon_tr.io_exception_bits_exceptionVec_2 = io_exception_bits_exceptionVec_2;
        //    mon_tr.io_exception_bits_exceptionVec_3 = io_exception_bits_exceptionVec_3;
        //    mon_tr.io_exception_bits_exceptionVec_4 = io_exception_bits_exceptionVec_4;
        //    mon_tr.io_exception_bits_exceptionVec_5 = io_exception_bits_exceptionVec_5;
        //    mon_tr.io_exception_bits_exceptionVec_6 = io_exception_bits_exceptionVec_6;
        //    mon_tr.io_exception_bits_exceptionVec_7 = io_exception_bits_exceptionVec_7;
        //    mon_tr.io_exception_bits_exceptionVec_8 = io_exception_bits_exceptionVec_8;
        //    mon_tr.io_exception_bits_exceptionVec_9 = io_exception_bits_exceptionVec_9;
        //    mon_tr.io_exception_bits_exceptionVec_10 = io_exception_bits_exceptionVec_10;
        //    mon_tr.io_exception_bits_exceptionVec_11 = io_exception_bits_exceptionVec_11;
        //    mon_tr.io_exception_bits_exceptionVec_12 = io_exception_bits_exceptionVec_12;
        //    mon_tr.io_exception_bits_exceptionVec_13 = io_exception_bits_exceptionVec_13;
        //    mon_tr.io_exception_bits_exceptionVec_14 = io_exception_bits_exceptionVec_14;
        //    mon_tr.io_exception_bits_exceptionVec_15 = io_exception_bits_exceptionVec_15;
        //    mon_tr.io_exception_bits_exceptionVec_16 = io_exception_bits_exceptionVec_16;
        //    mon_tr.io_exception_bits_exceptionVec_17 = io_exception_bits_exceptionVec_17;
        //    mon_tr.io_exception_bits_exceptionVec_18 = io_exception_bits_exceptionVec_18;
        //    mon_tr.io_exception_bits_exceptionVec_19 = io_exception_bits_exceptionVec_19;
        //    mon_tr.io_exception_bits_exceptionVec_20 = io_exception_bits_exceptionVec_20;
        //    mon_tr.io_exception_bits_exceptionVec_21 = io_exception_bits_exceptionVec_21;
        //    mon_tr.io_exception_bits_exceptionVec_22 = io_exception_bits_exceptionVec_22;
        //    mon_tr.io_exception_bits_exceptionVec_23 = io_exception_bits_exceptionVec_23;
        //    mon_tr.io_exception_bits_isPcBkpt = io_exception_bits_isPcBkpt;
        //    mon_tr.io_exception_bits_isFetchMalAddr = io_exception_bits_isFetchMalAddr;
        //    mon_tr.io_exception_bits_gpaddr = io_exception_bits_gpaddr;
        //    mon_tr.io_exception_bits_singleStep = io_exception_bits_singleStep;
        //    mon_tr.io_exception_bits_crossPageIPFFix = io_exception_bits_crossPageIPFFix;
        //    mon_tr.io_exception_bits_isInterrupt = io_exception_bits_isInterrupt;
        //    mon_tr.io_exception_bits_isHls = io_exception_bits_isHls;
        //    mon_tr.io_exception_bits_trigger = io_exception_bits_trigger;
        //    mon_tr.io_exception_bits_isForVSnonLeafPTE = io_exception_bits_isForVSnonLeafPTE;
        //    mon_tr.io_commits_isCommit = io_commits_isCommit;
        //    mon_tr.io_commits_commitValid_0 = io_commits_commitValid_0;
        //    mon_tr.io_commits_commitValid_1 = io_commits_commitValid_1;
        //    mon_tr.io_commits_commitValid_2 = io_commits_commitValid_2;
        //    mon_tr.io_commits_commitValid_3 = io_commits_commitValid_3;
        //    mon_tr.io_commits_commitValid_4 = io_commits_commitValid_4;
        //    mon_tr.io_commits_commitValid_5 = io_commits_commitValid_5;
        //    mon_tr.io_commits_commitValid_6 = io_commits_commitValid_6;
        //    mon_tr.io_commits_commitValid_7 = io_commits_commitValid_7;
        //    mon_tr.io_commits_isWalk = io_commits_isWalk;
        //    mon_tr.io_commits_walkValid_0 = io_commits_walkValid_0;
        //    mon_tr.io_commits_walkValid_1 = io_commits_walkValid_1;
        //    mon_tr.io_commits_walkValid_2 = io_commits_walkValid_2;
        //    mon_tr.io_commits_walkValid_3 = io_commits_walkValid_3;
        //    mon_tr.io_commits_walkValid_4 = io_commits_walkValid_4;
        //    mon_tr.io_commits_walkValid_5 = io_commits_walkValid_5;
        //    mon_tr.io_commits_walkValid_6 = io_commits_walkValid_6;
        //    mon_tr.io_commits_walkValid_7 = io_commits_walkValid_7;
        //    mon_tr.io_commits_info_0_walk_v = io_commits_info_0_walk_v;
        //    mon_tr.io_commits_info_0_commit_v = io_commits_info_0_commit_v;
        //    mon_tr.io_commits_info_0_commit_w = io_commits_info_0_commit_w;
        //    mon_tr.io_commits_info_0_realDestSize = io_commits_info_0_realDestSize;
        //    mon_tr.io_commits_info_0_interrupt_safe = io_commits_info_0_interrupt_safe;
        //    mon_tr.io_commits_info_0_wflags = io_commits_info_0_wflags;
        //    mon_tr.io_commits_info_0_fflags = io_commits_info_0_fflags;
        //    mon_tr.io_commits_info_0_vxsat = io_commits_info_0_vxsat;
        //    mon_tr.io_commits_info_0_isRVC = io_commits_info_0_isRVC;
        //    mon_tr.io_commits_info_0_isVset = io_commits_info_0_isVset;
        //    mon_tr.io_commits_info_0_isHls = io_commits_info_0_isHls;
        //    mon_tr.io_commits_info_0_isVls = io_commits_info_0_isVls;
        //    mon_tr.io_commits_info_0_vls = io_commits_info_0_vls;
        //    mon_tr.io_commits_info_0_mmio = io_commits_info_0_mmio;
        //    mon_tr.io_commits_info_0_commitType = io_commits_info_0_commitType;
        //    mon_tr.io_commits_info_0_ftqIdx_flag = io_commits_info_0_ftqIdx_flag;
        //    mon_tr.io_commits_info_0_ftqIdx_value = io_commits_info_0_ftqIdx_value;
        //    mon_tr.io_commits_info_0_ftqOffset = io_commits_info_0_ftqOffset;
        //    mon_tr.io_commits_info_0_instrSize = io_commits_info_0_instrSize;
        //    mon_tr.io_commits_info_0_fpWen = io_commits_info_0_fpWen;
        //    mon_tr.io_commits_info_0_rfWen = io_commits_info_0_rfWen;
        //    mon_tr.io_commits_info_0_needFlush = io_commits_info_0_needFlush;
        //    mon_tr.io_commits_info_0_traceBlockInPipe_itype = io_commits_info_0_traceBlockInPipe_itype;
        //    mon_tr.io_commits_info_0_traceBlockInPipe_iretire = io_commits_info_0_traceBlockInPipe_iretire;
        //    mon_tr.io_commits_info_0_traceBlockInPipe_ilastsize = io_commits_info_0_traceBlockInPipe_ilastsize;
        //    mon_tr.io_commits_info_0_debug_pc = io_commits_info_0_debug_pc;
        //    mon_tr.io_commits_info_0_debug_instr = io_commits_info_0_debug_instr;
        //    mon_tr.io_commits_info_0_debug_ldest = io_commits_info_0_debug_ldest;
        //    mon_tr.io_commits_info_0_debug_pdest = io_commits_info_0_debug_pdest;
        //    mon_tr.io_commits_info_0_debug_otherPdest_0 = io_commits_info_0_debug_otherPdest_0;
        //    mon_tr.io_commits_info_0_debug_otherPdest_1 = io_commits_info_0_debug_otherPdest_1;
        //    mon_tr.io_commits_info_0_debug_otherPdest_2 = io_commits_info_0_debug_otherPdest_2;
        //    mon_tr.io_commits_info_0_debug_otherPdest_3 = io_commits_info_0_debug_otherPdest_3;
        //    mon_tr.io_commits_info_0_debug_otherPdest_4 = io_commits_info_0_debug_otherPdest_4;
        //    mon_tr.io_commits_info_0_debug_otherPdest_5 = io_commits_info_0_debug_otherPdest_5;
        //    mon_tr.io_commits_info_0_debug_otherPdest_6 = io_commits_info_0_debug_otherPdest_6;
        //    mon_tr.io_commits_info_0_debug_fuType = io_commits_info_0_debug_fuType;
        //    mon_tr.io_commits_info_0_dirtyFs = io_commits_info_0_dirtyFs;
        //    mon_tr.io_commits_info_0_dirtyVs = io_commits_info_0_dirtyVs;
        //    mon_tr.io_commits_info_1_walk_v = io_commits_info_1_walk_v;
        //    mon_tr.io_commits_info_1_commit_v = io_commits_info_1_commit_v;
        //    mon_tr.io_commits_info_1_commit_w = io_commits_info_1_commit_w;
        //    mon_tr.io_commits_info_1_realDestSize = io_commits_info_1_realDestSize;
        //    mon_tr.io_commits_info_1_interrupt_safe = io_commits_info_1_interrupt_safe;
        //    mon_tr.io_commits_info_1_wflags = io_commits_info_1_wflags;
        //    mon_tr.io_commits_info_1_fflags = io_commits_info_1_fflags;
        //    mon_tr.io_commits_info_1_vxsat = io_commits_info_1_vxsat;
        //    mon_tr.io_commits_info_1_isRVC = io_commits_info_1_isRVC;
        //    mon_tr.io_commits_info_1_isVset = io_commits_info_1_isVset;
        //    mon_tr.io_commits_info_1_isHls = io_commits_info_1_isHls;
        //    mon_tr.io_commits_info_1_isVls = io_commits_info_1_isVls;
        //    mon_tr.io_commits_info_1_vls = io_commits_info_1_vls;
        //    mon_tr.io_commits_info_1_mmio = io_commits_info_1_mmio;
        //    mon_tr.io_commits_info_1_commitType = io_commits_info_1_commitType;
        //    mon_tr.io_commits_info_1_ftqIdx_flag = io_commits_info_1_ftqIdx_flag;
        //    mon_tr.io_commits_info_1_ftqIdx_value = io_commits_info_1_ftqIdx_value;
        //    mon_tr.io_commits_info_1_ftqOffset = io_commits_info_1_ftqOffset;
        //    mon_tr.io_commits_info_1_instrSize = io_commits_info_1_instrSize;
        //    mon_tr.io_commits_info_1_fpWen = io_commits_info_1_fpWen;
        //    mon_tr.io_commits_info_1_rfWen = io_commits_info_1_rfWen;
        //    mon_tr.io_commits_info_1_needFlush = io_commits_info_1_needFlush;
        //    mon_tr.io_commits_info_1_traceBlockInPipe_itype = io_commits_info_1_traceBlockInPipe_itype;
        //    mon_tr.io_commits_info_1_traceBlockInPipe_iretire = io_commits_info_1_traceBlockInPipe_iretire;
        //    mon_tr.io_commits_info_1_traceBlockInPipe_ilastsize = io_commits_info_1_traceBlockInPipe_ilastsize;
        //    mon_tr.io_commits_info_1_debug_pc = io_commits_info_1_debug_pc;
        //    mon_tr.io_commits_info_1_debug_instr = io_commits_info_1_debug_instr;
        //    mon_tr.io_commits_info_1_debug_ldest = io_commits_info_1_debug_ldest;
        //    mon_tr.io_commits_info_1_debug_pdest = io_commits_info_1_debug_pdest;
        //    mon_tr.io_commits_info_1_debug_otherPdest_0 = io_commits_info_1_debug_otherPdest_0;
        //    mon_tr.io_commits_info_1_debug_otherPdest_1 = io_commits_info_1_debug_otherPdest_1;
        //    mon_tr.io_commits_info_1_debug_otherPdest_2 = io_commits_info_1_debug_otherPdest_2;
        //    mon_tr.io_commits_info_1_debug_otherPdest_3 = io_commits_info_1_debug_otherPdest_3;
        //    mon_tr.io_commits_info_1_debug_otherPdest_4 = io_commits_info_1_debug_otherPdest_4;
        //    mon_tr.io_commits_info_1_debug_otherPdest_5 = io_commits_info_1_debug_otherPdest_5;
        //    mon_tr.io_commits_info_1_debug_otherPdest_6 = io_commits_info_1_debug_otherPdest_6;
        //    mon_tr.io_commits_info_1_debug_fuType = io_commits_info_1_debug_fuType;
        //    mon_tr.io_commits_info_1_dirtyFs = io_commits_info_1_dirtyFs;
        //    mon_tr.io_commits_info_1_dirtyVs = io_commits_info_1_dirtyVs;
        //    mon_tr.io_commits_info_2_walk_v = io_commits_info_2_walk_v;
        //    mon_tr.io_commits_info_2_commit_v = io_commits_info_2_commit_v;
        //    mon_tr.io_commits_info_2_commit_w = io_commits_info_2_commit_w;
        //    mon_tr.io_commits_info_2_realDestSize = io_commits_info_2_realDestSize;
        //    mon_tr.io_commits_info_2_interrupt_safe = io_commits_info_2_interrupt_safe;
        //    mon_tr.io_commits_info_2_wflags = io_commits_info_2_wflags;
        //    mon_tr.io_commits_info_2_fflags = io_commits_info_2_fflags;
        //    mon_tr.io_commits_info_2_vxsat = io_commits_info_2_vxsat;
        //    mon_tr.io_commits_info_2_isRVC = io_commits_info_2_isRVC;
        //    mon_tr.io_commits_info_2_isVset = io_commits_info_2_isVset;
        //    mon_tr.io_commits_info_2_isHls = io_commits_info_2_isHls;
        //    mon_tr.io_commits_info_2_isVls = io_commits_info_2_isVls;
        //    mon_tr.io_commits_info_2_vls = io_commits_info_2_vls;
        //    mon_tr.io_commits_info_2_mmio = io_commits_info_2_mmio;
        //    mon_tr.io_commits_info_2_commitType = io_commits_info_2_commitType;
        //    mon_tr.io_commits_info_2_ftqIdx_flag = io_commits_info_2_ftqIdx_flag;
        //    mon_tr.io_commits_info_2_ftqIdx_value = io_commits_info_2_ftqIdx_value;
        //    mon_tr.io_commits_info_2_ftqOffset = io_commits_info_2_ftqOffset;
        //    mon_tr.io_commits_info_2_instrSize = io_commits_info_2_instrSize;
        //    mon_tr.io_commits_info_2_fpWen = io_commits_info_2_fpWen;
        //    mon_tr.io_commits_info_2_rfWen = io_commits_info_2_rfWen;
        //    mon_tr.io_commits_info_2_needFlush = io_commits_info_2_needFlush;
        //    mon_tr.io_commits_info_2_traceBlockInPipe_itype = io_commits_info_2_traceBlockInPipe_itype;
        //    mon_tr.io_commits_info_2_traceBlockInPipe_iretire = io_commits_info_2_traceBlockInPipe_iretire;
        //    mon_tr.io_commits_info_2_traceBlockInPipe_ilastsize = io_commits_info_2_traceBlockInPipe_ilastsize;
        //    mon_tr.io_commits_info_2_debug_pc = io_commits_info_2_debug_pc;
        //    mon_tr.io_commits_info_2_debug_instr = io_commits_info_2_debug_instr;
        //    mon_tr.io_commits_info_2_debug_ldest = io_commits_info_2_debug_ldest;
        //    mon_tr.io_commits_info_2_debug_pdest = io_commits_info_2_debug_pdest;
        //    mon_tr.io_commits_info_2_debug_otherPdest_0 = io_commits_info_2_debug_otherPdest_0;
        //    mon_tr.io_commits_info_2_debug_otherPdest_1 = io_commits_info_2_debug_otherPdest_1;
        //    mon_tr.io_commits_info_2_debug_otherPdest_2 = io_commits_info_2_debug_otherPdest_2;
        //    mon_tr.io_commits_info_2_debug_otherPdest_3 = io_commits_info_2_debug_otherPdest_3;
        //    mon_tr.io_commits_info_2_debug_otherPdest_4 = io_commits_info_2_debug_otherPdest_4;
        //    mon_tr.io_commits_info_2_debug_otherPdest_5 = io_commits_info_2_debug_otherPdest_5;
        //    mon_tr.io_commits_info_2_debug_otherPdest_6 = io_commits_info_2_debug_otherPdest_6;
        //    mon_tr.io_commits_info_2_debug_fuType = io_commits_info_2_debug_fuType;
        //    mon_tr.io_commits_info_2_dirtyFs = io_commits_info_2_dirtyFs;
        //    mon_tr.io_commits_info_2_dirtyVs = io_commits_info_2_dirtyVs;
        //    mon_tr.io_commits_info_3_walk_v = io_commits_info_3_walk_v;
        //    mon_tr.io_commits_info_3_commit_v = io_commits_info_3_commit_v;
        //    mon_tr.io_commits_info_3_commit_w = io_commits_info_3_commit_w;
        //    mon_tr.io_commits_info_3_realDestSize = io_commits_info_3_realDestSize;
        //    mon_tr.io_commits_info_3_interrupt_safe = io_commits_info_3_interrupt_safe;
        //    mon_tr.io_commits_info_3_wflags = io_commits_info_3_wflags;
        //    mon_tr.io_commits_info_3_fflags = io_commits_info_3_fflags;
        //    mon_tr.io_commits_info_3_vxsat = io_commits_info_3_vxsat;
        //    mon_tr.io_commits_info_3_isRVC = io_commits_info_3_isRVC;
        //    mon_tr.io_commits_info_3_isVset = io_commits_info_3_isVset;
        //    mon_tr.io_commits_info_3_isHls = io_commits_info_3_isHls;
        //    mon_tr.io_commits_info_3_isVls = io_commits_info_3_isVls;
        //    mon_tr.io_commits_info_3_vls = io_commits_info_3_vls;
        //    mon_tr.io_commits_info_3_mmio = io_commits_info_3_mmio;
        //    mon_tr.io_commits_info_3_commitType = io_commits_info_3_commitType;
        //    mon_tr.io_commits_info_3_ftqIdx_flag = io_commits_info_3_ftqIdx_flag;
        //    mon_tr.io_commits_info_3_ftqIdx_value = io_commits_info_3_ftqIdx_value;
        //    mon_tr.io_commits_info_3_ftqOffset = io_commits_info_3_ftqOffset;
        //    mon_tr.io_commits_info_3_instrSize = io_commits_info_3_instrSize;
        //    mon_tr.io_commits_info_3_fpWen = io_commits_info_3_fpWen;
        //    mon_tr.io_commits_info_3_rfWen = io_commits_info_3_rfWen;
        //    mon_tr.io_commits_info_3_needFlush = io_commits_info_3_needFlush;
        //    mon_tr.io_commits_info_3_traceBlockInPipe_itype = io_commits_info_3_traceBlockInPipe_itype;
        //    mon_tr.io_commits_info_3_traceBlockInPipe_iretire = io_commits_info_3_traceBlockInPipe_iretire;
        //    mon_tr.io_commits_info_3_traceBlockInPipe_ilastsize = io_commits_info_3_traceBlockInPipe_ilastsize;
        //    mon_tr.io_commits_info_3_debug_pc = io_commits_info_3_debug_pc;
        //    mon_tr.io_commits_info_3_debug_instr = io_commits_info_3_debug_instr;
        //    mon_tr.io_commits_info_3_debug_ldest = io_commits_info_3_debug_ldest;
        //    mon_tr.io_commits_info_3_debug_pdest = io_commits_info_3_debug_pdest;
        //    mon_tr.io_commits_info_3_debug_otherPdest_0 = io_commits_info_3_debug_otherPdest_0;
        //    mon_tr.io_commits_info_3_debug_otherPdest_1 = io_commits_info_3_debug_otherPdest_1;
        //    mon_tr.io_commits_info_3_debug_otherPdest_2 = io_commits_info_3_debug_otherPdest_2;
        //    mon_tr.io_commits_info_3_debug_otherPdest_3 = io_commits_info_3_debug_otherPdest_3;
        //    mon_tr.io_commits_info_3_debug_otherPdest_4 = io_commits_info_3_debug_otherPdest_4;
        //    mon_tr.io_commits_info_3_debug_otherPdest_5 = io_commits_info_3_debug_otherPdest_5;
        //    mon_tr.io_commits_info_3_debug_otherPdest_6 = io_commits_info_3_debug_otherPdest_6;
        //    mon_tr.io_commits_info_3_debug_fuType = io_commits_info_3_debug_fuType;
        //    mon_tr.io_commits_info_3_dirtyFs = io_commits_info_3_dirtyFs;
        //    mon_tr.io_commits_info_3_dirtyVs = io_commits_info_3_dirtyVs;
        //    mon_tr.io_commits_info_4_walk_v = io_commits_info_4_walk_v;
        //    mon_tr.io_commits_info_4_commit_v = io_commits_info_4_commit_v;
        //    mon_tr.io_commits_info_4_commit_w = io_commits_info_4_commit_w;
        //    mon_tr.io_commits_info_4_realDestSize = io_commits_info_4_realDestSize;
        //    mon_tr.io_commits_info_4_interrupt_safe = io_commits_info_4_interrupt_safe;
        //    mon_tr.io_commits_info_4_wflags = io_commits_info_4_wflags;
        //    mon_tr.io_commits_info_4_fflags = io_commits_info_4_fflags;
        //    mon_tr.io_commits_info_4_vxsat = io_commits_info_4_vxsat;
        //    mon_tr.io_commits_info_4_isRVC = io_commits_info_4_isRVC;
        //    mon_tr.io_commits_info_4_isVset = io_commits_info_4_isVset;
        //    mon_tr.io_commits_info_4_isHls = io_commits_info_4_isHls;
        //    mon_tr.io_commits_info_4_isVls = io_commits_info_4_isVls;
        //    mon_tr.io_commits_info_4_vls = io_commits_info_4_vls;
        //    mon_tr.io_commits_info_4_mmio = io_commits_info_4_mmio;
        //    mon_tr.io_commits_info_4_commitType = io_commits_info_4_commitType;
        //    mon_tr.io_commits_info_4_ftqIdx_flag = io_commits_info_4_ftqIdx_flag;
        //    mon_tr.io_commits_info_4_ftqIdx_value = io_commits_info_4_ftqIdx_value;
        //    mon_tr.io_commits_info_4_ftqOffset = io_commits_info_4_ftqOffset;
        //    mon_tr.io_commits_info_4_instrSize = io_commits_info_4_instrSize;
        //    mon_tr.io_commits_info_4_fpWen = io_commits_info_4_fpWen;
        //    mon_tr.io_commits_info_4_rfWen = io_commits_info_4_rfWen;
        //    mon_tr.io_commits_info_4_needFlush = io_commits_info_4_needFlush;
        //    mon_tr.io_commits_info_4_traceBlockInPipe_itype = io_commits_info_4_traceBlockInPipe_itype;
        //    mon_tr.io_commits_info_4_traceBlockInPipe_iretire = io_commits_info_4_traceBlockInPipe_iretire;
        //    mon_tr.io_commits_info_4_traceBlockInPipe_ilastsize = io_commits_info_4_traceBlockInPipe_ilastsize;
        //    mon_tr.io_commits_info_4_debug_pc = io_commits_info_4_debug_pc;
        //    mon_tr.io_commits_info_4_debug_instr = io_commits_info_4_debug_instr;
        //    mon_tr.io_commits_info_4_debug_ldest = io_commits_info_4_debug_ldest;
        //    mon_tr.io_commits_info_4_debug_pdest = io_commits_info_4_debug_pdest;
        //    mon_tr.io_commits_info_4_debug_otherPdest_0 = io_commits_info_4_debug_otherPdest_0;
        //    mon_tr.io_commits_info_4_debug_otherPdest_1 = io_commits_info_4_debug_otherPdest_1;
        //    mon_tr.io_commits_info_4_debug_otherPdest_2 = io_commits_info_4_debug_otherPdest_2;
        //    mon_tr.io_commits_info_4_debug_otherPdest_3 = io_commits_info_4_debug_otherPdest_3;
        //    mon_tr.io_commits_info_4_debug_otherPdest_4 = io_commits_info_4_debug_otherPdest_4;
        //    mon_tr.io_commits_info_4_debug_otherPdest_5 = io_commits_info_4_debug_otherPdest_5;
        //    mon_tr.io_commits_info_4_debug_otherPdest_6 = io_commits_info_4_debug_otherPdest_6;
        //    mon_tr.io_commits_info_4_debug_fuType = io_commits_info_4_debug_fuType;
        //    mon_tr.io_commits_info_4_dirtyFs = io_commits_info_4_dirtyFs;
        //    mon_tr.io_commits_info_4_dirtyVs = io_commits_info_4_dirtyVs;
        //    mon_tr.io_commits_info_5_walk_v = io_commits_info_5_walk_v;
        //    mon_tr.io_commits_info_5_commit_v = io_commits_info_5_commit_v;
        //    mon_tr.io_commits_info_5_commit_w = io_commits_info_5_commit_w;
        //    mon_tr.io_commits_info_5_realDestSize = io_commits_info_5_realDestSize;
        //    mon_tr.io_commits_info_5_interrupt_safe = io_commits_info_5_interrupt_safe;
        //    mon_tr.io_commits_info_5_wflags = io_commits_info_5_wflags;
        //    mon_tr.io_commits_info_5_fflags = io_commits_info_5_fflags;
        //    mon_tr.io_commits_info_5_vxsat = io_commits_info_5_vxsat;
        //    mon_tr.io_commits_info_5_isRVC = io_commits_info_5_isRVC;
        //    mon_tr.io_commits_info_5_isVset = io_commits_info_5_isVset;
        //    mon_tr.io_commits_info_5_isHls = io_commits_info_5_isHls;
        //    mon_tr.io_commits_info_5_isVls = io_commits_info_5_isVls;
        //    mon_tr.io_commits_info_5_vls = io_commits_info_5_vls;
        //    mon_tr.io_commits_info_5_mmio = io_commits_info_5_mmio;
        //    mon_tr.io_commits_info_5_commitType = io_commits_info_5_commitType;
        //    mon_tr.io_commits_info_5_ftqIdx_flag = io_commits_info_5_ftqIdx_flag;
        //    mon_tr.io_commits_info_5_ftqIdx_value = io_commits_info_5_ftqIdx_value;
        //    mon_tr.io_commits_info_5_ftqOffset = io_commits_info_5_ftqOffset;
        //    mon_tr.io_commits_info_5_instrSize = io_commits_info_5_instrSize;
        //    mon_tr.io_commits_info_5_fpWen = io_commits_info_5_fpWen;
        //    mon_tr.io_commits_info_5_rfWen = io_commits_info_5_rfWen;
        //    mon_tr.io_commits_info_5_needFlush = io_commits_info_5_needFlush;
        //    mon_tr.io_commits_info_5_traceBlockInPipe_itype = io_commits_info_5_traceBlockInPipe_itype;
        //    mon_tr.io_commits_info_5_traceBlockInPipe_iretire = io_commits_info_5_traceBlockInPipe_iretire;
        //    mon_tr.io_commits_info_5_traceBlockInPipe_ilastsize = io_commits_info_5_traceBlockInPipe_ilastsize;
        //    mon_tr.io_commits_info_5_debug_pc = io_commits_info_5_debug_pc;
        //    mon_tr.io_commits_info_5_debug_instr = io_commits_info_5_debug_instr;
        //    mon_tr.io_commits_info_5_debug_ldest = io_commits_info_5_debug_ldest;
        //    mon_tr.io_commits_info_5_debug_pdest = io_commits_info_5_debug_pdest;
        //    mon_tr.io_commits_info_5_debug_otherPdest_0 = io_commits_info_5_debug_otherPdest_0;
        //    mon_tr.io_commits_info_5_debug_otherPdest_1 = io_commits_info_5_debug_otherPdest_1;
        //    mon_tr.io_commits_info_5_debug_otherPdest_2 = io_commits_info_5_debug_otherPdest_2;
        //    mon_tr.io_commits_info_5_debug_otherPdest_3 = io_commits_info_5_debug_otherPdest_3;
        //    mon_tr.io_commits_info_5_debug_otherPdest_4 = io_commits_info_5_debug_otherPdest_4;
        //    mon_tr.io_commits_info_5_debug_otherPdest_5 = io_commits_info_5_debug_otherPdest_5;
        //    mon_tr.io_commits_info_5_debug_otherPdest_6 = io_commits_info_5_debug_otherPdest_6;
        //    mon_tr.io_commits_info_5_debug_fuType = io_commits_info_5_debug_fuType;
        //    mon_tr.io_commits_info_5_dirtyFs = io_commits_info_5_dirtyFs;
        //    mon_tr.io_commits_info_5_dirtyVs = io_commits_info_5_dirtyVs;
        //    mon_tr.io_commits_info_6_walk_v = io_commits_info_6_walk_v;
        //    mon_tr.io_commits_info_6_commit_v = io_commits_info_6_commit_v;
        //    mon_tr.io_commits_info_6_commit_w = io_commits_info_6_commit_w;
        //    mon_tr.io_commits_info_6_realDestSize = io_commits_info_6_realDestSize;
        //    mon_tr.io_commits_info_6_interrupt_safe = io_commits_info_6_interrupt_safe;
        //    mon_tr.io_commits_info_6_wflags = io_commits_info_6_wflags;
        //    mon_tr.io_commits_info_6_fflags = io_commits_info_6_fflags;
        //    mon_tr.io_commits_info_6_vxsat = io_commits_info_6_vxsat;
        //    mon_tr.io_commits_info_6_isRVC = io_commits_info_6_isRVC;
        //    mon_tr.io_commits_info_6_isVset = io_commits_info_6_isVset;
        //    mon_tr.io_commits_info_6_isHls = io_commits_info_6_isHls;
        //    mon_tr.io_commits_info_6_isVls = io_commits_info_6_isVls;
        //    mon_tr.io_commits_info_6_vls = io_commits_info_6_vls;
        //    mon_tr.io_commits_info_6_mmio = io_commits_info_6_mmio;
        //    mon_tr.io_commits_info_6_commitType = io_commits_info_6_commitType;
        //    mon_tr.io_commits_info_6_ftqIdx_flag = io_commits_info_6_ftqIdx_flag;
        //    mon_tr.io_commits_info_6_ftqIdx_value = io_commits_info_6_ftqIdx_value;
        //    mon_tr.io_commits_info_6_ftqOffset = io_commits_info_6_ftqOffset;
        //    mon_tr.io_commits_info_6_instrSize = io_commits_info_6_instrSize;
        //    mon_tr.io_commits_info_6_fpWen = io_commits_info_6_fpWen;
        //    mon_tr.io_commits_info_6_rfWen = io_commits_info_6_rfWen;
        //    mon_tr.io_commits_info_6_needFlush = io_commits_info_6_needFlush;
        //    mon_tr.io_commits_info_6_traceBlockInPipe_itype = io_commits_info_6_traceBlockInPipe_itype;
        //    mon_tr.io_commits_info_6_traceBlockInPipe_iretire = io_commits_info_6_traceBlockInPipe_iretire;
        //    mon_tr.io_commits_info_6_traceBlockInPipe_ilastsize = io_commits_info_6_traceBlockInPipe_ilastsize;
        //    mon_tr.io_commits_info_6_debug_pc = io_commits_info_6_debug_pc;
        //    mon_tr.io_commits_info_6_debug_instr = io_commits_info_6_debug_instr;
        //    mon_tr.io_commits_info_6_debug_ldest = io_commits_info_6_debug_ldest;
        //    mon_tr.io_commits_info_6_debug_pdest = io_commits_info_6_debug_pdest;
        //    mon_tr.io_commits_info_6_debug_otherPdest_0 = io_commits_info_6_debug_otherPdest_0;
        //    mon_tr.io_commits_info_6_debug_otherPdest_1 = io_commits_info_6_debug_otherPdest_1;
        //    mon_tr.io_commits_info_6_debug_otherPdest_2 = io_commits_info_6_debug_otherPdest_2;
        //    mon_tr.io_commits_info_6_debug_otherPdest_3 = io_commits_info_6_debug_otherPdest_3;
        //    mon_tr.io_commits_info_6_debug_otherPdest_4 = io_commits_info_6_debug_otherPdest_4;
        //    mon_tr.io_commits_info_6_debug_otherPdest_5 = io_commits_info_6_debug_otherPdest_5;
        //    mon_tr.io_commits_info_6_debug_otherPdest_6 = io_commits_info_6_debug_otherPdest_6;
        //    mon_tr.io_commits_info_6_debug_fuType = io_commits_info_6_debug_fuType;
        //    mon_tr.io_commits_info_6_dirtyFs = io_commits_info_6_dirtyFs;
        //    mon_tr.io_commits_info_6_dirtyVs = io_commits_info_6_dirtyVs;
        //    mon_tr.io_commits_info_7_walk_v = io_commits_info_7_walk_v;
        //    mon_tr.io_commits_info_7_commit_v = io_commits_info_7_commit_v;
        //    mon_tr.io_commits_info_7_commit_w = io_commits_info_7_commit_w;
        //    mon_tr.io_commits_info_7_realDestSize = io_commits_info_7_realDestSize;
        //    mon_tr.io_commits_info_7_interrupt_safe = io_commits_info_7_interrupt_safe;
        //    mon_tr.io_commits_info_7_wflags = io_commits_info_7_wflags;
        //    mon_tr.io_commits_info_7_fflags = io_commits_info_7_fflags;
        //    mon_tr.io_commits_info_7_vxsat = io_commits_info_7_vxsat;
        //    mon_tr.io_commits_info_7_isRVC = io_commits_info_7_isRVC;
        //    mon_tr.io_commits_info_7_isVset = io_commits_info_7_isVset;
        //    mon_tr.io_commits_info_7_isHls = io_commits_info_7_isHls;
        //    mon_tr.io_commits_info_7_isVls = io_commits_info_7_isVls;
        //    mon_tr.io_commits_info_7_vls = io_commits_info_7_vls;
        //    mon_tr.io_commits_info_7_mmio = io_commits_info_7_mmio;
        //    mon_tr.io_commits_info_7_commitType = io_commits_info_7_commitType;
        //    mon_tr.io_commits_info_7_ftqIdx_flag = io_commits_info_7_ftqIdx_flag;
        //    mon_tr.io_commits_info_7_ftqIdx_value = io_commits_info_7_ftqIdx_value;
        //    mon_tr.io_commits_info_7_ftqOffset = io_commits_info_7_ftqOffset;
        //    mon_tr.io_commits_info_7_instrSize = io_commits_info_7_instrSize;
        //    mon_tr.io_commits_info_7_fpWen = io_commits_info_7_fpWen;
        //    mon_tr.io_commits_info_7_rfWen = io_commits_info_7_rfWen;
        //    mon_tr.io_commits_info_7_needFlush = io_commits_info_7_needFlush;
        //    mon_tr.io_commits_info_7_traceBlockInPipe_itype = io_commits_info_7_traceBlockInPipe_itype;
        //    mon_tr.io_commits_info_7_traceBlockInPipe_iretire = io_commits_info_7_traceBlockInPipe_iretire;
        //    mon_tr.io_commits_info_7_traceBlockInPipe_ilastsize = io_commits_info_7_traceBlockInPipe_ilastsize;
        //    mon_tr.io_commits_info_7_debug_pc = io_commits_info_7_debug_pc;
        //    mon_tr.io_commits_info_7_debug_instr = io_commits_info_7_debug_instr;
        //    mon_tr.io_commits_info_7_debug_ldest = io_commits_info_7_debug_ldest;
        //    mon_tr.io_commits_info_7_debug_pdest = io_commits_info_7_debug_pdest;
        //    mon_tr.io_commits_info_7_debug_otherPdest_0 = io_commits_info_7_debug_otherPdest_0;
        //    mon_tr.io_commits_info_7_debug_otherPdest_1 = io_commits_info_7_debug_otherPdest_1;
        //    mon_tr.io_commits_info_7_debug_otherPdest_2 = io_commits_info_7_debug_otherPdest_2;
        //    mon_tr.io_commits_info_7_debug_otherPdest_3 = io_commits_info_7_debug_otherPdest_3;
        //    mon_tr.io_commits_info_7_debug_otherPdest_4 = io_commits_info_7_debug_otherPdest_4;
        //    mon_tr.io_commits_info_7_debug_otherPdest_5 = io_commits_info_7_debug_otherPdest_5;
        //    mon_tr.io_commits_info_7_debug_otherPdest_6 = io_commits_info_7_debug_otherPdest_6;
        //    mon_tr.io_commits_info_7_debug_fuType = io_commits_info_7_debug_fuType;
        //    mon_tr.io_commits_info_7_dirtyFs = io_commits_info_7_dirtyFs;
        //    mon_tr.io_commits_info_7_dirtyVs = io_commits_info_7_dirtyVs;
        //    mon_tr.io_commits_robIdx_0_flag = io_commits_robIdx_0_flag;
        //    mon_tr.io_commits_robIdx_0_value = io_commits_robIdx_0_value;
        //    mon_tr.io_commits_robIdx_1_flag = io_commits_robIdx_1_flag;
        //    mon_tr.io_commits_robIdx_1_value = io_commits_robIdx_1_value;
        //    mon_tr.io_commits_robIdx_2_flag = io_commits_robIdx_2_flag;
        //    mon_tr.io_commits_robIdx_2_value = io_commits_robIdx_2_value;
        //    mon_tr.io_commits_robIdx_3_flag = io_commits_robIdx_3_flag;
        //    mon_tr.io_commits_robIdx_3_value = io_commits_robIdx_3_value;
        //    mon_tr.io_commits_robIdx_4_flag = io_commits_robIdx_4_flag;
        //    mon_tr.io_commits_robIdx_4_value = io_commits_robIdx_4_value;
        //    mon_tr.io_commits_robIdx_5_flag = io_commits_robIdx_5_flag;
        //    mon_tr.io_commits_robIdx_5_value = io_commits_robIdx_5_value;
        //    mon_tr.io_commits_robIdx_6_flag = io_commits_robIdx_6_flag;
        //    mon_tr.io_commits_robIdx_6_value = io_commits_robIdx_6_value;
        //    mon_tr.io_commits_robIdx_7_flag = io_commits_robIdx_7_flag;
        //    mon_tr.io_commits_robIdx_7_value = io_commits_robIdx_7_value;
        //    mon_tr.io_trace_blockCommit = io_trace_blockCommit;
        //    mon_tr.io_trace_traceCommitInfo_blocks_0_valid = io_trace_traceCommitInfo_blocks_0_valid;
        //    mon_tr.io_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value = io_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value;
        //    mon_tr.io_trace_traceCommitInfo_blocks_0_bits_ftqOffset = io_trace_traceCommitInfo_blocks_0_bits_ftqOffset;
        //    mon_tr.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype = io_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype;
        //    mon_tr.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire = io_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire;
        //    mon_tr.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize = io_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize;
        //    mon_tr.io_trace_traceCommitInfo_blocks_1_valid = io_trace_traceCommitInfo_blocks_1_valid;
        //    mon_tr.io_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value = io_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value;
        //    mon_tr.io_trace_traceCommitInfo_blocks_1_bits_ftqOffset = io_trace_traceCommitInfo_blocks_1_bits_ftqOffset;
        //    mon_tr.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype = io_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype;
        //    mon_tr.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire = io_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire;
        //    mon_tr.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize = io_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize;
        //    mon_tr.io_trace_traceCommitInfo_blocks_2_valid = io_trace_traceCommitInfo_blocks_2_valid;
        //    mon_tr.io_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value = io_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value;
        //    mon_tr.io_trace_traceCommitInfo_blocks_2_bits_ftqOffset = io_trace_traceCommitInfo_blocks_2_bits_ftqOffset;
        //    mon_tr.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype = io_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype;
        //    mon_tr.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire = io_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire;
        //    mon_tr.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize = io_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize;
        //    mon_tr.io_trace_traceCommitInfo_blocks_3_valid = io_trace_traceCommitInfo_blocks_3_valid;
        //    mon_tr.io_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value = io_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value;
        //    mon_tr.io_trace_traceCommitInfo_blocks_3_bits_ftqOffset = io_trace_traceCommitInfo_blocks_3_bits_ftqOffset;
        //    mon_tr.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype = io_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype;
        //    mon_tr.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire = io_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire;
        //    mon_tr.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize = io_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize;
        //    mon_tr.io_trace_traceCommitInfo_blocks_4_valid = io_trace_traceCommitInfo_blocks_4_valid;
        //    mon_tr.io_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value = io_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value;
        //    mon_tr.io_trace_traceCommitInfo_blocks_4_bits_ftqOffset = io_trace_traceCommitInfo_blocks_4_bits_ftqOffset;
        //    mon_tr.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype = io_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype;
        //    mon_tr.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire = io_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire;
        //    mon_tr.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize = io_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize;
        //    mon_tr.io_trace_traceCommitInfo_blocks_5_valid = io_trace_traceCommitInfo_blocks_5_valid;
        //    mon_tr.io_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value = io_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value;
        //    mon_tr.io_trace_traceCommitInfo_blocks_5_bits_ftqOffset = io_trace_traceCommitInfo_blocks_5_bits_ftqOffset;
        //    mon_tr.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype = io_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype;
        //    mon_tr.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire = io_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire;
        //    mon_tr.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize = io_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize;
        //    mon_tr.io_trace_traceCommitInfo_blocks_6_valid = io_trace_traceCommitInfo_blocks_6_valid;
        //    mon_tr.io_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value = io_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value;
        //    mon_tr.io_trace_traceCommitInfo_blocks_6_bits_ftqOffset = io_trace_traceCommitInfo_blocks_6_bits_ftqOffset;
        //    mon_tr.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype = io_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype;
        //    mon_tr.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire = io_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire;
        //    mon_tr.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize = io_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize;
        //    mon_tr.io_trace_traceCommitInfo_blocks_7_valid = io_trace_traceCommitInfo_blocks_7_valid;
        //    mon_tr.io_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value = io_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value;
        //    mon_tr.io_trace_traceCommitInfo_blocks_7_bits_ftqOffset = io_trace_traceCommitInfo_blocks_7_bits_ftqOffset;
        //    mon_tr.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype = io_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype;
        //    mon_tr.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire = io_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire;
        //    mon_tr.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize = io_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize;
        //    mon_tr.io_rabCommits_isCommit = io_rabCommits_isCommit;
        //    mon_tr.io_rabCommits_commitValid_0 = io_rabCommits_commitValid_0;
        //    mon_tr.io_rabCommits_commitValid_1 = io_rabCommits_commitValid_1;
        //    mon_tr.io_rabCommits_commitValid_2 = io_rabCommits_commitValid_2;
        //    mon_tr.io_rabCommits_commitValid_3 = io_rabCommits_commitValid_3;
        //    mon_tr.io_rabCommits_commitValid_4 = io_rabCommits_commitValid_4;
        //    mon_tr.io_rabCommits_commitValid_5 = io_rabCommits_commitValid_5;
        //    mon_tr.io_rabCommits_isWalk = io_rabCommits_isWalk;
        //    mon_tr.io_rabCommits_walkValid_0 = io_rabCommits_walkValid_0;
        //    mon_tr.io_rabCommits_walkValid_1 = io_rabCommits_walkValid_1;
        //    mon_tr.io_rabCommits_walkValid_2 = io_rabCommits_walkValid_2;
        //    mon_tr.io_rabCommits_walkValid_3 = io_rabCommits_walkValid_3;
        //    mon_tr.io_rabCommits_walkValid_4 = io_rabCommits_walkValid_4;
        //    mon_tr.io_rabCommits_walkValid_5 = io_rabCommits_walkValid_5;
        //    mon_tr.io_rabCommits_info_0_ldest = io_rabCommits_info_0_ldest;
        //    mon_tr.io_rabCommits_info_0_pdest = io_rabCommits_info_0_pdest;
        //    mon_tr.io_rabCommits_info_0_rfWen = io_rabCommits_info_0_rfWen;
        //    mon_tr.io_rabCommits_info_0_fpWen = io_rabCommits_info_0_fpWen;
        //    mon_tr.io_rabCommits_info_0_vecWen = io_rabCommits_info_0_vecWen;
        //    mon_tr.io_rabCommits_info_0_v0Wen = io_rabCommits_info_0_v0Wen;
        //    mon_tr.io_rabCommits_info_0_vlWen = io_rabCommits_info_0_vlWen;
        //    mon_tr.io_rabCommits_info_0_isMove = io_rabCommits_info_0_isMove;
        //    mon_tr.io_rabCommits_info_1_ldest = io_rabCommits_info_1_ldest;
        //    mon_tr.io_rabCommits_info_1_pdest = io_rabCommits_info_1_pdest;
        //    mon_tr.io_rabCommits_info_1_rfWen = io_rabCommits_info_1_rfWen;
        //    mon_tr.io_rabCommits_info_1_fpWen = io_rabCommits_info_1_fpWen;
        //    mon_tr.io_rabCommits_info_1_vecWen = io_rabCommits_info_1_vecWen;
        //    mon_tr.io_rabCommits_info_1_v0Wen = io_rabCommits_info_1_v0Wen;
        //    mon_tr.io_rabCommits_info_1_vlWen = io_rabCommits_info_1_vlWen;
        //    mon_tr.io_rabCommits_info_1_isMove = io_rabCommits_info_1_isMove;
        //    mon_tr.io_rabCommits_info_2_ldest = io_rabCommits_info_2_ldest;
        //    mon_tr.io_rabCommits_info_2_pdest = io_rabCommits_info_2_pdest;
        //    mon_tr.io_rabCommits_info_2_rfWen = io_rabCommits_info_2_rfWen;
        //    mon_tr.io_rabCommits_info_2_fpWen = io_rabCommits_info_2_fpWen;
        //    mon_tr.io_rabCommits_info_2_vecWen = io_rabCommits_info_2_vecWen;
        //    mon_tr.io_rabCommits_info_2_v0Wen = io_rabCommits_info_2_v0Wen;
        //    mon_tr.io_rabCommits_info_2_vlWen = io_rabCommits_info_2_vlWen;
        //    mon_tr.io_rabCommits_info_2_isMove = io_rabCommits_info_2_isMove;
        //    mon_tr.io_rabCommits_info_3_ldest = io_rabCommits_info_3_ldest;
        //    mon_tr.io_rabCommits_info_3_pdest = io_rabCommits_info_3_pdest;
        //    mon_tr.io_rabCommits_info_3_rfWen = io_rabCommits_info_3_rfWen;
        //    mon_tr.io_rabCommits_info_3_fpWen = io_rabCommits_info_3_fpWen;
        //    mon_tr.io_rabCommits_info_3_vecWen = io_rabCommits_info_3_vecWen;
        //    mon_tr.io_rabCommits_info_3_v0Wen = io_rabCommits_info_3_v0Wen;
        //    mon_tr.io_rabCommits_info_3_vlWen = io_rabCommits_info_3_vlWen;
        //    mon_tr.io_rabCommits_info_3_isMove = io_rabCommits_info_3_isMove;
        //    mon_tr.io_rabCommits_info_4_ldest = io_rabCommits_info_4_ldest;
        //    mon_tr.io_rabCommits_info_4_pdest = io_rabCommits_info_4_pdest;
        //    mon_tr.io_rabCommits_info_4_rfWen = io_rabCommits_info_4_rfWen;
        //    mon_tr.io_rabCommits_info_4_fpWen = io_rabCommits_info_4_fpWen;
        //    mon_tr.io_rabCommits_info_4_vecWen = io_rabCommits_info_4_vecWen;
        //    mon_tr.io_rabCommits_info_4_v0Wen = io_rabCommits_info_4_v0Wen;
        //    mon_tr.io_rabCommits_info_4_vlWen = io_rabCommits_info_4_vlWen;
        //    mon_tr.io_rabCommits_info_4_isMove = io_rabCommits_info_4_isMove;
        //    mon_tr.io_rabCommits_info_5_ldest = io_rabCommits_info_5_ldest;
        //    mon_tr.io_rabCommits_info_5_pdest = io_rabCommits_info_5_pdest;
        //    mon_tr.io_rabCommits_info_5_rfWen = io_rabCommits_info_5_rfWen;
        //    mon_tr.io_rabCommits_info_5_fpWen = io_rabCommits_info_5_fpWen;
        //    mon_tr.io_rabCommits_info_5_vecWen = io_rabCommits_info_5_vecWen;
        //    mon_tr.io_rabCommits_info_5_v0Wen = io_rabCommits_info_5_v0Wen;
        //    mon_tr.io_rabCommits_info_5_vlWen = io_rabCommits_info_5_vlWen;
        //    mon_tr.io_rabCommits_info_5_isMove = io_rabCommits_info_5_isMove;
        //    mon_tr.io_diffCommits_commitValid_0 = io_diffCommits_commitValid_0;
        //    mon_tr.io_diffCommits_commitValid_1 = io_diffCommits_commitValid_1;
        //    mon_tr.io_diffCommits_commitValid_2 = io_diffCommits_commitValid_2;
        //    mon_tr.io_diffCommits_commitValid_3 = io_diffCommits_commitValid_3;
        //    mon_tr.io_diffCommits_commitValid_4 = io_diffCommits_commitValid_4;
        //    mon_tr.io_diffCommits_commitValid_5 = io_diffCommits_commitValid_5;
        //    mon_tr.io_diffCommits_commitValid_6 = io_diffCommits_commitValid_6;
        //    mon_tr.io_diffCommits_commitValid_7 = io_diffCommits_commitValid_7;
        //    mon_tr.io_diffCommits_commitValid_8 = io_diffCommits_commitValid_8;
        //    mon_tr.io_diffCommits_commitValid_9 = io_diffCommits_commitValid_9;
        //    mon_tr.io_diffCommits_commitValid_10 = io_diffCommits_commitValid_10;
        //    mon_tr.io_diffCommits_commitValid_11 = io_diffCommits_commitValid_11;
        //    mon_tr.io_diffCommits_commitValid_12 = io_diffCommits_commitValid_12;
        //    mon_tr.io_diffCommits_commitValid_13 = io_diffCommits_commitValid_13;
        //    mon_tr.io_diffCommits_commitValid_14 = io_diffCommits_commitValid_14;
        //    mon_tr.io_diffCommits_commitValid_15 = io_diffCommits_commitValid_15;
        //    mon_tr.io_diffCommits_commitValid_16 = io_diffCommits_commitValid_16;
        //    mon_tr.io_diffCommits_commitValid_17 = io_diffCommits_commitValid_17;
        //    mon_tr.io_diffCommits_commitValid_18 = io_diffCommits_commitValid_18;
        //    mon_tr.io_diffCommits_commitValid_19 = io_diffCommits_commitValid_19;
        //    mon_tr.io_diffCommits_commitValid_20 = io_diffCommits_commitValid_20;
        //    mon_tr.io_diffCommits_commitValid_21 = io_diffCommits_commitValid_21;
        //    mon_tr.io_diffCommits_commitValid_22 = io_diffCommits_commitValid_22;
        //    mon_tr.io_diffCommits_commitValid_23 = io_diffCommits_commitValid_23;
        //    mon_tr.io_diffCommits_commitValid_24 = io_diffCommits_commitValid_24;
        //    mon_tr.io_diffCommits_commitValid_25 = io_diffCommits_commitValid_25;
        //    mon_tr.io_diffCommits_commitValid_26 = io_diffCommits_commitValid_26;
        //    mon_tr.io_diffCommits_commitValid_27 = io_diffCommits_commitValid_27;
        //    mon_tr.io_diffCommits_commitValid_28 = io_diffCommits_commitValid_28;
        //    mon_tr.io_diffCommits_commitValid_29 = io_diffCommits_commitValid_29;
        //    mon_tr.io_diffCommits_commitValid_30 = io_diffCommits_commitValid_30;
        //    mon_tr.io_diffCommits_commitValid_31 = io_diffCommits_commitValid_31;
        //    mon_tr.io_diffCommits_commitValid_32 = io_diffCommits_commitValid_32;
        //    mon_tr.io_diffCommits_commitValid_33 = io_diffCommits_commitValid_33;
        //    mon_tr.io_diffCommits_commitValid_34 = io_diffCommits_commitValid_34;
        //    mon_tr.io_diffCommits_commitValid_35 = io_diffCommits_commitValid_35;
        //    mon_tr.io_diffCommits_commitValid_36 = io_diffCommits_commitValid_36;
        //    mon_tr.io_diffCommits_commitValid_37 = io_diffCommits_commitValid_37;
        //    mon_tr.io_diffCommits_commitValid_38 = io_diffCommits_commitValid_38;
        //    mon_tr.io_diffCommits_commitValid_39 = io_diffCommits_commitValid_39;
        //    mon_tr.io_diffCommits_commitValid_40 = io_diffCommits_commitValid_40;
        //    mon_tr.io_diffCommits_commitValid_41 = io_diffCommits_commitValid_41;
        //    mon_tr.io_diffCommits_commitValid_42 = io_diffCommits_commitValid_42;
        //    mon_tr.io_diffCommits_commitValid_43 = io_diffCommits_commitValid_43;
        //    mon_tr.io_diffCommits_commitValid_44 = io_diffCommits_commitValid_44;
        //    mon_tr.io_diffCommits_commitValid_45 = io_diffCommits_commitValid_45;
        //    mon_tr.io_diffCommits_commitValid_46 = io_diffCommits_commitValid_46;
        //    mon_tr.io_diffCommits_commitValid_47 = io_diffCommits_commitValid_47;
        //    mon_tr.io_diffCommits_commitValid_48 = io_diffCommits_commitValid_48;
        //    mon_tr.io_diffCommits_commitValid_49 = io_diffCommits_commitValid_49;
        //    mon_tr.io_diffCommits_commitValid_50 = io_diffCommits_commitValid_50;
        //    mon_tr.io_diffCommits_commitValid_51 = io_diffCommits_commitValid_51;
        //    mon_tr.io_diffCommits_commitValid_52 = io_diffCommits_commitValid_52;
        //    mon_tr.io_diffCommits_commitValid_53 = io_diffCommits_commitValid_53;
        //    mon_tr.io_diffCommits_commitValid_54 = io_diffCommits_commitValid_54;
        //    mon_tr.io_diffCommits_commitValid_55 = io_diffCommits_commitValid_55;
        //    mon_tr.io_diffCommits_commitValid_56 = io_diffCommits_commitValid_56;
        //    mon_tr.io_diffCommits_commitValid_57 = io_diffCommits_commitValid_57;
        //    mon_tr.io_diffCommits_commitValid_58 = io_diffCommits_commitValid_58;
        //    mon_tr.io_diffCommits_commitValid_59 = io_diffCommits_commitValid_59;
        //    mon_tr.io_diffCommits_commitValid_60 = io_diffCommits_commitValid_60;
        //    mon_tr.io_diffCommits_commitValid_61 = io_diffCommits_commitValid_61;
        //    mon_tr.io_diffCommits_commitValid_62 = io_diffCommits_commitValid_62;
        //    mon_tr.io_diffCommits_commitValid_63 = io_diffCommits_commitValid_63;
        //    mon_tr.io_diffCommits_commitValid_64 = io_diffCommits_commitValid_64;
        //    mon_tr.io_diffCommits_commitValid_65 = io_diffCommits_commitValid_65;
        //    mon_tr.io_diffCommits_commitValid_66 = io_diffCommits_commitValid_66;
        //    mon_tr.io_diffCommits_commitValid_67 = io_diffCommits_commitValid_67;
        //    mon_tr.io_diffCommits_commitValid_68 = io_diffCommits_commitValid_68;
        //    mon_tr.io_diffCommits_commitValid_69 = io_diffCommits_commitValid_69;
        //    mon_tr.io_diffCommits_commitValid_70 = io_diffCommits_commitValid_70;
        //    mon_tr.io_diffCommits_commitValid_71 = io_diffCommits_commitValid_71;
        //    mon_tr.io_diffCommits_commitValid_72 = io_diffCommits_commitValid_72;
        //    mon_tr.io_diffCommits_commitValid_73 = io_diffCommits_commitValid_73;
        //    mon_tr.io_diffCommits_commitValid_74 = io_diffCommits_commitValid_74;
        //    mon_tr.io_diffCommits_commitValid_75 = io_diffCommits_commitValid_75;
        //    mon_tr.io_diffCommits_commitValid_76 = io_diffCommits_commitValid_76;
        //    mon_tr.io_diffCommits_commitValid_77 = io_diffCommits_commitValid_77;
        //    mon_tr.io_diffCommits_commitValid_78 = io_diffCommits_commitValid_78;
        //    mon_tr.io_diffCommits_commitValid_79 = io_diffCommits_commitValid_79;
        //    mon_tr.io_diffCommits_commitValid_80 = io_diffCommits_commitValid_80;
        //    mon_tr.io_diffCommits_commitValid_81 = io_diffCommits_commitValid_81;
        //    mon_tr.io_diffCommits_commitValid_82 = io_diffCommits_commitValid_82;
        //    mon_tr.io_diffCommits_commitValid_83 = io_diffCommits_commitValid_83;
        //    mon_tr.io_diffCommits_commitValid_84 = io_diffCommits_commitValid_84;
        //    mon_tr.io_diffCommits_commitValid_85 = io_diffCommits_commitValid_85;
        //    mon_tr.io_diffCommits_commitValid_86 = io_diffCommits_commitValid_86;
        //    mon_tr.io_diffCommits_commitValid_87 = io_diffCommits_commitValid_87;
        //    mon_tr.io_diffCommits_commitValid_88 = io_diffCommits_commitValid_88;
        //    mon_tr.io_diffCommits_commitValid_89 = io_diffCommits_commitValid_89;
        //    mon_tr.io_diffCommits_commitValid_90 = io_diffCommits_commitValid_90;
        //    mon_tr.io_diffCommits_commitValid_91 = io_diffCommits_commitValid_91;
        //    mon_tr.io_diffCommits_commitValid_92 = io_diffCommits_commitValid_92;
        //    mon_tr.io_diffCommits_commitValid_93 = io_diffCommits_commitValid_93;
        //    mon_tr.io_diffCommits_commitValid_94 = io_diffCommits_commitValid_94;
        //    mon_tr.io_diffCommits_commitValid_95 = io_diffCommits_commitValid_95;
        //    mon_tr.io_diffCommits_commitValid_96 = io_diffCommits_commitValid_96;
        //    mon_tr.io_diffCommits_commitValid_97 = io_diffCommits_commitValid_97;
        //    mon_tr.io_diffCommits_commitValid_98 = io_diffCommits_commitValid_98;
        //    mon_tr.io_diffCommits_commitValid_99 = io_diffCommits_commitValid_99;
        //    mon_tr.io_diffCommits_commitValid_100 = io_diffCommits_commitValid_100;
        //    mon_tr.io_diffCommits_commitValid_101 = io_diffCommits_commitValid_101;
        //    mon_tr.io_diffCommits_commitValid_102 = io_diffCommits_commitValid_102;
        //    mon_tr.io_diffCommits_commitValid_103 = io_diffCommits_commitValid_103;
        //    mon_tr.io_diffCommits_commitValid_104 = io_diffCommits_commitValid_104;
        //    mon_tr.io_diffCommits_commitValid_105 = io_diffCommits_commitValid_105;
        //    mon_tr.io_diffCommits_commitValid_106 = io_diffCommits_commitValid_106;
        //    mon_tr.io_diffCommits_commitValid_107 = io_diffCommits_commitValid_107;
        //    mon_tr.io_diffCommits_commitValid_108 = io_diffCommits_commitValid_108;
        //    mon_tr.io_diffCommits_commitValid_109 = io_diffCommits_commitValid_109;
        //    mon_tr.io_diffCommits_commitValid_110 = io_diffCommits_commitValid_110;
        //    mon_tr.io_diffCommits_commitValid_111 = io_diffCommits_commitValid_111;
        //    mon_tr.io_diffCommits_commitValid_112 = io_diffCommits_commitValid_112;
        //    mon_tr.io_diffCommits_commitValid_113 = io_diffCommits_commitValid_113;
        //    mon_tr.io_diffCommits_commitValid_114 = io_diffCommits_commitValid_114;
        //    mon_tr.io_diffCommits_commitValid_115 = io_diffCommits_commitValid_115;
        //    mon_tr.io_diffCommits_commitValid_116 = io_diffCommits_commitValid_116;
        //    mon_tr.io_diffCommits_commitValid_117 = io_diffCommits_commitValid_117;
        //    mon_tr.io_diffCommits_commitValid_118 = io_diffCommits_commitValid_118;
        //    mon_tr.io_diffCommits_commitValid_119 = io_diffCommits_commitValid_119;
        //    mon_tr.io_diffCommits_commitValid_120 = io_diffCommits_commitValid_120;
        //    mon_tr.io_diffCommits_commitValid_121 = io_diffCommits_commitValid_121;
        //    mon_tr.io_diffCommits_commitValid_122 = io_diffCommits_commitValid_122;
        //    mon_tr.io_diffCommits_commitValid_123 = io_diffCommits_commitValid_123;
        //    mon_tr.io_diffCommits_commitValid_124 = io_diffCommits_commitValid_124;
        //    mon_tr.io_diffCommits_commitValid_125 = io_diffCommits_commitValid_125;
        //    mon_tr.io_diffCommits_commitValid_126 = io_diffCommits_commitValid_126;
        //    mon_tr.io_diffCommits_commitValid_127 = io_diffCommits_commitValid_127;
        //    mon_tr.io_diffCommits_commitValid_128 = io_diffCommits_commitValid_128;
        //    mon_tr.io_diffCommits_commitValid_129 = io_diffCommits_commitValid_129;
        //    mon_tr.io_diffCommits_commitValid_130 = io_diffCommits_commitValid_130;
        //    mon_tr.io_diffCommits_commitValid_131 = io_diffCommits_commitValid_131;
        //    mon_tr.io_diffCommits_commitValid_132 = io_diffCommits_commitValid_132;
        //    mon_tr.io_diffCommits_commitValid_133 = io_diffCommits_commitValid_133;
        //    mon_tr.io_diffCommits_commitValid_134 = io_diffCommits_commitValid_134;
        //    mon_tr.io_diffCommits_commitValid_135 = io_diffCommits_commitValid_135;
        //    mon_tr.io_diffCommits_commitValid_136 = io_diffCommits_commitValid_136;
        //    mon_tr.io_diffCommits_commitValid_137 = io_diffCommits_commitValid_137;
        //    mon_tr.io_diffCommits_commitValid_138 = io_diffCommits_commitValid_138;
        //    mon_tr.io_diffCommits_commitValid_139 = io_diffCommits_commitValid_139;
        //    mon_tr.io_diffCommits_commitValid_140 = io_diffCommits_commitValid_140;
        //    mon_tr.io_diffCommits_commitValid_141 = io_diffCommits_commitValid_141;
        //    mon_tr.io_diffCommits_commitValid_142 = io_diffCommits_commitValid_142;
        //    mon_tr.io_diffCommits_commitValid_143 = io_diffCommits_commitValid_143;
        //    mon_tr.io_diffCommits_commitValid_144 = io_diffCommits_commitValid_144;
        //    mon_tr.io_diffCommits_commitValid_145 = io_diffCommits_commitValid_145;
        //    mon_tr.io_diffCommits_commitValid_146 = io_diffCommits_commitValid_146;
        //    mon_tr.io_diffCommits_commitValid_147 = io_diffCommits_commitValid_147;
        //    mon_tr.io_diffCommits_commitValid_148 = io_diffCommits_commitValid_148;
        //    mon_tr.io_diffCommits_commitValid_149 = io_diffCommits_commitValid_149;
        //    mon_tr.io_diffCommits_commitValid_150 = io_diffCommits_commitValid_150;
        //    mon_tr.io_diffCommits_commitValid_151 = io_diffCommits_commitValid_151;
        //    mon_tr.io_diffCommits_commitValid_152 = io_diffCommits_commitValid_152;
        //    mon_tr.io_diffCommits_commitValid_153 = io_diffCommits_commitValid_153;
        //    mon_tr.io_diffCommits_commitValid_154 = io_diffCommits_commitValid_154;
        //    mon_tr.io_diffCommits_commitValid_155 = io_diffCommits_commitValid_155;
        //    mon_tr.io_diffCommits_commitValid_156 = io_diffCommits_commitValid_156;
        //    mon_tr.io_diffCommits_commitValid_157 = io_diffCommits_commitValid_157;
        //    mon_tr.io_diffCommits_commitValid_158 = io_diffCommits_commitValid_158;
        //    mon_tr.io_diffCommits_commitValid_159 = io_diffCommits_commitValid_159;
        //    mon_tr.io_diffCommits_commitValid_160 = io_diffCommits_commitValid_160;
        //    mon_tr.io_diffCommits_commitValid_161 = io_diffCommits_commitValid_161;
        //    mon_tr.io_diffCommits_commitValid_162 = io_diffCommits_commitValid_162;
        //    mon_tr.io_diffCommits_commitValid_163 = io_diffCommits_commitValid_163;
        //    mon_tr.io_diffCommits_commitValid_164 = io_diffCommits_commitValid_164;
        //    mon_tr.io_diffCommits_commitValid_165 = io_diffCommits_commitValid_165;
        //    mon_tr.io_diffCommits_commitValid_166 = io_diffCommits_commitValid_166;
        //    mon_tr.io_diffCommits_commitValid_167 = io_diffCommits_commitValid_167;
        //    mon_tr.io_diffCommits_commitValid_168 = io_diffCommits_commitValid_168;
        //    mon_tr.io_diffCommits_commitValid_169 = io_diffCommits_commitValid_169;
        //    mon_tr.io_diffCommits_commitValid_170 = io_diffCommits_commitValid_170;
        //    mon_tr.io_diffCommits_commitValid_171 = io_diffCommits_commitValid_171;
        //    mon_tr.io_diffCommits_commitValid_172 = io_diffCommits_commitValid_172;
        //    mon_tr.io_diffCommits_commitValid_173 = io_diffCommits_commitValid_173;
        //    mon_tr.io_diffCommits_commitValid_174 = io_diffCommits_commitValid_174;
        //    mon_tr.io_diffCommits_commitValid_175 = io_diffCommits_commitValid_175;
        //    mon_tr.io_diffCommits_commitValid_176 = io_diffCommits_commitValid_176;
        //    mon_tr.io_diffCommits_commitValid_177 = io_diffCommits_commitValid_177;
        //    mon_tr.io_diffCommits_commitValid_178 = io_diffCommits_commitValid_178;
        //    mon_tr.io_diffCommits_commitValid_179 = io_diffCommits_commitValid_179;
        //    mon_tr.io_diffCommits_commitValid_180 = io_diffCommits_commitValid_180;
        //    mon_tr.io_diffCommits_commitValid_181 = io_diffCommits_commitValid_181;
        //    mon_tr.io_diffCommits_commitValid_182 = io_diffCommits_commitValid_182;
        //    mon_tr.io_diffCommits_commitValid_183 = io_diffCommits_commitValid_183;
        //    mon_tr.io_diffCommits_commitValid_184 = io_diffCommits_commitValid_184;
        //    mon_tr.io_diffCommits_commitValid_185 = io_diffCommits_commitValid_185;
        //    mon_tr.io_diffCommits_commitValid_186 = io_diffCommits_commitValid_186;
        //    mon_tr.io_diffCommits_commitValid_187 = io_diffCommits_commitValid_187;
        //    mon_tr.io_diffCommits_commitValid_188 = io_diffCommits_commitValid_188;
        //    mon_tr.io_diffCommits_commitValid_189 = io_diffCommits_commitValid_189;
        //    mon_tr.io_diffCommits_commitValid_190 = io_diffCommits_commitValid_190;
        //    mon_tr.io_diffCommits_commitValid_191 = io_diffCommits_commitValid_191;
        //    mon_tr.io_diffCommits_commitValid_192 = io_diffCommits_commitValid_192;
        //    mon_tr.io_diffCommits_commitValid_193 = io_diffCommits_commitValid_193;
        //    mon_tr.io_diffCommits_commitValid_194 = io_diffCommits_commitValid_194;
        //    mon_tr.io_diffCommits_commitValid_195 = io_diffCommits_commitValid_195;
        //    mon_tr.io_diffCommits_commitValid_196 = io_diffCommits_commitValid_196;
        //    mon_tr.io_diffCommits_commitValid_197 = io_diffCommits_commitValid_197;
        //    mon_tr.io_diffCommits_commitValid_198 = io_diffCommits_commitValid_198;
        //    mon_tr.io_diffCommits_commitValid_199 = io_diffCommits_commitValid_199;
        //    mon_tr.io_diffCommits_commitValid_200 = io_diffCommits_commitValid_200;
        //    mon_tr.io_diffCommits_commitValid_201 = io_diffCommits_commitValid_201;
        //    mon_tr.io_diffCommits_commitValid_202 = io_diffCommits_commitValid_202;
        //    mon_tr.io_diffCommits_commitValid_203 = io_diffCommits_commitValid_203;
        //    mon_tr.io_diffCommits_commitValid_204 = io_diffCommits_commitValid_204;
        //    mon_tr.io_diffCommits_commitValid_205 = io_diffCommits_commitValid_205;
        //    mon_tr.io_diffCommits_commitValid_206 = io_diffCommits_commitValid_206;
        //    mon_tr.io_diffCommits_commitValid_207 = io_diffCommits_commitValid_207;
        //    mon_tr.io_diffCommits_commitValid_208 = io_diffCommits_commitValid_208;
        //    mon_tr.io_diffCommits_commitValid_209 = io_diffCommits_commitValid_209;
        //    mon_tr.io_diffCommits_commitValid_210 = io_diffCommits_commitValid_210;
        //    mon_tr.io_diffCommits_commitValid_211 = io_diffCommits_commitValid_211;
        //    mon_tr.io_diffCommits_commitValid_212 = io_diffCommits_commitValid_212;
        //    mon_tr.io_diffCommits_commitValid_213 = io_diffCommits_commitValid_213;
        //    mon_tr.io_diffCommits_commitValid_214 = io_diffCommits_commitValid_214;
        //    mon_tr.io_diffCommits_commitValid_215 = io_diffCommits_commitValid_215;
        //    mon_tr.io_diffCommits_commitValid_216 = io_diffCommits_commitValid_216;
        //    mon_tr.io_diffCommits_commitValid_217 = io_diffCommits_commitValid_217;
        //    mon_tr.io_diffCommits_commitValid_218 = io_diffCommits_commitValid_218;
        //    mon_tr.io_diffCommits_commitValid_219 = io_diffCommits_commitValid_219;
        //    mon_tr.io_diffCommits_commitValid_220 = io_diffCommits_commitValid_220;
        //    mon_tr.io_diffCommits_commitValid_221 = io_diffCommits_commitValid_221;
        //    mon_tr.io_diffCommits_commitValid_222 = io_diffCommits_commitValid_222;
        //    mon_tr.io_diffCommits_commitValid_223 = io_diffCommits_commitValid_223;
        //    mon_tr.io_diffCommits_commitValid_224 = io_diffCommits_commitValid_224;
        //    mon_tr.io_diffCommits_commitValid_225 = io_diffCommits_commitValid_225;
        //    mon_tr.io_diffCommits_commitValid_226 = io_diffCommits_commitValid_226;
        //    mon_tr.io_diffCommits_commitValid_227 = io_diffCommits_commitValid_227;
        //    mon_tr.io_diffCommits_commitValid_228 = io_diffCommits_commitValid_228;
        //    mon_tr.io_diffCommits_commitValid_229 = io_diffCommits_commitValid_229;
        //    mon_tr.io_diffCommits_commitValid_230 = io_diffCommits_commitValid_230;
        //    mon_tr.io_diffCommits_commitValid_231 = io_diffCommits_commitValid_231;
        //    mon_tr.io_diffCommits_commitValid_232 = io_diffCommits_commitValid_232;
        //    mon_tr.io_diffCommits_commitValid_233 = io_diffCommits_commitValid_233;
        //    mon_tr.io_diffCommits_commitValid_234 = io_diffCommits_commitValid_234;
        //    mon_tr.io_diffCommits_commitValid_235 = io_diffCommits_commitValid_235;
        //    mon_tr.io_diffCommits_commitValid_236 = io_diffCommits_commitValid_236;
        //    mon_tr.io_diffCommits_commitValid_237 = io_diffCommits_commitValid_237;
        //    mon_tr.io_diffCommits_commitValid_238 = io_diffCommits_commitValid_238;
        //    mon_tr.io_diffCommits_commitValid_239 = io_diffCommits_commitValid_239;
        //    mon_tr.io_diffCommits_commitValid_240 = io_diffCommits_commitValid_240;
        //    mon_tr.io_diffCommits_commitValid_241 = io_diffCommits_commitValid_241;
        //    mon_tr.io_diffCommits_commitValid_242 = io_diffCommits_commitValid_242;
        //    mon_tr.io_diffCommits_commitValid_243 = io_diffCommits_commitValid_243;
        //    mon_tr.io_diffCommits_commitValid_244 = io_diffCommits_commitValid_244;
        //    mon_tr.io_diffCommits_commitValid_245 = io_diffCommits_commitValid_245;
        //    mon_tr.io_diffCommits_commitValid_246 = io_diffCommits_commitValid_246;
        //    mon_tr.io_diffCommits_commitValid_247 = io_diffCommits_commitValid_247;
        //    mon_tr.io_diffCommits_commitValid_248 = io_diffCommits_commitValid_248;
        //    mon_tr.io_diffCommits_commitValid_249 = io_diffCommits_commitValid_249;
        //    mon_tr.io_diffCommits_commitValid_250 = io_diffCommits_commitValid_250;
        //    mon_tr.io_diffCommits_commitValid_251 = io_diffCommits_commitValid_251;
        //    mon_tr.io_diffCommits_commitValid_252 = io_diffCommits_commitValid_252;
        //    mon_tr.io_diffCommits_commitValid_253 = io_diffCommits_commitValid_253;
        //    mon_tr.io_diffCommits_commitValid_254 = io_diffCommits_commitValid_254;
        //    mon_tr.io_diffCommits_info_0_ldest = io_diffCommits_info_0_ldest;
        //    mon_tr.io_diffCommits_info_0_pdest = io_diffCommits_info_0_pdest;
        //    mon_tr.io_diffCommits_info_0_rfWen = io_diffCommits_info_0_rfWen;
        //    mon_tr.io_diffCommits_info_0_fpWen = io_diffCommits_info_0_fpWen;
        //    mon_tr.io_diffCommits_info_0_vecWen = io_diffCommits_info_0_vecWen;
        //    mon_tr.io_diffCommits_info_0_v0Wen = io_diffCommits_info_0_v0Wen;
        //    mon_tr.io_diffCommits_info_0_vlWen = io_diffCommits_info_0_vlWen;
        //    mon_tr.io_diffCommits_info_1_ldest = io_diffCommits_info_1_ldest;
        //    mon_tr.io_diffCommits_info_1_pdest = io_diffCommits_info_1_pdest;
        //    mon_tr.io_diffCommits_info_1_rfWen = io_diffCommits_info_1_rfWen;
        //    mon_tr.io_diffCommits_info_1_fpWen = io_diffCommits_info_1_fpWen;
        //    mon_tr.io_diffCommits_info_1_vecWen = io_diffCommits_info_1_vecWen;
        //    mon_tr.io_diffCommits_info_1_v0Wen = io_diffCommits_info_1_v0Wen;
        //    mon_tr.io_diffCommits_info_1_vlWen = io_diffCommits_info_1_vlWen;
        //    mon_tr.io_diffCommits_info_2_ldest = io_diffCommits_info_2_ldest;
        //    mon_tr.io_diffCommits_info_2_pdest = io_diffCommits_info_2_pdest;
        //    mon_tr.io_diffCommits_info_2_rfWen = io_diffCommits_info_2_rfWen;
        //    mon_tr.io_diffCommits_info_2_fpWen = io_diffCommits_info_2_fpWen;
        //    mon_tr.io_diffCommits_info_2_vecWen = io_diffCommits_info_2_vecWen;
        //    mon_tr.io_diffCommits_info_2_v0Wen = io_diffCommits_info_2_v0Wen;
        //    mon_tr.io_diffCommits_info_2_vlWen = io_diffCommits_info_2_vlWen;
        //    mon_tr.io_diffCommits_info_3_ldest = io_diffCommits_info_3_ldest;
        //    mon_tr.io_diffCommits_info_3_pdest = io_diffCommits_info_3_pdest;
        //    mon_tr.io_diffCommits_info_3_rfWen = io_diffCommits_info_3_rfWen;
        //    mon_tr.io_diffCommits_info_3_fpWen = io_diffCommits_info_3_fpWen;
        //    mon_tr.io_diffCommits_info_3_vecWen = io_diffCommits_info_3_vecWen;
        //    mon_tr.io_diffCommits_info_3_v0Wen = io_diffCommits_info_3_v0Wen;
        //    mon_tr.io_diffCommits_info_3_vlWen = io_diffCommits_info_3_vlWen;
        //    mon_tr.io_diffCommits_info_4_ldest = io_diffCommits_info_4_ldest;
        //    mon_tr.io_diffCommits_info_4_pdest = io_diffCommits_info_4_pdest;
        //    mon_tr.io_diffCommits_info_4_rfWen = io_diffCommits_info_4_rfWen;
        //    mon_tr.io_diffCommits_info_4_fpWen = io_diffCommits_info_4_fpWen;
        //    mon_tr.io_diffCommits_info_4_vecWen = io_diffCommits_info_4_vecWen;
        //    mon_tr.io_diffCommits_info_4_v0Wen = io_diffCommits_info_4_v0Wen;
        //    mon_tr.io_diffCommits_info_4_vlWen = io_diffCommits_info_4_vlWen;
        //    mon_tr.io_diffCommits_info_5_ldest = io_diffCommits_info_5_ldest;
        //    mon_tr.io_diffCommits_info_5_pdest = io_diffCommits_info_5_pdest;
        //    mon_tr.io_diffCommits_info_5_rfWen = io_diffCommits_info_5_rfWen;
        //    mon_tr.io_diffCommits_info_5_fpWen = io_diffCommits_info_5_fpWen;
        //    mon_tr.io_diffCommits_info_5_vecWen = io_diffCommits_info_5_vecWen;
        //    mon_tr.io_diffCommits_info_5_v0Wen = io_diffCommits_info_5_v0Wen;
        //    mon_tr.io_diffCommits_info_5_vlWen = io_diffCommits_info_5_vlWen;
        //    mon_tr.io_diffCommits_info_6_ldest = io_diffCommits_info_6_ldest;
        //    mon_tr.io_diffCommits_info_6_pdest = io_diffCommits_info_6_pdest;
        //    mon_tr.io_diffCommits_info_6_rfWen = io_diffCommits_info_6_rfWen;
        //    mon_tr.io_diffCommits_info_6_fpWen = io_diffCommits_info_6_fpWen;
        //    mon_tr.io_diffCommits_info_6_vecWen = io_diffCommits_info_6_vecWen;
        //    mon_tr.io_diffCommits_info_6_v0Wen = io_diffCommits_info_6_v0Wen;
        //    mon_tr.io_diffCommits_info_6_vlWen = io_diffCommits_info_6_vlWen;
        //    mon_tr.io_diffCommits_info_7_ldest = io_diffCommits_info_7_ldest;
        //    mon_tr.io_diffCommits_info_7_pdest = io_diffCommits_info_7_pdest;
        //    mon_tr.io_diffCommits_info_7_rfWen = io_diffCommits_info_7_rfWen;
        //    mon_tr.io_diffCommits_info_7_fpWen = io_diffCommits_info_7_fpWen;
        //    mon_tr.io_diffCommits_info_7_vecWen = io_diffCommits_info_7_vecWen;
        //    mon_tr.io_diffCommits_info_7_v0Wen = io_diffCommits_info_7_v0Wen;
        //    mon_tr.io_diffCommits_info_7_vlWen = io_diffCommits_info_7_vlWen;
        //    mon_tr.io_diffCommits_info_8_ldest = io_diffCommits_info_8_ldest;
        //    mon_tr.io_diffCommits_info_8_pdest = io_diffCommits_info_8_pdest;
        //    mon_tr.io_diffCommits_info_8_rfWen = io_diffCommits_info_8_rfWen;
        //    mon_tr.io_diffCommits_info_8_fpWen = io_diffCommits_info_8_fpWen;
        //    mon_tr.io_diffCommits_info_8_vecWen = io_diffCommits_info_8_vecWen;
        //    mon_tr.io_diffCommits_info_8_v0Wen = io_diffCommits_info_8_v0Wen;
        //    mon_tr.io_diffCommits_info_8_vlWen = io_diffCommits_info_8_vlWen;
        //    mon_tr.io_diffCommits_info_9_ldest = io_diffCommits_info_9_ldest;
        //    mon_tr.io_diffCommits_info_9_pdest = io_diffCommits_info_9_pdest;
        //    mon_tr.io_diffCommits_info_9_rfWen = io_diffCommits_info_9_rfWen;
        //    mon_tr.io_diffCommits_info_9_fpWen = io_diffCommits_info_9_fpWen;
        //    mon_tr.io_diffCommits_info_9_vecWen = io_diffCommits_info_9_vecWen;
        //    mon_tr.io_diffCommits_info_9_v0Wen = io_diffCommits_info_9_v0Wen;
        //    mon_tr.io_diffCommits_info_9_vlWen = io_diffCommits_info_9_vlWen;
        //    mon_tr.io_diffCommits_info_10_ldest = io_diffCommits_info_10_ldest;
        //    mon_tr.io_diffCommits_info_10_pdest = io_diffCommits_info_10_pdest;
        //    mon_tr.io_diffCommits_info_10_rfWen = io_diffCommits_info_10_rfWen;
        //    mon_tr.io_diffCommits_info_10_fpWen = io_diffCommits_info_10_fpWen;
        //    mon_tr.io_diffCommits_info_10_vecWen = io_diffCommits_info_10_vecWen;
        //    mon_tr.io_diffCommits_info_10_v0Wen = io_diffCommits_info_10_v0Wen;
        //    mon_tr.io_diffCommits_info_10_vlWen = io_diffCommits_info_10_vlWen;
        //    mon_tr.io_diffCommits_info_11_ldest = io_diffCommits_info_11_ldest;
        //    mon_tr.io_diffCommits_info_11_pdest = io_diffCommits_info_11_pdest;
        //    mon_tr.io_diffCommits_info_11_rfWen = io_diffCommits_info_11_rfWen;
        //    mon_tr.io_diffCommits_info_11_fpWen = io_diffCommits_info_11_fpWen;
        //    mon_tr.io_diffCommits_info_11_vecWen = io_diffCommits_info_11_vecWen;
        //    mon_tr.io_diffCommits_info_11_v0Wen = io_diffCommits_info_11_v0Wen;
        //    mon_tr.io_diffCommits_info_11_vlWen = io_diffCommits_info_11_vlWen;
        //    mon_tr.io_diffCommits_info_12_ldest = io_diffCommits_info_12_ldest;
        //    mon_tr.io_diffCommits_info_12_pdest = io_diffCommits_info_12_pdest;
        //    mon_tr.io_diffCommits_info_12_rfWen = io_diffCommits_info_12_rfWen;
        //    mon_tr.io_diffCommits_info_12_fpWen = io_diffCommits_info_12_fpWen;
        //    mon_tr.io_diffCommits_info_12_vecWen = io_diffCommits_info_12_vecWen;
        //    mon_tr.io_diffCommits_info_12_v0Wen = io_diffCommits_info_12_v0Wen;
        //    mon_tr.io_diffCommits_info_12_vlWen = io_diffCommits_info_12_vlWen;
        //    mon_tr.io_diffCommits_info_13_ldest = io_diffCommits_info_13_ldest;
        //    mon_tr.io_diffCommits_info_13_pdest = io_diffCommits_info_13_pdest;
        //    mon_tr.io_diffCommits_info_13_rfWen = io_diffCommits_info_13_rfWen;
        //    mon_tr.io_diffCommits_info_13_fpWen = io_diffCommits_info_13_fpWen;
        //    mon_tr.io_diffCommits_info_13_vecWen = io_diffCommits_info_13_vecWen;
        //    mon_tr.io_diffCommits_info_13_v0Wen = io_diffCommits_info_13_v0Wen;
        //    mon_tr.io_diffCommits_info_13_vlWen = io_diffCommits_info_13_vlWen;
        //    mon_tr.io_diffCommits_info_14_ldest = io_diffCommits_info_14_ldest;
        //    mon_tr.io_diffCommits_info_14_pdest = io_diffCommits_info_14_pdest;
        //    mon_tr.io_diffCommits_info_14_rfWen = io_diffCommits_info_14_rfWen;
        //    mon_tr.io_diffCommits_info_14_fpWen = io_diffCommits_info_14_fpWen;
        //    mon_tr.io_diffCommits_info_14_vecWen = io_diffCommits_info_14_vecWen;
        //    mon_tr.io_diffCommits_info_14_v0Wen = io_diffCommits_info_14_v0Wen;
        //    mon_tr.io_diffCommits_info_14_vlWen = io_diffCommits_info_14_vlWen;
        //    mon_tr.io_diffCommits_info_15_ldest = io_diffCommits_info_15_ldest;
        //    mon_tr.io_diffCommits_info_15_pdest = io_diffCommits_info_15_pdest;
        //    mon_tr.io_diffCommits_info_15_rfWen = io_diffCommits_info_15_rfWen;
        //    mon_tr.io_diffCommits_info_15_fpWen = io_diffCommits_info_15_fpWen;
        //    mon_tr.io_diffCommits_info_15_vecWen = io_diffCommits_info_15_vecWen;
        //    mon_tr.io_diffCommits_info_15_v0Wen = io_diffCommits_info_15_v0Wen;
        //    mon_tr.io_diffCommits_info_15_vlWen = io_diffCommits_info_15_vlWen;
        //    mon_tr.io_diffCommits_info_16_ldest = io_diffCommits_info_16_ldest;
        //    mon_tr.io_diffCommits_info_16_pdest = io_diffCommits_info_16_pdest;
        //    mon_tr.io_diffCommits_info_16_rfWen = io_diffCommits_info_16_rfWen;
        //    mon_tr.io_diffCommits_info_16_fpWen = io_diffCommits_info_16_fpWen;
        //    mon_tr.io_diffCommits_info_16_vecWen = io_diffCommits_info_16_vecWen;
        //    mon_tr.io_diffCommits_info_16_v0Wen = io_diffCommits_info_16_v0Wen;
        //    mon_tr.io_diffCommits_info_16_vlWen = io_diffCommits_info_16_vlWen;
        //    mon_tr.io_diffCommits_info_17_ldest = io_diffCommits_info_17_ldest;
        //    mon_tr.io_diffCommits_info_17_pdest = io_diffCommits_info_17_pdest;
        //    mon_tr.io_diffCommits_info_17_rfWen = io_diffCommits_info_17_rfWen;
        //    mon_tr.io_diffCommits_info_17_fpWen = io_diffCommits_info_17_fpWen;
        //    mon_tr.io_diffCommits_info_17_vecWen = io_diffCommits_info_17_vecWen;
        //    mon_tr.io_diffCommits_info_17_v0Wen = io_diffCommits_info_17_v0Wen;
        //    mon_tr.io_diffCommits_info_17_vlWen = io_diffCommits_info_17_vlWen;
        //    mon_tr.io_diffCommits_info_18_ldest = io_diffCommits_info_18_ldest;
        //    mon_tr.io_diffCommits_info_18_pdest = io_diffCommits_info_18_pdest;
        //    mon_tr.io_diffCommits_info_18_rfWen = io_diffCommits_info_18_rfWen;
        //    mon_tr.io_diffCommits_info_18_fpWen = io_diffCommits_info_18_fpWen;
        //    mon_tr.io_diffCommits_info_18_vecWen = io_diffCommits_info_18_vecWen;
        //    mon_tr.io_diffCommits_info_18_v0Wen = io_diffCommits_info_18_v0Wen;
        //    mon_tr.io_diffCommits_info_18_vlWen = io_diffCommits_info_18_vlWen;
        //    mon_tr.io_diffCommits_info_19_ldest = io_diffCommits_info_19_ldest;
        //    mon_tr.io_diffCommits_info_19_pdest = io_diffCommits_info_19_pdest;
        //    mon_tr.io_diffCommits_info_19_rfWen = io_diffCommits_info_19_rfWen;
        //    mon_tr.io_diffCommits_info_19_fpWen = io_diffCommits_info_19_fpWen;
        //    mon_tr.io_diffCommits_info_19_vecWen = io_diffCommits_info_19_vecWen;
        //    mon_tr.io_diffCommits_info_19_v0Wen = io_diffCommits_info_19_v0Wen;
        //    mon_tr.io_diffCommits_info_19_vlWen = io_diffCommits_info_19_vlWen;
        //    mon_tr.io_diffCommits_info_20_ldest = io_diffCommits_info_20_ldest;
        //    mon_tr.io_diffCommits_info_20_pdest = io_diffCommits_info_20_pdest;
        //    mon_tr.io_diffCommits_info_20_rfWen = io_diffCommits_info_20_rfWen;
        //    mon_tr.io_diffCommits_info_20_fpWen = io_diffCommits_info_20_fpWen;
        //    mon_tr.io_diffCommits_info_20_vecWen = io_diffCommits_info_20_vecWen;
        //    mon_tr.io_diffCommits_info_20_v0Wen = io_diffCommits_info_20_v0Wen;
        //    mon_tr.io_diffCommits_info_20_vlWen = io_diffCommits_info_20_vlWen;
        //    mon_tr.io_diffCommits_info_21_ldest = io_diffCommits_info_21_ldest;
        //    mon_tr.io_diffCommits_info_21_pdest = io_diffCommits_info_21_pdest;
        //    mon_tr.io_diffCommits_info_21_rfWen = io_diffCommits_info_21_rfWen;
        //    mon_tr.io_diffCommits_info_21_fpWen = io_diffCommits_info_21_fpWen;
        //    mon_tr.io_diffCommits_info_21_vecWen = io_diffCommits_info_21_vecWen;
        //    mon_tr.io_diffCommits_info_21_v0Wen = io_diffCommits_info_21_v0Wen;
        //    mon_tr.io_diffCommits_info_21_vlWen = io_diffCommits_info_21_vlWen;
        //    mon_tr.io_diffCommits_info_22_ldest = io_diffCommits_info_22_ldest;
        //    mon_tr.io_diffCommits_info_22_pdest = io_diffCommits_info_22_pdest;
        //    mon_tr.io_diffCommits_info_22_rfWen = io_diffCommits_info_22_rfWen;
        //    mon_tr.io_diffCommits_info_22_fpWen = io_diffCommits_info_22_fpWen;
        //    mon_tr.io_diffCommits_info_22_vecWen = io_diffCommits_info_22_vecWen;
        //    mon_tr.io_diffCommits_info_22_v0Wen = io_diffCommits_info_22_v0Wen;
        //    mon_tr.io_diffCommits_info_22_vlWen = io_diffCommits_info_22_vlWen;
        //    mon_tr.io_diffCommits_info_23_ldest = io_diffCommits_info_23_ldest;
        //    mon_tr.io_diffCommits_info_23_pdest = io_diffCommits_info_23_pdest;
        //    mon_tr.io_diffCommits_info_23_rfWen = io_diffCommits_info_23_rfWen;
        //    mon_tr.io_diffCommits_info_23_fpWen = io_diffCommits_info_23_fpWen;
        //    mon_tr.io_diffCommits_info_23_vecWen = io_diffCommits_info_23_vecWen;
        //    mon_tr.io_diffCommits_info_23_v0Wen = io_diffCommits_info_23_v0Wen;
        //    mon_tr.io_diffCommits_info_23_vlWen = io_diffCommits_info_23_vlWen;
        //    mon_tr.io_diffCommits_info_24_ldest = io_diffCommits_info_24_ldest;
        //    mon_tr.io_diffCommits_info_24_pdest = io_diffCommits_info_24_pdest;
        //    mon_tr.io_diffCommits_info_24_rfWen = io_diffCommits_info_24_rfWen;
        //    mon_tr.io_diffCommits_info_24_fpWen = io_diffCommits_info_24_fpWen;
        //    mon_tr.io_diffCommits_info_24_vecWen = io_diffCommits_info_24_vecWen;
        //    mon_tr.io_diffCommits_info_24_v0Wen = io_diffCommits_info_24_v0Wen;
        //    mon_tr.io_diffCommits_info_24_vlWen = io_diffCommits_info_24_vlWen;
        //    mon_tr.io_diffCommits_info_25_ldest = io_diffCommits_info_25_ldest;
        //    mon_tr.io_diffCommits_info_25_pdest = io_diffCommits_info_25_pdest;
        //    mon_tr.io_diffCommits_info_25_rfWen = io_diffCommits_info_25_rfWen;
        //    mon_tr.io_diffCommits_info_25_fpWen = io_diffCommits_info_25_fpWen;
        //    mon_tr.io_diffCommits_info_25_vecWen = io_diffCommits_info_25_vecWen;
        //    mon_tr.io_diffCommits_info_25_v0Wen = io_diffCommits_info_25_v0Wen;
        //    mon_tr.io_diffCommits_info_25_vlWen = io_diffCommits_info_25_vlWen;
        //    mon_tr.io_diffCommits_info_26_ldest = io_diffCommits_info_26_ldest;
        //    mon_tr.io_diffCommits_info_26_pdest = io_diffCommits_info_26_pdest;
        //    mon_tr.io_diffCommits_info_26_rfWen = io_diffCommits_info_26_rfWen;
        //    mon_tr.io_diffCommits_info_26_fpWen = io_diffCommits_info_26_fpWen;
        //    mon_tr.io_diffCommits_info_26_vecWen = io_diffCommits_info_26_vecWen;
        //    mon_tr.io_diffCommits_info_26_v0Wen = io_diffCommits_info_26_v0Wen;
        //    mon_tr.io_diffCommits_info_26_vlWen = io_diffCommits_info_26_vlWen;
        //    mon_tr.io_diffCommits_info_27_ldest = io_diffCommits_info_27_ldest;
        //    mon_tr.io_diffCommits_info_27_pdest = io_diffCommits_info_27_pdest;
        //    mon_tr.io_diffCommits_info_27_rfWen = io_diffCommits_info_27_rfWen;
        //    mon_tr.io_diffCommits_info_27_fpWen = io_diffCommits_info_27_fpWen;
        //    mon_tr.io_diffCommits_info_27_vecWen = io_diffCommits_info_27_vecWen;
        //    mon_tr.io_diffCommits_info_27_v0Wen = io_diffCommits_info_27_v0Wen;
        //    mon_tr.io_diffCommits_info_27_vlWen = io_diffCommits_info_27_vlWen;
        //    mon_tr.io_diffCommits_info_28_ldest = io_diffCommits_info_28_ldest;
        //    mon_tr.io_diffCommits_info_28_pdest = io_diffCommits_info_28_pdest;
        //    mon_tr.io_diffCommits_info_28_rfWen = io_diffCommits_info_28_rfWen;
        //    mon_tr.io_diffCommits_info_28_fpWen = io_diffCommits_info_28_fpWen;
        //    mon_tr.io_diffCommits_info_28_vecWen = io_diffCommits_info_28_vecWen;
        //    mon_tr.io_diffCommits_info_28_v0Wen = io_diffCommits_info_28_v0Wen;
        //    mon_tr.io_diffCommits_info_28_vlWen = io_diffCommits_info_28_vlWen;
        //    mon_tr.io_diffCommits_info_29_ldest = io_diffCommits_info_29_ldest;
        //    mon_tr.io_diffCommits_info_29_pdest = io_diffCommits_info_29_pdest;
        //    mon_tr.io_diffCommits_info_29_rfWen = io_diffCommits_info_29_rfWen;
        //    mon_tr.io_diffCommits_info_29_fpWen = io_diffCommits_info_29_fpWen;
        //    mon_tr.io_diffCommits_info_29_vecWen = io_diffCommits_info_29_vecWen;
        //    mon_tr.io_diffCommits_info_29_v0Wen = io_diffCommits_info_29_v0Wen;
        //    mon_tr.io_diffCommits_info_29_vlWen = io_diffCommits_info_29_vlWen;
        //    mon_tr.io_diffCommits_info_30_ldest = io_diffCommits_info_30_ldest;
        //    mon_tr.io_diffCommits_info_30_pdest = io_diffCommits_info_30_pdest;
        //    mon_tr.io_diffCommits_info_30_rfWen = io_diffCommits_info_30_rfWen;
        //    mon_tr.io_diffCommits_info_30_fpWen = io_diffCommits_info_30_fpWen;
        //    mon_tr.io_diffCommits_info_30_vecWen = io_diffCommits_info_30_vecWen;
        //    mon_tr.io_diffCommits_info_30_v0Wen = io_diffCommits_info_30_v0Wen;
        //    mon_tr.io_diffCommits_info_30_vlWen = io_diffCommits_info_30_vlWen;
        //    mon_tr.io_diffCommits_info_31_ldest = io_diffCommits_info_31_ldest;
        //    mon_tr.io_diffCommits_info_31_pdest = io_diffCommits_info_31_pdest;
        //    mon_tr.io_diffCommits_info_31_rfWen = io_diffCommits_info_31_rfWen;
        //    mon_tr.io_diffCommits_info_31_fpWen = io_diffCommits_info_31_fpWen;
        //    mon_tr.io_diffCommits_info_31_vecWen = io_diffCommits_info_31_vecWen;
        //    mon_tr.io_diffCommits_info_31_v0Wen = io_diffCommits_info_31_v0Wen;
        //    mon_tr.io_diffCommits_info_31_vlWen = io_diffCommits_info_31_vlWen;
        //    mon_tr.io_diffCommits_info_32_ldest = io_diffCommits_info_32_ldest;
        //    mon_tr.io_diffCommits_info_32_pdest = io_diffCommits_info_32_pdest;
        //    mon_tr.io_diffCommits_info_32_rfWen = io_diffCommits_info_32_rfWen;
        //    mon_tr.io_diffCommits_info_32_fpWen = io_diffCommits_info_32_fpWen;
        //    mon_tr.io_diffCommits_info_32_vecWen = io_diffCommits_info_32_vecWen;
        //    mon_tr.io_diffCommits_info_32_v0Wen = io_diffCommits_info_32_v0Wen;
        //    mon_tr.io_diffCommits_info_32_vlWen = io_diffCommits_info_32_vlWen;
        //    mon_tr.io_diffCommits_info_33_ldest = io_diffCommits_info_33_ldest;
        //    mon_tr.io_diffCommits_info_33_pdest = io_diffCommits_info_33_pdest;
        //    mon_tr.io_diffCommits_info_33_rfWen = io_diffCommits_info_33_rfWen;
        //    mon_tr.io_diffCommits_info_33_fpWen = io_diffCommits_info_33_fpWen;
        //    mon_tr.io_diffCommits_info_33_vecWen = io_diffCommits_info_33_vecWen;
        //    mon_tr.io_diffCommits_info_33_v0Wen = io_diffCommits_info_33_v0Wen;
        //    mon_tr.io_diffCommits_info_33_vlWen = io_diffCommits_info_33_vlWen;
        //    mon_tr.io_diffCommits_info_34_ldest = io_diffCommits_info_34_ldest;
        //    mon_tr.io_diffCommits_info_34_pdest = io_diffCommits_info_34_pdest;
        //    mon_tr.io_diffCommits_info_34_rfWen = io_diffCommits_info_34_rfWen;
        //    mon_tr.io_diffCommits_info_34_fpWen = io_diffCommits_info_34_fpWen;
        //    mon_tr.io_diffCommits_info_34_vecWen = io_diffCommits_info_34_vecWen;
        //    mon_tr.io_diffCommits_info_34_v0Wen = io_diffCommits_info_34_v0Wen;
        //    mon_tr.io_diffCommits_info_34_vlWen = io_diffCommits_info_34_vlWen;
        //    mon_tr.io_diffCommits_info_35_ldest = io_diffCommits_info_35_ldest;
        //    mon_tr.io_diffCommits_info_35_pdest = io_diffCommits_info_35_pdest;
        //    mon_tr.io_diffCommits_info_35_rfWen = io_diffCommits_info_35_rfWen;
        //    mon_tr.io_diffCommits_info_35_fpWen = io_diffCommits_info_35_fpWen;
        //    mon_tr.io_diffCommits_info_35_vecWen = io_diffCommits_info_35_vecWen;
        //    mon_tr.io_diffCommits_info_35_v0Wen = io_diffCommits_info_35_v0Wen;
        //    mon_tr.io_diffCommits_info_35_vlWen = io_diffCommits_info_35_vlWen;
        //    mon_tr.io_diffCommits_info_36_ldest = io_diffCommits_info_36_ldest;
        //    mon_tr.io_diffCommits_info_36_pdest = io_diffCommits_info_36_pdest;
        //    mon_tr.io_diffCommits_info_36_rfWen = io_diffCommits_info_36_rfWen;
        //    mon_tr.io_diffCommits_info_36_fpWen = io_diffCommits_info_36_fpWen;
        //    mon_tr.io_diffCommits_info_36_vecWen = io_diffCommits_info_36_vecWen;
        //    mon_tr.io_diffCommits_info_36_v0Wen = io_diffCommits_info_36_v0Wen;
        //    mon_tr.io_diffCommits_info_36_vlWen = io_diffCommits_info_36_vlWen;
        //    mon_tr.io_diffCommits_info_37_ldest = io_diffCommits_info_37_ldest;
        //    mon_tr.io_diffCommits_info_37_pdest = io_diffCommits_info_37_pdest;
        //    mon_tr.io_diffCommits_info_37_rfWen = io_diffCommits_info_37_rfWen;
        //    mon_tr.io_diffCommits_info_37_fpWen = io_diffCommits_info_37_fpWen;
        //    mon_tr.io_diffCommits_info_37_vecWen = io_diffCommits_info_37_vecWen;
        //    mon_tr.io_diffCommits_info_37_v0Wen = io_diffCommits_info_37_v0Wen;
        //    mon_tr.io_diffCommits_info_37_vlWen = io_diffCommits_info_37_vlWen;
        //    mon_tr.io_diffCommits_info_38_ldest = io_diffCommits_info_38_ldest;
        //    mon_tr.io_diffCommits_info_38_pdest = io_diffCommits_info_38_pdest;
        //    mon_tr.io_diffCommits_info_38_rfWen = io_diffCommits_info_38_rfWen;
        //    mon_tr.io_diffCommits_info_38_fpWen = io_diffCommits_info_38_fpWen;
        //    mon_tr.io_diffCommits_info_38_vecWen = io_diffCommits_info_38_vecWen;
        //    mon_tr.io_diffCommits_info_38_v0Wen = io_diffCommits_info_38_v0Wen;
        //    mon_tr.io_diffCommits_info_38_vlWen = io_diffCommits_info_38_vlWen;
        //    mon_tr.io_diffCommits_info_39_ldest = io_diffCommits_info_39_ldest;
        //    mon_tr.io_diffCommits_info_39_pdest = io_diffCommits_info_39_pdest;
        //    mon_tr.io_diffCommits_info_39_rfWen = io_diffCommits_info_39_rfWen;
        //    mon_tr.io_diffCommits_info_39_fpWen = io_diffCommits_info_39_fpWen;
        //    mon_tr.io_diffCommits_info_39_vecWen = io_diffCommits_info_39_vecWen;
        //    mon_tr.io_diffCommits_info_39_v0Wen = io_diffCommits_info_39_v0Wen;
        //    mon_tr.io_diffCommits_info_39_vlWen = io_diffCommits_info_39_vlWen;
        //    mon_tr.io_diffCommits_info_40_ldest = io_diffCommits_info_40_ldest;
        //    mon_tr.io_diffCommits_info_40_pdest = io_diffCommits_info_40_pdest;
        //    mon_tr.io_diffCommits_info_40_rfWen = io_diffCommits_info_40_rfWen;
        //    mon_tr.io_diffCommits_info_40_fpWen = io_diffCommits_info_40_fpWen;
        //    mon_tr.io_diffCommits_info_40_vecWen = io_diffCommits_info_40_vecWen;
        //    mon_tr.io_diffCommits_info_40_v0Wen = io_diffCommits_info_40_v0Wen;
        //    mon_tr.io_diffCommits_info_40_vlWen = io_diffCommits_info_40_vlWen;
        //    mon_tr.io_diffCommits_info_41_ldest = io_diffCommits_info_41_ldest;
        //    mon_tr.io_diffCommits_info_41_pdest = io_diffCommits_info_41_pdest;
        //    mon_tr.io_diffCommits_info_41_rfWen = io_diffCommits_info_41_rfWen;
        //    mon_tr.io_diffCommits_info_41_fpWen = io_diffCommits_info_41_fpWen;
        //    mon_tr.io_diffCommits_info_41_vecWen = io_diffCommits_info_41_vecWen;
        //    mon_tr.io_diffCommits_info_41_v0Wen = io_diffCommits_info_41_v0Wen;
        //    mon_tr.io_diffCommits_info_41_vlWen = io_diffCommits_info_41_vlWen;
        //    mon_tr.io_diffCommits_info_42_ldest = io_diffCommits_info_42_ldest;
        //    mon_tr.io_diffCommits_info_42_pdest = io_diffCommits_info_42_pdest;
        //    mon_tr.io_diffCommits_info_42_rfWen = io_diffCommits_info_42_rfWen;
        //    mon_tr.io_diffCommits_info_42_fpWen = io_diffCommits_info_42_fpWen;
        //    mon_tr.io_diffCommits_info_42_vecWen = io_diffCommits_info_42_vecWen;
        //    mon_tr.io_diffCommits_info_42_v0Wen = io_diffCommits_info_42_v0Wen;
        //    mon_tr.io_diffCommits_info_42_vlWen = io_diffCommits_info_42_vlWen;
        //    mon_tr.io_diffCommits_info_43_ldest = io_diffCommits_info_43_ldest;
        //    mon_tr.io_diffCommits_info_43_pdest = io_diffCommits_info_43_pdest;
        //    mon_tr.io_diffCommits_info_43_rfWen = io_diffCommits_info_43_rfWen;
        //    mon_tr.io_diffCommits_info_43_fpWen = io_diffCommits_info_43_fpWen;
        //    mon_tr.io_diffCommits_info_43_vecWen = io_diffCommits_info_43_vecWen;
        //    mon_tr.io_diffCommits_info_43_v0Wen = io_diffCommits_info_43_v0Wen;
        //    mon_tr.io_diffCommits_info_43_vlWen = io_diffCommits_info_43_vlWen;
        //    mon_tr.io_diffCommits_info_44_ldest = io_diffCommits_info_44_ldest;
        //    mon_tr.io_diffCommits_info_44_pdest = io_diffCommits_info_44_pdest;
        //    mon_tr.io_diffCommits_info_44_rfWen = io_diffCommits_info_44_rfWen;
        //    mon_tr.io_diffCommits_info_44_fpWen = io_diffCommits_info_44_fpWen;
        //    mon_tr.io_diffCommits_info_44_vecWen = io_diffCommits_info_44_vecWen;
        //    mon_tr.io_diffCommits_info_44_v0Wen = io_diffCommits_info_44_v0Wen;
        //    mon_tr.io_diffCommits_info_44_vlWen = io_diffCommits_info_44_vlWen;
        //    mon_tr.io_diffCommits_info_45_ldest = io_diffCommits_info_45_ldest;
        //    mon_tr.io_diffCommits_info_45_pdest = io_diffCommits_info_45_pdest;
        //    mon_tr.io_diffCommits_info_45_rfWen = io_diffCommits_info_45_rfWen;
        //    mon_tr.io_diffCommits_info_45_fpWen = io_diffCommits_info_45_fpWen;
        //    mon_tr.io_diffCommits_info_45_vecWen = io_diffCommits_info_45_vecWen;
        //    mon_tr.io_diffCommits_info_45_v0Wen = io_diffCommits_info_45_v0Wen;
        //    mon_tr.io_diffCommits_info_45_vlWen = io_diffCommits_info_45_vlWen;
        //    mon_tr.io_diffCommits_info_46_ldest = io_diffCommits_info_46_ldest;
        //    mon_tr.io_diffCommits_info_46_pdest = io_diffCommits_info_46_pdest;
        //    mon_tr.io_diffCommits_info_46_rfWen = io_diffCommits_info_46_rfWen;
        //    mon_tr.io_diffCommits_info_46_fpWen = io_diffCommits_info_46_fpWen;
        //    mon_tr.io_diffCommits_info_46_vecWen = io_diffCommits_info_46_vecWen;
        //    mon_tr.io_diffCommits_info_46_v0Wen = io_diffCommits_info_46_v0Wen;
        //    mon_tr.io_diffCommits_info_46_vlWen = io_diffCommits_info_46_vlWen;
        //    mon_tr.io_diffCommits_info_47_ldest = io_diffCommits_info_47_ldest;
        //    mon_tr.io_diffCommits_info_47_pdest = io_diffCommits_info_47_pdest;
        //    mon_tr.io_diffCommits_info_47_rfWen = io_diffCommits_info_47_rfWen;
        //    mon_tr.io_diffCommits_info_47_fpWen = io_diffCommits_info_47_fpWen;
        //    mon_tr.io_diffCommits_info_47_vecWen = io_diffCommits_info_47_vecWen;
        //    mon_tr.io_diffCommits_info_47_v0Wen = io_diffCommits_info_47_v0Wen;
        //    mon_tr.io_diffCommits_info_47_vlWen = io_diffCommits_info_47_vlWen;
        //    mon_tr.io_diffCommits_info_48_ldest = io_diffCommits_info_48_ldest;
        //    mon_tr.io_diffCommits_info_48_pdest = io_diffCommits_info_48_pdest;
        //    mon_tr.io_diffCommits_info_48_rfWen = io_diffCommits_info_48_rfWen;
        //    mon_tr.io_diffCommits_info_48_fpWen = io_diffCommits_info_48_fpWen;
        //    mon_tr.io_diffCommits_info_48_vecWen = io_diffCommits_info_48_vecWen;
        //    mon_tr.io_diffCommits_info_48_v0Wen = io_diffCommits_info_48_v0Wen;
        //    mon_tr.io_diffCommits_info_48_vlWen = io_diffCommits_info_48_vlWen;
        //    mon_tr.io_diffCommits_info_49_ldest = io_diffCommits_info_49_ldest;
        //    mon_tr.io_diffCommits_info_49_pdest = io_diffCommits_info_49_pdest;
        //    mon_tr.io_diffCommits_info_49_rfWen = io_diffCommits_info_49_rfWen;
        //    mon_tr.io_diffCommits_info_49_fpWen = io_diffCommits_info_49_fpWen;
        //    mon_tr.io_diffCommits_info_49_vecWen = io_diffCommits_info_49_vecWen;
        //    mon_tr.io_diffCommits_info_49_v0Wen = io_diffCommits_info_49_v0Wen;
        //    mon_tr.io_diffCommits_info_49_vlWen = io_diffCommits_info_49_vlWen;
        //    mon_tr.io_diffCommits_info_50_ldest = io_diffCommits_info_50_ldest;
        //    mon_tr.io_diffCommits_info_50_pdest = io_diffCommits_info_50_pdest;
        //    mon_tr.io_diffCommits_info_50_rfWen = io_diffCommits_info_50_rfWen;
        //    mon_tr.io_diffCommits_info_50_fpWen = io_diffCommits_info_50_fpWen;
        //    mon_tr.io_diffCommits_info_50_vecWen = io_diffCommits_info_50_vecWen;
        //    mon_tr.io_diffCommits_info_50_v0Wen = io_diffCommits_info_50_v0Wen;
        //    mon_tr.io_diffCommits_info_50_vlWen = io_diffCommits_info_50_vlWen;
        //    mon_tr.io_diffCommits_info_51_ldest = io_diffCommits_info_51_ldest;
        //    mon_tr.io_diffCommits_info_51_pdest = io_diffCommits_info_51_pdest;
        //    mon_tr.io_diffCommits_info_51_rfWen = io_diffCommits_info_51_rfWen;
        //    mon_tr.io_diffCommits_info_51_fpWen = io_diffCommits_info_51_fpWen;
        //    mon_tr.io_diffCommits_info_51_vecWen = io_diffCommits_info_51_vecWen;
        //    mon_tr.io_diffCommits_info_51_v0Wen = io_diffCommits_info_51_v0Wen;
        //    mon_tr.io_diffCommits_info_51_vlWen = io_diffCommits_info_51_vlWen;
        //    mon_tr.io_diffCommits_info_52_ldest = io_diffCommits_info_52_ldest;
        //    mon_tr.io_diffCommits_info_52_pdest = io_diffCommits_info_52_pdest;
        //    mon_tr.io_diffCommits_info_52_rfWen = io_diffCommits_info_52_rfWen;
        //    mon_tr.io_diffCommits_info_52_fpWen = io_diffCommits_info_52_fpWen;
        //    mon_tr.io_diffCommits_info_52_vecWen = io_diffCommits_info_52_vecWen;
        //    mon_tr.io_diffCommits_info_52_v0Wen = io_diffCommits_info_52_v0Wen;
        //    mon_tr.io_diffCommits_info_52_vlWen = io_diffCommits_info_52_vlWen;
        //    mon_tr.io_diffCommits_info_53_ldest = io_diffCommits_info_53_ldest;
        //    mon_tr.io_diffCommits_info_53_pdest = io_diffCommits_info_53_pdest;
        //    mon_tr.io_diffCommits_info_53_rfWen = io_diffCommits_info_53_rfWen;
        //    mon_tr.io_diffCommits_info_53_fpWen = io_diffCommits_info_53_fpWen;
        //    mon_tr.io_diffCommits_info_53_vecWen = io_diffCommits_info_53_vecWen;
        //    mon_tr.io_diffCommits_info_53_v0Wen = io_diffCommits_info_53_v0Wen;
        //    mon_tr.io_diffCommits_info_53_vlWen = io_diffCommits_info_53_vlWen;
        //    mon_tr.io_diffCommits_info_54_ldest = io_diffCommits_info_54_ldest;
        //    mon_tr.io_diffCommits_info_54_pdest = io_diffCommits_info_54_pdest;
        //    mon_tr.io_diffCommits_info_54_rfWen = io_diffCommits_info_54_rfWen;
        //    mon_tr.io_diffCommits_info_54_fpWen = io_diffCommits_info_54_fpWen;
        //    mon_tr.io_diffCommits_info_54_vecWen = io_diffCommits_info_54_vecWen;
        //    mon_tr.io_diffCommits_info_54_v0Wen = io_diffCommits_info_54_v0Wen;
        //    mon_tr.io_diffCommits_info_54_vlWen = io_diffCommits_info_54_vlWen;
        //    mon_tr.io_diffCommits_info_55_ldest = io_diffCommits_info_55_ldest;
        //    mon_tr.io_diffCommits_info_55_pdest = io_diffCommits_info_55_pdest;
        //    mon_tr.io_diffCommits_info_55_rfWen = io_diffCommits_info_55_rfWen;
        //    mon_tr.io_diffCommits_info_55_fpWen = io_diffCommits_info_55_fpWen;
        //    mon_tr.io_diffCommits_info_55_vecWen = io_diffCommits_info_55_vecWen;
        //    mon_tr.io_diffCommits_info_55_v0Wen = io_diffCommits_info_55_v0Wen;
        //    mon_tr.io_diffCommits_info_55_vlWen = io_diffCommits_info_55_vlWen;
        //    mon_tr.io_diffCommits_info_56_ldest = io_diffCommits_info_56_ldest;
        //    mon_tr.io_diffCommits_info_56_pdest = io_diffCommits_info_56_pdest;
        //    mon_tr.io_diffCommits_info_56_rfWen = io_diffCommits_info_56_rfWen;
        //    mon_tr.io_diffCommits_info_56_fpWen = io_diffCommits_info_56_fpWen;
        //    mon_tr.io_diffCommits_info_56_vecWen = io_diffCommits_info_56_vecWen;
        //    mon_tr.io_diffCommits_info_56_v0Wen = io_diffCommits_info_56_v0Wen;
        //    mon_tr.io_diffCommits_info_56_vlWen = io_diffCommits_info_56_vlWen;
        //    mon_tr.io_diffCommits_info_57_ldest = io_diffCommits_info_57_ldest;
        //    mon_tr.io_diffCommits_info_57_pdest = io_diffCommits_info_57_pdest;
        //    mon_tr.io_diffCommits_info_57_rfWen = io_diffCommits_info_57_rfWen;
        //    mon_tr.io_diffCommits_info_57_fpWen = io_diffCommits_info_57_fpWen;
        //    mon_tr.io_diffCommits_info_57_vecWen = io_diffCommits_info_57_vecWen;
        //    mon_tr.io_diffCommits_info_57_v0Wen = io_diffCommits_info_57_v0Wen;
        //    mon_tr.io_diffCommits_info_57_vlWen = io_diffCommits_info_57_vlWen;
        //    mon_tr.io_diffCommits_info_58_ldest = io_diffCommits_info_58_ldest;
        //    mon_tr.io_diffCommits_info_58_pdest = io_diffCommits_info_58_pdest;
        //    mon_tr.io_diffCommits_info_58_rfWen = io_diffCommits_info_58_rfWen;
        //    mon_tr.io_diffCommits_info_58_fpWen = io_diffCommits_info_58_fpWen;
        //    mon_tr.io_diffCommits_info_58_vecWen = io_diffCommits_info_58_vecWen;
        //    mon_tr.io_diffCommits_info_58_v0Wen = io_diffCommits_info_58_v0Wen;
        //    mon_tr.io_diffCommits_info_58_vlWen = io_diffCommits_info_58_vlWen;
        //    mon_tr.io_diffCommits_info_59_ldest = io_diffCommits_info_59_ldest;
        //    mon_tr.io_diffCommits_info_59_pdest = io_diffCommits_info_59_pdest;
        //    mon_tr.io_diffCommits_info_59_rfWen = io_diffCommits_info_59_rfWen;
        //    mon_tr.io_diffCommits_info_59_fpWen = io_diffCommits_info_59_fpWen;
        //    mon_tr.io_diffCommits_info_59_vecWen = io_diffCommits_info_59_vecWen;
        //    mon_tr.io_diffCommits_info_59_v0Wen = io_diffCommits_info_59_v0Wen;
        //    mon_tr.io_diffCommits_info_59_vlWen = io_diffCommits_info_59_vlWen;
        //    mon_tr.io_diffCommits_info_60_ldest = io_diffCommits_info_60_ldest;
        //    mon_tr.io_diffCommits_info_60_pdest = io_diffCommits_info_60_pdest;
        //    mon_tr.io_diffCommits_info_60_rfWen = io_diffCommits_info_60_rfWen;
        //    mon_tr.io_diffCommits_info_60_fpWen = io_diffCommits_info_60_fpWen;
        //    mon_tr.io_diffCommits_info_60_vecWen = io_diffCommits_info_60_vecWen;
        //    mon_tr.io_diffCommits_info_60_v0Wen = io_diffCommits_info_60_v0Wen;
        //    mon_tr.io_diffCommits_info_60_vlWen = io_diffCommits_info_60_vlWen;
        //    mon_tr.io_diffCommits_info_61_ldest = io_diffCommits_info_61_ldest;
        //    mon_tr.io_diffCommits_info_61_pdest = io_diffCommits_info_61_pdest;
        //    mon_tr.io_diffCommits_info_61_rfWen = io_diffCommits_info_61_rfWen;
        //    mon_tr.io_diffCommits_info_61_fpWen = io_diffCommits_info_61_fpWen;
        //    mon_tr.io_diffCommits_info_61_vecWen = io_diffCommits_info_61_vecWen;
        //    mon_tr.io_diffCommits_info_61_v0Wen = io_diffCommits_info_61_v0Wen;
        //    mon_tr.io_diffCommits_info_61_vlWen = io_diffCommits_info_61_vlWen;
        //    mon_tr.io_diffCommits_info_62_ldest = io_diffCommits_info_62_ldest;
        //    mon_tr.io_diffCommits_info_62_pdest = io_diffCommits_info_62_pdest;
        //    mon_tr.io_diffCommits_info_62_rfWen = io_diffCommits_info_62_rfWen;
        //    mon_tr.io_diffCommits_info_62_fpWen = io_diffCommits_info_62_fpWen;
        //    mon_tr.io_diffCommits_info_62_vecWen = io_diffCommits_info_62_vecWen;
        //    mon_tr.io_diffCommits_info_62_v0Wen = io_diffCommits_info_62_v0Wen;
        //    mon_tr.io_diffCommits_info_62_vlWen = io_diffCommits_info_62_vlWen;
        //    mon_tr.io_diffCommits_info_63_ldest = io_diffCommits_info_63_ldest;
        //    mon_tr.io_diffCommits_info_63_pdest = io_diffCommits_info_63_pdest;
        //    mon_tr.io_diffCommits_info_63_rfWen = io_diffCommits_info_63_rfWen;
        //    mon_tr.io_diffCommits_info_63_fpWen = io_diffCommits_info_63_fpWen;
        //    mon_tr.io_diffCommits_info_63_vecWen = io_diffCommits_info_63_vecWen;
        //    mon_tr.io_diffCommits_info_63_v0Wen = io_diffCommits_info_63_v0Wen;
        //    mon_tr.io_diffCommits_info_63_vlWen = io_diffCommits_info_63_vlWen;
        //    mon_tr.io_diffCommits_info_64_ldest = io_diffCommits_info_64_ldest;
        //    mon_tr.io_diffCommits_info_64_pdest = io_diffCommits_info_64_pdest;
        //    mon_tr.io_diffCommits_info_64_rfWen = io_diffCommits_info_64_rfWen;
        //    mon_tr.io_diffCommits_info_64_fpWen = io_diffCommits_info_64_fpWen;
        //    mon_tr.io_diffCommits_info_64_vecWen = io_diffCommits_info_64_vecWen;
        //    mon_tr.io_diffCommits_info_64_v0Wen = io_diffCommits_info_64_v0Wen;
        //    mon_tr.io_diffCommits_info_64_vlWen = io_diffCommits_info_64_vlWen;
        //    mon_tr.io_diffCommits_info_65_ldest = io_diffCommits_info_65_ldest;
        //    mon_tr.io_diffCommits_info_65_pdest = io_diffCommits_info_65_pdest;
        //    mon_tr.io_diffCommits_info_65_rfWen = io_diffCommits_info_65_rfWen;
        //    mon_tr.io_diffCommits_info_65_fpWen = io_diffCommits_info_65_fpWen;
        //    mon_tr.io_diffCommits_info_65_vecWen = io_diffCommits_info_65_vecWen;
        //    mon_tr.io_diffCommits_info_65_v0Wen = io_diffCommits_info_65_v0Wen;
        //    mon_tr.io_diffCommits_info_65_vlWen = io_diffCommits_info_65_vlWen;
        //    mon_tr.io_diffCommits_info_66_ldest = io_diffCommits_info_66_ldest;
        //    mon_tr.io_diffCommits_info_66_pdest = io_diffCommits_info_66_pdest;
        //    mon_tr.io_diffCommits_info_66_rfWen = io_diffCommits_info_66_rfWen;
        //    mon_tr.io_diffCommits_info_66_fpWen = io_diffCommits_info_66_fpWen;
        //    mon_tr.io_diffCommits_info_66_vecWen = io_diffCommits_info_66_vecWen;
        //    mon_tr.io_diffCommits_info_66_v0Wen = io_diffCommits_info_66_v0Wen;
        //    mon_tr.io_diffCommits_info_66_vlWen = io_diffCommits_info_66_vlWen;
        //    mon_tr.io_diffCommits_info_67_ldest = io_diffCommits_info_67_ldest;
        //    mon_tr.io_diffCommits_info_67_pdest = io_diffCommits_info_67_pdest;
        //    mon_tr.io_diffCommits_info_67_rfWen = io_diffCommits_info_67_rfWen;
        //    mon_tr.io_diffCommits_info_67_fpWen = io_diffCommits_info_67_fpWen;
        //    mon_tr.io_diffCommits_info_67_vecWen = io_diffCommits_info_67_vecWen;
        //    mon_tr.io_diffCommits_info_67_v0Wen = io_diffCommits_info_67_v0Wen;
        //    mon_tr.io_diffCommits_info_67_vlWen = io_diffCommits_info_67_vlWen;
        //    mon_tr.io_diffCommits_info_68_ldest = io_diffCommits_info_68_ldest;
        //    mon_tr.io_diffCommits_info_68_pdest = io_diffCommits_info_68_pdest;
        //    mon_tr.io_diffCommits_info_68_rfWen = io_diffCommits_info_68_rfWen;
        //    mon_tr.io_diffCommits_info_68_fpWen = io_diffCommits_info_68_fpWen;
        //    mon_tr.io_diffCommits_info_68_vecWen = io_diffCommits_info_68_vecWen;
        //    mon_tr.io_diffCommits_info_68_v0Wen = io_diffCommits_info_68_v0Wen;
        //    mon_tr.io_diffCommits_info_68_vlWen = io_diffCommits_info_68_vlWen;
        //    mon_tr.io_diffCommits_info_69_ldest = io_diffCommits_info_69_ldest;
        //    mon_tr.io_diffCommits_info_69_pdest = io_diffCommits_info_69_pdest;
        //    mon_tr.io_diffCommits_info_69_rfWen = io_diffCommits_info_69_rfWen;
        //    mon_tr.io_diffCommits_info_69_fpWen = io_diffCommits_info_69_fpWen;
        //    mon_tr.io_diffCommits_info_69_vecWen = io_diffCommits_info_69_vecWen;
        //    mon_tr.io_diffCommits_info_69_v0Wen = io_diffCommits_info_69_v0Wen;
        //    mon_tr.io_diffCommits_info_69_vlWen = io_diffCommits_info_69_vlWen;
        //    mon_tr.io_diffCommits_info_70_ldest = io_diffCommits_info_70_ldest;
        //    mon_tr.io_diffCommits_info_70_pdest = io_diffCommits_info_70_pdest;
        //    mon_tr.io_diffCommits_info_70_rfWen = io_diffCommits_info_70_rfWen;
        //    mon_tr.io_diffCommits_info_70_fpWen = io_diffCommits_info_70_fpWen;
        //    mon_tr.io_diffCommits_info_70_vecWen = io_diffCommits_info_70_vecWen;
        //    mon_tr.io_diffCommits_info_70_v0Wen = io_diffCommits_info_70_v0Wen;
        //    mon_tr.io_diffCommits_info_70_vlWen = io_diffCommits_info_70_vlWen;
        //    mon_tr.io_diffCommits_info_71_ldest = io_diffCommits_info_71_ldest;
        //    mon_tr.io_diffCommits_info_71_pdest = io_diffCommits_info_71_pdest;
        //    mon_tr.io_diffCommits_info_71_rfWen = io_diffCommits_info_71_rfWen;
        //    mon_tr.io_diffCommits_info_71_fpWen = io_diffCommits_info_71_fpWen;
        //    mon_tr.io_diffCommits_info_71_vecWen = io_diffCommits_info_71_vecWen;
        //    mon_tr.io_diffCommits_info_71_v0Wen = io_diffCommits_info_71_v0Wen;
        //    mon_tr.io_diffCommits_info_71_vlWen = io_diffCommits_info_71_vlWen;
        //    mon_tr.io_diffCommits_info_72_ldest = io_diffCommits_info_72_ldest;
        //    mon_tr.io_diffCommits_info_72_pdest = io_diffCommits_info_72_pdest;
        //    mon_tr.io_diffCommits_info_72_rfWen = io_diffCommits_info_72_rfWen;
        //    mon_tr.io_diffCommits_info_72_fpWen = io_diffCommits_info_72_fpWen;
        //    mon_tr.io_diffCommits_info_72_vecWen = io_diffCommits_info_72_vecWen;
        //    mon_tr.io_diffCommits_info_72_v0Wen = io_diffCommits_info_72_v0Wen;
        //    mon_tr.io_diffCommits_info_72_vlWen = io_diffCommits_info_72_vlWen;
        //    mon_tr.io_diffCommits_info_73_ldest = io_diffCommits_info_73_ldest;
        //    mon_tr.io_diffCommits_info_73_pdest = io_diffCommits_info_73_pdest;
        //    mon_tr.io_diffCommits_info_73_rfWen = io_diffCommits_info_73_rfWen;
        //    mon_tr.io_diffCommits_info_73_fpWen = io_diffCommits_info_73_fpWen;
        //    mon_tr.io_diffCommits_info_73_vecWen = io_diffCommits_info_73_vecWen;
        //    mon_tr.io_diffCommits_info_73_v0Wen = io_diffCommits_info_73_v0Wen;
        //    mon_tr.io_diffCommits_info_73_vlWen = io_diffCommits_info_73_vlWen;
        //    mon_tr.io_diffCommits_info_74_ldest = io_diffCommits_info_74_ldest;
        //    mon_tr.io_diffCommits_info_74_pdest = io_diffCommits_info_74_pdest;
        //    mon_tr.io_diffCommits_info_74_rfWen = io_diffCommits_info_74_rfWen;
        //    mon_tr.io_diffCommits_info_74_fpWen = io_diffCommits_info_74_fpWen;
        //    mon_tr.io_diffCommits_info_74_vecWen = io_diffCommits_info_74_vecWen;
        //    mon_tr.io_diffCommits_info_74_v0Wen = io_diffCommits_info_74_v0Wen;
        //    mon_tr.io_diffCommits_info_74_vlWen = io_diffCommits_info_74_vlWen;
        //    mon_tr.io_diffCommits_info_75_ldest = io_diffCommits_info_75_ldest;
        //    mon_tr.io_diffCommits_info_75_pdest = io_diffCommits_info_75_pdest;
        //    mon_tr.io_diffCommits_info_75_rfWen = io_diffCommits_info_75_rfWen;
        //    mon_tr.io_diffCommits_info_75_fpWen = io_diffCommits_info_75_fpWen;
        //    mon_tr.io_diffCommits_info_75_vecWen = io_diffCommits_info_75_vecWen;
        //    mon_tr.io_diffCommits_info_75_v0Wen = io_diffCommits_info_75_v0Wen;
        //    mon_tr.io_diffCommits_info_75_vlWen = io_diffCommits_info_75_vlWen;
        //    mon_tr.io_diffCommits_info_76_ldest = io_diffCommits_info_76_ldest;
        //    mon_tr.io_diffCommits_info_76_pdest = io_diffCommits_info_76_pdest;
        //    mon_tr.io_diffCommits_info_76_rfWen = io_diffCommits_info_76_rfWen;
        //    mon_tr.io_diffCommits_info_76_fpWen = io_diffCommits_info_76_fpWen;
        //    mon_tr.io_diffCommits_info_76_vecWen = io_diffCommits_info_76_vecWen;
        //    mon_tr.io_diffCommits_info_76_v0Wen = io_diffCommits_info_76_v0Wen;
        //    mon_tr.io_diffCommits_info_76_vlWen = io_diffCommits_info_76_vlWen;
        //    mon_tr.io_diffCommits_info_77_ldest = io_diffCommits_info_77_ldest;
        //    mon_tr.io_diffCommits_info_77_pdest = io_diffCommits_info_77_pdest;
        //    mon_tr.io_diffCommits_info_77_rfWen = io_diffCommits_info_77_rfWen;
        //    mon_tr.io_diffCommits_info_77_fpWen = io_diffCommits_info_77_fpWen;
        //    mon_tr.io_diffCommits_info_77_vecWen = io_diffCommits_info_77_vecWen;
        //    mon_tr.io_diffCommits_info_77_v0Wen = io_diffCommits_info_77_v0Wen;
        //    mon_tr.io_diffCommits_info_77_vlWen = io_diffCommits_info_77_vlWen;
        //    mon_tr.io_diffCommits_info_78_ldest = io_diffCommits_info_78_ldest;
        //    mon_tr.io_diffCommits_info_78_pdest = io_diffCommits_info_78_pdest;
        //    mon_tr.io_diffCommits_info_78_rfWen = io_diffCommits_info_78_rfWen;
        //    mon_tr.io_diffCommits_info_78_fpWen = io_diffCommits_info_78_fpWen;
        //    mon_tr.io_diffCommits_info_78_vecWen = io_diffCommits_info_78_vecWen;
        //    mon_tr.io_diffCommits_info_78_v0Wen = io_diffCommits_info_78_v0Wen;
        //    mon_tr.io_diffCommits_info_78_vlWen = io_diffCommits_info_78_vlWen;
        //    mon_tr.io_diffCommits_info_79_ldest = io_diffCommits_info_79_ldest;
        //    mon_tr.io_diffCommits_info_79_pdest = io_diffCommits_info_79_pdest;
        //    mon_tr.io_diffCommits_info_79_rfWen = io_diffCommits_info_79_rfWen;
        //    mon_tr.io_diffCommits_info_79_fpWen = io_diffCommits_info_79_fpWen;
        //    mon_tr.io_diffCommits_info_79_vecWen = io_diffCommits_info_79_vecWen;
        //    mon_tr.io_diffCommits_info_79_v0Wen = io_diffCommits_info_79_v0Wen;
        //    mon_tr.io_diffCommits_info_79_vlWen = io_diffCommits_info_79_vlWen;
        //    mon_tr.io_diffCommits_info_80_ldest = io_diffCommits_info_80_ldest;
        //    mon_tr.io_diffCommits_info_80_pdest = io_diffCommits_info_80_pdest;
        //    mon_tr.io_diffCommits_info_80_rfWen = io_diffCommits_info_80_rfWen;
        //    mon_tr.io_diffCommits_info_80_fpWen = io_diffCommits_info_80_fpWen;
        //    mon_tr.io_diffCommits_info_80_vecWen = io_diffCommits_info_80_vecWen;
        //    mon_tr.io_diffCommits_info_80_v0Wen = io_diffCommits_info_80_v0Wen;
        //    mon_tr.io_diffCommits_info_80_vlWen = io_diffCommits_info_80_vlWen;
        //    mon_tr.io_diffCommits_info_81_ldest = io_diffCommits_info_81_ldest;
        //    mon_tr.io_diffCommits_info_81_pdest = io_diffCommits_info_81_pdest;
        //    mon_tr.io_diffCommits_info_81_rfWen = io_diffCommits_info_81_rfWen;
        //    mon_tr.io_diffCommits_info_81_fpWen = io_diffCommits_info_81_fpWen;
        //    mon_tr.io_diffCommits_info_81_vecWen = io_diffCommits_info_81_vecWen;
        //    mon_tr.io_diffCommits_info_81_v0Wen = io_diffCommits_info_81_v0Wen;
        //    mon_tr.io_diffCommits_info_81_vlWen = io_diffCommits_info_81_vlWen;
        //    mon_tr.io_diffCommits_info_82_ldest = io_diffCommits_info_82_ldest;
        //    mon_tr.io_diffCommits_info_82_pdest = io_diffCommits_info_82_pdest;
        //    mon_tr.io_diffCommits_info_82_rfWen = io_diffCommits_info_82_rfWen;
        //    mon_tr.io_diffCommits_info_82_fpWen = io_diffCommits_info_82_fpWen;
        //    mon_tr.io_diffCommits_info_82_vecWen = io_diffCommits_info_82_vecWen;
        //    mon_tr.io_diffCommits_info_82_v0Wen = io_diffCommits_info_82_v0Wen;
        //    mon_tr.io_diffCommits_info_82_vlWen = io_diffCommits_info_82_vlWen;
        //    mon_tr.io_diffCommits_info_83_ldest = io_diffCommits_info_83_ldest;
        //    mon_tr.io_diffCommits_info_83_pdest = io_diffCommits_info_83_pdest;
        //    mon_tr.io_diffCommits_info_83_rfWen = io_diffCommits_info_83_rfWen;
        //    mon_tr.io_diffCommits_info_83_fpWen = io_diffCommits_info_83_fpWen;
        //    mon_tr.io_diffCommits_info_83_vecWen = io_diffCommits_info_83_vecWen;
        //    mon_tr.io_diffCommits_info_83_v0Wen = io_diffCommits_info_83_v0Wen;
        //    mon_tr.io_diffCommits_info_83_vlWen = io_diffCommits_info_83_vlWen;
        //    mon_tr.io_diffCommits_info_84_ldest = io_diffCommits_info_84_ldest;
        //    mon_tr.io_diffCommits_info_84_pdest = io_diffCommits_info_84_pdest;
        //    mon_tr.io_diffCommits_info_84_rfWen = io_diffCommits_info_84_rfWen;
        //    mon_tr.io_diffCommits_info_84_fpWen = io_diffCommits_info_84_fpWen;
        //    mon_tr.io_diffCommits_info_84_vecWen = io_diffCommits_info_84_vecWen;
        //    mon_tr.io_diffCommits_info_84_v0Wen = io_diffCommits_info_84_v0Wen;
        //    mon_tr.io_diffCommits_info_84_vlWen = io_diffCommits_info_84_vlWen;
        //    mon_tr.io_diffCommits_info_85_ldest = io_diffCommits_info_85_ldest;
        //    mon_tr.io_diffCommits_info_85_pdest = io_diffCommits_info_85_pdest;
        //    mon_tr.io_diffCommits_info_85_rfWen = io_diffCommits_info_85_rfWen;
        //    mon_tr.io_diffCommits_info_85_fpWen = io_diffCommits_info_85_fpWen;
        //    mon_tr.io_diffCommits_info_85_vecWen = io_diffCommits_info_85_vecWen;
        //    mon_tr.io_diffCommits_info_85_v0Wen = io_diffCommits_info_85_v0Wen;
        //    mon_tr.io_diffCommits_info_85_vlWen = io_diffCommits_info_85_vlWen;
        //    mon_tr.io_diffCommits_info_86_ldest = io_diffCommits_info_86_ldest;
        //    mon_tr.io_diffCommits_info_86_pdest = io_diffCommits_info_86_pdest;
        //    mon_tr.io_diffCommits_info_86_rfWen = io_diffCommits_info_86_rfWen;
        //    mon_tr.io_diffCommits_info_86_fpWen = io_diffCommits_info_86_fpWen;
        //    mon_tr.io_diffCommits_info_86_vecWen = io_diffCommits_info_86_vecWen;
        //    mon_tr.io_diffCommits_info_86_v0Wen = io_diffCommits_info_86_v0Wen;
        //    mon_tr.io_diffCommits_info_86_vlWen = io_diffCommits_info_86_vlWen;
        //    mon_tr.io_diffCommits_info_87_ldest = io_diffCommits_info_87_ldest;
        //    mon_tr.io_diffCommits_info_87_pdest = io_diffCommits_info_87_pdest;
        //    mon_tr.io_diffCommits_info_87_rfWen = io_diffCommits_info_87_rfWen;
        //    mon_tr.io_diffCommits_info_87_fpWen = io_diffCommits_info_87_fpWen;
        //    mon_tr.io_diffCommits_info_87_vecWen = io_diffCommits_info_87_vecWen;
        //    mon_tr.io_diffCommits_info_87_v0Wen = io_diffCommits_info_87_v0Wen;
        //    mon_tr.io_diffCommits_info_87_vlWen = io_diffCommits_info_87_vlWen;
        //    mon_tr.io_diffCommits_info_88_ldest = io_diffCommits_info_88_ldest;
        //    mon_tr.io_diffCommits_info_88_pdest = io_diffCommits_info_88_pdest;
        //    mon_tr.io_diffCommits_info_88_rfWen = io_diffCommits_info_88_rfWen;
        //    mon_tr.io_diffCommits_info_88_fpWen = io_diffCommits_info_88_fpWen;
        //    mon_tr.io_diffCommits_info_88_vecWen = io_diffCommits_info_88_vecWen;
        //    mon_tr.io_diffCommits_info_88_v0Wen = io_diffCommits_info_88_v0Wen;
        //    mon_tr.io_diffCommits_info_88_vlWen = io_diffCommits_info_88_vlWen;
        //    mon_tr.io_diffCommits_info_89_ldest = io_diffCommits_info_89_ldest;
        //    mon_tr.io_diffCommits_info_89_pdest = io_diffCommits_info_89_pdest;
        //    mon_tr.io_diffCommits_info_89_rfWen = io_diffCommits_info_89_rfWen;
        //    mon_tr.io_diffCommits_info_89_fpWen = io_diffCommits_info_89_fpWen;
        //    mon_tr.io_diffCommits_info_89_vecWen = io_diffCommits_info_89_vecWen;
        //    mon_tr.io_diffCommits_info_89_v0Wen = io_diffCommits_info_89_v0Wen;
        //    mon_tr.io_diffCommits_info_89_vlWen = io_diffCommits_info_89_vlWen;
        //    mon_tr.io_diffCommits_info_90_ldest = io_diffCommits_info_90_ldest;
        //    mon_tr.io_diffCommits_info_90_pdest = io_diffCommits_info_90_pdest;
        //    mon_tr.io_diffCommits_info_90_rfWen = io_diffCommits_info_90_rfWen;
        //    mon_tr.io_diffCommits_info_90_fpWen = io_diffCommits_info_90_fpWen;
        //    mon_tr.io_diffCommits_info_90_vecWen = io_diffCommits_info_90_vecWen;
        //    mon_tr.io_diffCommits_info_90_v0Wen = io_diffCommits_info_90_v0Wen;
        //    mon_tr.io_diffCommits_info_90_vlWen = io_diffCommits_info_90_vlWen;
        //    mon_tr.io_diffCommits_info_91_ldest = io_diffCommits_info_91_ldest;
        //    mon_tr.io_diffCommits_info_91_pdest = io_diffCommits_info_91_pdest;
        //    mon_tr.io_diffCommits_info_91_rfWen = io_diffCommits_info_91_rfWen;
        //    mon_tr.io_diffCommits_info_91_fpWen = io_diffCommits_info_91_fpWen;
        //    mon_tr.io_diffCommits_info_91_vecWen = io_diffCommits_info_91_vecWen;
        //    mon_tr.io_diffCommits_info_91_v0Wen = io_diffCommits_info_91_v0Wen;
        //    mon_tr.io_diffCommits_info_91_vlWen = io_diffCommits_info_91_vlWen;
        //    mon_tr.io_diffCommits_info_92_ldest = io_diffCommits_info_92_ldest;
        //    mon_tr.io_diffCommits_info_92_pdest = io_diffCommits_info_92_pdest;
        //    mon_tr.io_diffCommits_info_92_rfWen = io_diffCommits_info_92_rfWen;
        //    mon_tr.io_diffCommits_info_92_fpWen = io_diffCommits_info_92_fpWen;
        //    mon_tr.io_diffCommits_info_92_vecWen = io_diffCommits_info_92_vecWen;
        //    mon_tr.io_diffCommits_info_92_v0Wen = io_diffCommits_info_92_v0Wen;
        //    mon_tr.io_diffCommits_info_92_vlWen = io_diffCommits_info_92_vlWen;
        //    mon_tr.io_diffCommits_info_93_ldest = io_diffCommits_info_93_ldest;
        //    mon_tr.io_diffCommits_info_93_pdest = io_diffCommits_info_93_pdest;
        //    mon_tr.io_diffCommits_info_93_rfWen = io_diffCommits_info_93_rfWen;
        //    mon_tr.io_diffCommits_info_93_fpWen = io_diffCommits_info_93_fpWen;
        //    mon_tr.io_diffCommits_info_93_vecWen = io_diffCommits_info_93_vecWen;
        //    mon_tr.io_diffCommits_info_93_v0Wen = io_diffCommits_info_93_v0Wen;
        //    mon_tr.io_diffCommits_info_93_vlWen = io_diffCommits_info_93_vlWen;
        //    mon_tr.io_diffCommits_info_94_ldest = io_diffCommits_info_94_ldest;
        //    mon_tr.io_diffCommits_info_94_pdest = io_diffCommits_info_94_pdest;
        //    mon_tr.io_diffCommits_info_94_rfWen = io_diffCommits_info_94_rfWen;
        //    mon_tr.io_diffCommits_info_94_fpWen = io_diffCommits_info_94_fpWen;
        //    mon_tr.io_diffCommits_info_94_vecWen = io_diffCommits_info_94_vecWen;
        //    mon_tr.io_diffCommits_info_94_v0Wen = io_diffCommits_info_94_v0Wen;
        //    mon_tr.io_diffCommits_info_94_vlWen = io_diffCommits_info_94_vlWen;
        //    mon_tr.io_diffCommits_info_95_ldest = io_diffCommits_info_95_ldest;
        //    mon_tr.io_diffCommits_info_95_pdest = io_diffCommits_info_95_pdest;
        //    mon_tr.io_diffCommits_info_95_rfWen = io_diffCommits_info_95_rfWen;
        //    mon_tr.io_diffCommits_info_95_fpWen = io_diffCommits_info_95_fpWen;
        //    mon_tr.io_diffCommits_info_95_vecWen = io_diffCommits_info_95_vecWen;
        //    mon_tr.io_diffCommits_info_95_v0Wen = io_diffCommits_info_95_v0Wen;
        //    mon_tr.io_diffCommits_info_95_vlWen = io_diffCommits_info_95_vlWen;
        //    mon_tr.io_diffCommits_info_96_ldest = io_diffCommits_info_96_ldest;
        //    mon_tr.io_diffCommits_info_96_pdest = io_diffCommits_info_96_pdest;
        //    mon_tr.io_diffCommits_info_96_rfWen = io_diffCommits_info_96_rfWen;
        //    mon_tr.io_diffCommits_info_96_fpWen = io_diffCommits_info_96_fpWen;
        //    mon_tr.io_diffCommits_info_96_vecWen = io_diffCommits_info_96_vecWen;
        //    mon_tr.io_diffCommits_info_96_v0Wen = io_diffCommits_info_96_v0Wen;
        //    mon_tr.io_diffCommits_info_96_vlWen = io_diffCommits_info_96_vlWen;
        //    mon_tr.io_diffCommits_info_97_ldest = io_diffCommits_info_97_ldest;
        //    mon_tr.io_diffCommits_info_97_pdest = io_diffCommits_info_97_pdest;
        //    mon_tr.io_diffCommits_info_97_rfWen = io_diffCommits_info_97_rfWen;
        //    mon_tr.io_diffCommits_info_97_fpWen = io_diffCommits_info_97_fpWen;
        //    mon_tr.io_diffCommits_info_97_vecWen = io_diffCommits_info_97_vecWen;
        //    mon_tr.io_diffCommits_info_97_v0Wen = io_diffCommits_info_97_v0Wen;
        //    mon_tr.io_diffCommits_info_97_vlWen = io_diffCommits_info_97_vlWen;
        //    mon_tr.io_diffCommits_info_98_ldest = io_diffCommits_info_98_ldest;
        //    mon_tr.io_diffCommits_info_98_pdest = io_diffCommits_info_98_pdest;
        //    mon_tr.io_diffCommits_info_98_rfWen = io_diffCommits_info_98_rfWen;
        //    mon_tr.io_diffCommits_info_98_fpWen = io_diffCommits_info_98_fpWen;
        //    mon_tr.io_diffCommits_info_98_vecWen = io_diffCommits_info_98_vecWen;
        //    mon_tr.io_diffCommits_info_98_v0Wen = io_diffCommits_info_98_v0Wen;
        //    mon_tr.io_diffCommits_info_98_vlWen = io_diffCommits_info_98_vlWen;
        //    mon_tr.io_diffCommits_info_99_ldest = io_diffCommits_info_99_ldest;
        //    mon_tr.io_diffCommits_info_99_pdest = io_diffCommits_info_99_pdest;
        //    mon_tr.io_diffCommits_info_99_rfWen = io_diffCommits_info_99_rfWen;
        //    mon_tr.io_diffCommits_info_99_fpWen = io_diffCommits_info_99_fpWen;
        //    mon_tr.io_diffCommits_info_99_vecWen = io_diffCommits_info_99_vecWen;
        //    mon_tr.io_diffCommits_info_99_v0Wen = io_diffCommits_info_99_v0Wen;
        //    mon_tr.io_diffCommits_info_99_vlWen = io_diffCommits_info_99_vlWen;
        //    mon_tr.io_diffCommits_info_100_ldest = io_diffCommits_info_100_ldest;
        //    mon_tr.io_diffCommits_info_100_pdest = io_diffCommits_info_100_pdest;
        //    mon_tr.io_diffCommits_info_100_rfWen = io_diffCommits_info_100_rfWen;
        //    mon_tr.io_diffCommits_info_100_fpWen = io_diffCommits_info_100_fpWen;
        //    mon_tr.io_diffCommits_info_100_vecWen = io_diffCommits_info_100_vecWen;
        //    mon_tr.io_diffCommits_info_100_v0Wen = io_diffCommits_info_100_v0Wen;
        //    mon_tr.io_diffCommits_info_100_vlWen = io_diffCommits_info_100_vlWen;
        //    mon_tr.io_diffCommits_info_101_ldest = io_diffCommits_info_101_ldest;
        //    mon_tr.io_diffCommits_info_101_pdest = io_diffCommits_info_101_pdest;
        //    mon_tr.io_diffCommits_info_101_rfWen = io_diffCommits_info_101_rfWen;
        //    mon_tr.io_diffCommits_info_101_fpWen = io_diffCommits_info_101_fpWen;
        //    mon_tr.io_diffCommits_info_101_vecWen = io_diffCommits_info_101_vecWen;
        //    mon_tr.io_diffCommits_info_101_v0Wen = io_diffCommits_info_101_v0Wen;
        //    mon_tr.io_diffCommits_info_101_vlWen = io_diffCommits_info_101_vlWen;
        //    mon_tr.io_diffCommits_info_102_ldest = io_diffCommits_info_102_ldest;
        //    mon_tr.io_diffCommits_info_102_pdest = io_diffCommits_info_102_pdest;
        //    mon_tr.io_diffCommits_info_102_rfWen = io_diffCommits_info_102_rfWen;
        //    mon_tr.io_diffCommits_info_102_fpWen = io_diffCommits_info_102_fpWen;
        //    mon_tr.io_diffCommits_info_102_vecWen = io_diffCommits_info_102_vecWen;
        //    mon_tr.io_diffCommits_info_102_v0Wen = io_diffCommits_info_102_v0Wen;
        //    mon_tr.io_diffCommits_info_102_vlWen = io_diffCommits_info_102_vlWen;
        //    mon_tr.io_diffCommits_info_103_ldest = io_diffCommits_info_103_ldest;
        //    mon_tr.io_diffCommits_info_103_pdest = io_diffCommits_info_103_pdest;
        //    mon_tr.io_diffCommits_info_103_rfWen = io_diffCommits_info_103_rfWen;
        //    mon_tr.io_diffCommits_info_103_fpWen = io_diffCommits_info_103_fpWen;
        //    mon_tr.io_diffCommits_info_103_vecWen = io_diffCommits_info_103_vecWen;
        //    mon_tr.io_diffCommits_info_103_v0Wen = io_diffCommits_info_103_v0Wen;
        //    mon_tr.io_diffCommits_info_103_vlWen = io_diffCommits_info_103_vlWen;
        //    mon_tr.io_diffCommits_info_104_ldest = io_diffCommits_info_104_ldest;
        //    mon_tr.io_diffCommits_info_104_pdest = io_diffCommits_info_104_pdest;
        //    mon_tr.io_diffCommits_info_104_rfWen = io_diffCommits_info_104_rfWen;
        //    mon_tr.io_diffCommits_info_104_fpWen = io_diffCommits_info_104_fpWen;
        //    mon_tr.io_diffCommits_info_104_vecWen = io_diffCommits_info_104_vecWen;
        //    mon_tr.io_diffCommits_info_104_v0Wen = io_diffCommits_info_104_v0Wen;
        //    mon_tr.io_diffCommits_info_104_vlWen = io_diffCommits_info_104_vlWen;
        //    mon_tr.io_diffCommits_info_105_ldest = io_diffCommits_info_105_ldest;
        //    mon_tr.io_diffCommits_info_105_pdest = io_diffCommits_info_105_pdest;
        //    mon_tr.io_diffCommits_info_105_rfWen = io_diffCommits_info_105_rfWen;
        //    mon_tr.io_diffCommits_info_105_fpWen = io_diffCommits_info_105_fpWen;
        //    mon_tr.io_diffCommits_info_105_vecWen = io_diffCommits_info_105_vecWen;
        //    mon_tr.io_diffCommits_info_105_v0Wen = io_diffCommits_info_105_v0Wen;
        //    mon_tr.io_diffCommits_info_105_vlWen = io_diffCommits_info_105_vlWen;
        //    mon_tr.io_diffCommits_info_106_ldest = io_diffCommits_info_106_ldest;
        //    mon_tr.io_diffCommits_info_106_pdest = io_diffCommits_info_106_pdest;
        //    mon_tr.io_diffCommits_info_106_rfWen = io_diffCommits_info_106_rfWen;
        //    mon_tr.io_diffCommits_info_106_fpWen = io_diffCommits_info_106_fpWen;
        //    mon_tr.io_diffCommits_info_106_vecWen = io_diffCommits_info_106_vecWen;
        //    mon_tr.io_diffCommits_info_106_v0Wen = io_diffCommits_info_106_v0Wen;
        //    mon_tr.io_diffCommits_info_106_vlWen = io_diffCommits_info_106_vlWen;
        //    mon_tr.io_diffCommits_info_107_ldest = io_diffCommits_info_107_ldest;
        //    mon_tr.io_diffCommits_info_107_pdest = io_diffCommits_info_107_pdest;
        //    mon_tr.io_diffCommits_info_107_rfWen = io_diffCommits_info_107_rfWen;
        //    mon_tr.io_diffCommits_info_107_fpWen = io_diffCommits_info_107_fpWen;
        //    mon_tr.io_diffCommits_info_107_vecWen = io_diffCommits_info_107_vecWen;
        //    mon_tr.io_diffCommits_info_107_v0Wen = io_diffCommits_info_107_v0Wen;
        //    mon_tr.io_diffCommits_info_107_vlWen = io_diffCommits_info_107_vlWen;
        //    mon_tr.io_diffCommits_info_108_ldest = io_diffCommits_info_108_ldest;
        //    mon_tr.io_diffCommits_info_108_pdest = io_diffCommits_info_108_pdest;
        //    mon_tr.io_diffCommits_info_108_rfWen = io_diffCommits_info_108_rfWen;
        //    mon_tr.io_diffCommits_info_108_fpWen = io_diffCommits_info_108_fpWen;
        //    mon_tr.io_diffCommits_info_108_vecWen = io_diffCommits_info_108_vecWen;
        //    mon_tr.io_diffCommits_info_108_v0Wen = io_diffCommits_info_108_v0Wen;
        //    mon_tr.io_diffCommits_info_108_vlWen = io_diffCommits_info_108_vlWen;
        //    mon_tr.io_diffCommits_info_109_ldest = io_diffCommits_info_109_ldest;
        //    mon_tr.io_diffCommits_info_109_pdest = io_diffCommits_info_109_pdest;
        //    mon_tr.io_diffCommits_info_109_rfWen = io_diffCommits_info_109_rfWen;
        //    mon_tr.io_diffCommits_info_109_fpWen = io_diffCommits_info_109_fpWen;
        //    mon_tr.io_diffCommits_info_109_vecWen = io_diffCommits_info_109_vecWen;
        //    mon_tr.io_diffCommits_info_109_v0Wen = io_diffCommits_info_109_v0Wen;
        //    mon_tr.io_diffCommits_info_109_vlWen = io_diffCommits_info_109_vlWen;
        //    mon_tr.io_diffCommits_info_110_ldest = io_diffCommits_info_110_ldest;
        //    mon_tr.io_diffCommits_info_110_pdest = io_diffCommits_info_110_pdest;
        //    mon_tr.io_diffCommits_info_110_rfWen = io_diffCommits_info_110_rfWen;
        //    mon_tr.io_diffCommits_info_110_fpWen = io_diffCommits_info_110_fpWen;
        //    mon_tr.io_diffCommits_info_110_vecWen = io_diffCommits_info_110_vecWen;
        //    mon_tr.io_diffCommits_info_110_v0Wen = io_diffCommits_info_110_v0Wen;
        //    mon_tr.io_diffCommits_info_110_vlWen = io_diffCommits_info_110_vlWen;
        //    mon_tr.io_diffCommits_info_111_ldest = io_diffCommits_info_111_ldest;
        //    mon_tr.io_diffCommits_info_111_pdest = io_diffCommits_info_111_pdest;
        //    mon_tr.io_diffCommits_info_111_rfWen = io_diffCommits_info_111_rfWen;
        //    mon_tr.io_diffCommits_info_111_fpWen = io_diffCommits_info_111_fpWen;
        //    mon_tr.io_diffCommits_info_111_vecWen = io_diffCommits_info_111_vecWen;
        //    mon_tr.io_diffCommits_info_111_v0Wen = io_diffCommits_info_111_v0Wen;
        //    mon_tr.io_diffCommits_info_111_vlWen = io_diffCommits_info_111_vlWen;
        //    mon_tr.io_diffCommits_info_112_ldest = io_diffCommits_info_112_ldest;
        //    mon_tr.io_diffCommits_info_112_pdest = io_diffCommits_info_112_pdest;
        //    mon_tr.io_diffCommits_info_112_rfWen = io_diffCommits_info_112_rfWen;
        //    mon_tr.io_diffCommits_info_112_fpWen = io_diffCommits_info_112_fpWen;
        //    mon_tr.io_diffCommits_info_112_vecWen = io_diffCommits_info_112_vecWen;
        //    mon_tr.io_diffCommits_info_112_v0Wen = io_diffCommits_info_112_v0Wen;
        //    mon_tr.io_diffCommits_info_112_vlWen = io_diffCommits_info_112_vlWen;
        //    mon_tr.io_diffCommits_info_113_ldest = io_diffCommits_info_113_ldest;
        //    mon_tr.io_diffCommits_info_113_pdest = io_diffCommits_info_113_pdest;
        //    mon_tr.io_diffCommits_info_113_rfWen = io_diffCommits_info_113_rfWen;
        //    mon_tr.io_diffCommits_info_113_fpWen = io_diffCommits_info_113_fpWen;
        //    mon_tr.io_diffCommits_info_113_vecWen = io_diffCommits_info_113_vecWen;
        //    mon_tr.io_diffCommits_info_113_v0Wen = io_diffCommits_info_113_v0Wen;
        //    mon_tr.io_diffCommits_info_113_vlWen = io_diffCommits_info_113_vlWen;
        //    mon_tr.io_diffCommits_info_114_ldest = io_diffCommits_info_114_ldest;
        //    mon_tr.io_diffCommits_info_114_pdest = io_diffCommits_info_114_pdest;
        //    mon_tr.io_diffCommits_info_114_rfWen = io_diffCommits_info_114_rfWen;
        //    mon_tr.io_diffCommits_info_114_fpWen = io_diffCommits_info_114_fpWen;
        //    mon_tr.io_diffCommits_info_114_vecWen = io_diffCommits_info_114_vecWen;
        //    mon_tr.io_diffCommits_info_114_v0Wen = io_diffCommits_info_114_v0Wen;
        //    mon_tr.io_diffCommits_info_114_vlWen = io_diffCommits_info_114_vlWen;
        //    mon_tr.io_diffCommits_info_115_ldest = io_diffCommits_info_115_ldest;
        //    mon_tr.io_diffCommits_info_115_pdest = io_diffCommits_info_115_pdest;
        //    mon_tr.io_diffCommits_info_115_rfWen = io_diffCommits_info_115_rfWen;
        //    mon_tr.io_diffCommits_info_115_fpWen = io_diffCommits_info_115_fpWen;
        //    mon_tr.io_diffCommits_info_115_vecWen = io_diffCommits_info_115_vecWen;
        //    mon_tr.io_diffCommits_info_115_v0Wen = io_diffCommits_info_115_v0Wen;
        //    mon_tr.io_diffCommits_info_115_vlWen = io_diffCommits_info_115_vlWen;
        //    mon_tr.io_diffCommits_info_116_ldest = io_diffCommits_info_116_ldest;
        //    mon_tr.io_diffCommits_info_116_pdest = io_diffCommits_info_116_pdest;
        //    mon_tr.io_diffCommits_info_116_rfWen = io_diffCommits_info_116_rfWen;
        //    mon_tr.io_diffCommits_info_116_fpWen = io_diffCommits_info_116_fpWen;
        //    mon_tr.io_diffCommits_info_116_vecWen = io_diffCommits_info_116_vecWen;
        //    mon_tr.io_diffCommits_info_116_v0Wen = io_diffCommits_info_116_v0Wen;
        //    mon_tr.io_diffCommits_info_116_vlWen = io_diffCommits_info_116_vlWen;
        //    mon_tr.io_diffCommits_info_117_ldest = io_diffCommits_info_117_ldest;
        //    mon_tr.io_diffCommits_info_117_pdest = io_diffCommits_info_117_pdest;
        //    mon_tr.io_diffCommits_info_117_rfWen = io_diffCommits_info_117_rfWen;
        //    mon_tr.io_diffCommits_info_117_fpWen = io_diffCommits_info_117_fpWen;
        //    mon_tr.io_diffCommits_info_117_vecWen = io_diffCommits_info_117_vecWen;
        //    mon_tr.io_diffCommits_info_117_v0Wen = io_diffCommits_info_117_v0Wen;
        //    mon_tr.io_diffCommits_info_117_vlWen = io_diffCommits_info_117_vlWen;
        //    mon_tr.io_diffCommits_info_118_ldest = io_diffCommits_info_118_ldest;
        //    mon_tr.io_diffCommits_info_118_pdest = io_diffCommits_info_118_pdest;
        //    mon_tr.io_diffCommits_info_118_rfWen = io_diffCommits_info_118_rfWen;
        //    mon_tr.io_diffCommits_info_118_fpWen = io_diffCommits_info_118_fpWen;
        //    mon_tr.io_diffCommits_info_118_vecWen = io_diffCommits_info_118_vecWen;
        //    mon_tr.io_diffCommits_info_118_v0Wen = io_diffCommits_info_118_v0Wen;
        //    mon_tr.io_diffCommits_info_118_vlWen = io_diffCommits_info_118_vlWen;
        //    mon_tr.io_diffCommits_info_119_ldest = io_diffCommits_info_119_ldest;
        //    mon_tr.io_diffCommits_info_119_pdest = io_diffCommits_info_119_pdest;
        //    mon_tr.io_diffCommits_info_119_rfWen = io_diffCommits_info_119_rfWen;
        //    mon_tr.io_diffCommits_info_119_fpWen = io_diffCommits_info_119_fpWen;
        //    mon_tr.io_diffCommits_info_119_vecWen = io_diffCommits_info_119_vecWen;
        //    mon_tr.io_diffCommits_info_119_v0Wen = io_diffCommits_info_119_v0Wen;
        //    mon_tr.io_diffCommits_info_119_vlWen = io_diffCommits_info_119_vlWen;
        //    mon_tr.io_diffCommits_info_120_ldest = io_diffCommits_info_120_ldest;
        //    mon_tr.io_diffCommits_info_120_pdest = io_diffCommits_info_120_pdest;
        //    mon_tr.io_diffCommits_info_120_rfWen = io_diffCommits_info_120_rfWen;
        //    mon_tr.io_diffCommits_info_120_fpWen = io_diffCommits_info_120_fpWen;
        //    mon_tr.io_diffCommits_info_120_vecWen = io_diffCommits_info_120_vecWen;
        //    mon_tr.io_diffCommits_info_120_v0Wen = io_diffCommits_info_120_v0Wen;
        //    mon_tr.io_diffCommits_info_120_vlWen = io_diffCommits_info_120_vlWen;
        //    mon_tr.io_diffCommits_info_121_ldest = io_diffCommits_info_121_ldest;
        //    mon_tr.io_diffCommits_info_121_pdest = io_diffCommits_info_121_pdest;
        //    mon_tr.io_diffCommits_info_121_rfWen = io_diffCommits_info_121_rfWen;
        //    mon_tr.io_diffCommits_info_121_fpWen = io_diffCommits_info_121_fpWen;
        //    mon_tr.io_diffCommits_info_121_vecWen = io_diffCommits_info_121_vecWen;
        //    mon_tr.io_diffCommits_info_121_v0Wen = io_diffCommits_info_121_v0Wen;
        //    mon_tr.io_diffCommits_info_121_vlWen = io_diffCommits_info_121_vlWen;
        //    mon_tr.io_diffCommits_info_122_ldest = io_diffCommits_info_122_ldest;
        //    mon_tr.io_diffCommits_info_122_pdest = io_diffCommits_info_122_pdest;
        //    mon_tr.io_diffCommits_info_122_rfWen = io_diffCommits_info_122_rfWen;
        //    mon_tr.io_diffCommits_info_122_fpWen = io_diffCommits_info_122_fpWen;
        //    mon_tr.io_diffCommits_info_122_vecWen = io_diffCommits_info_122_vecWen;
        //    mon_tr.io_diffCommits_info_122_v0Wen = io_diffCommits_info_122_v0Wen;
        //    mon_tr.io_diffCommits_info_122_vlWen = io_diffCommits_info_122_vlWen;
        //    mon_tr.io_diffCommits_info_123_ldest = io_diffCommits_info_123_ldest;
        //    mon_tr.io_diffCommits_info_123_pdest = io_diffCommits_info_123_pdest;
        //    mon_tr.io_diffCommits_info_123_rfWen = io_diffCommits_info_123_rfWen;
        //    mon_tr.io_diffCommits_info_123_fpWen = io_diffCommits_info_123_fpWen;
        //    mon_tr.io_diffCommits_info_123_vecWen = io_diffCommits_info_123_vecWen;
        //    mon_tr.io_diffCommits_info_123_v0Wen = io_diffCommits_info_123_v0Wen;
        //    mon_tr.io_diffCommits_info_123_vlWen = io_diffCommits_info_123_vlWen;
        //    mon_tr.io_diffCommits_info_124_ldest = io_diffCommits_info_124_ldest;
        //    mon_tr.io_diffCommits_info_124_pdest = io_diffCommits_info_124_pdest;
        //    mon_tr.io_diffCommits_info_124_rfWen = io_diffCommits_info_124_rfWen;
        //    mon_tr.io_diffCommits_info_124_fpWen = io_diffCommits_info_124_fpWen;
        //    mon_tr.io_diffCommits_info_124_vecWen = io_diffCommits_info_124_vecWen;
        //    mon_tr.io_diffCommits_info_124_v0Wen = io_diffCommits_info_124_v0Wen;
        //    mon_tr.io_diffCommits_info_124_vlWen = io_diffCommits_info_124_vlWen;
        //    mon_tr.io_diffCommits_info_125_ldest = io_diffCommits_info_125_ldest;
        //    mon_tr.io_diffCommits_info_125_pdest = io_diffCommits_info_125_pdest;
        //    mon_tr.io_diffCommits_info_125_rfWen = io_diffCommits_info_125_rfWen;
        //    mon_tr.io_diffCommits_info_125_fpWen = io_diffCommits_info_125_fpWen;
        //    mon_tr.io_diffCommits_info_125_vecWen = io_diffCommits_info_125_vecWen;
        //    mon_tr.io_diffCommits_info_125_v0Wen = io_diffCommits_info_125_v0Wen;
        //    mon_tr.io_diffCommits_info_125_vlWen = io_diffCommits_info_125_vlWen;
        //    mon_tr.io_diffCommits_info_126_ldest = io_diffCommits_info_126_ldest;
        //    mon_tr.io_diffCommits_info_126_pdest = io_diffCommits_info_126_pdest;
        //    mon_tr.io_diffCommits_info_126_rfWen = io_diffCommits_info_126_rfWen;
        //    mon_tr.io_diffCommits_info_126_fpWen = io_diffCommits_info_126_fpWen;
        //    mon_tr.io_diffCommits_info_126_vecWen = io_diffCommits_info_126_vecWen;
        //    mon_tr.io_diffCommits_info_126_v0Wen = io_diffCommits_info_126_v0Wen;
        //    mon_tr.io_diffCommits_info_126_vlWen = io_diffCommits_info_126_vlWen;
        //    mon_tr.io_diffCommits_info_127_ldest = io_diffCommits_info_127_ldest;
        //    mon_tr.io_diffCommits_info_127_pdest = io_diffCommits_info_127_pdest;
        //    mon_tr.io_diffCommits_info_127_rfWen = io_diffCommits_info_127_rfWen;
        //    mon_tr.io_diffCommits_info_127_fpWen = io_diffCommits_info_127_fpWen;
        //    mon_tr.io_diffCommits_info_127_vecWen = io_diffCommits_info_127_vecWen;
        //    mon_tr.io_diffCommits_info_127_v0Wen = io_diffCommits_info_127_v0Wen;
        //    mon_tr.io_diffCommits_info_127_vlWen = io_diffCommits_info_127_vlWen;
        //    mon_tr.io_diffCommits_info_128_ldest = io_diffCommits_info_128_ldest;
        //    mon_tr.io_diffCommits_info_128_pdest = io_diffCommits_info_128_pdest;
        //    mon_tr.io_diffCommits_info_128_rfWen = io_diffCommits_info_128_rfWen;
        //    mon_tr.io_diffCommits_info_128_fpWen = io_diffCommits_info_128_fpWen;
        //    mon_tr.io_diffCommits_info_128_vecWen = io_diffCommits_info_128_vecWen;
        //    mon_tr.io_diffCommits_info_128_v0Wen = io_diffCommits_info_128_v0Wen;
        //    mon_tr.io_diffCommits_info_128_vlWen = io_diffCommits_info_128_vlWen;
        //    mon_tr.io_diffCommits_info_129_ldest = io_diffCommits_info_129_ldest;
        //    mon_tr.io_diffCommits_info_129_pdest = io_diffCommits_info_129_pdest;
        //    mon_tr.io_diffCommits_info_129_rfWen = io_diffCommits_info_129_rfWen;
        //    mon_tr.io_diffCommits_info_129_fpWen = io_diffCommits_info_129_fpWen;
        //    mon_tr.io_diffCommits_info_129_vecWen = io_diffCommits_info_129_vecWen;
        //    mon_tr.io_diffCommits_info_129_v0Wen = io_diffCommits_info_129_v0Wen;
        //    mon_tr.io_diffCommits_info_129_vlWen = io_diffCommits_info_129_vlWen;
        //    mon_tr.io_diffCommits_info_130_ldest = io_diffCommits_info_130_ldest;
        //    mon_tr.io_diffCommits_info_130_pdest = io_diffCommits_info_130_pdest;
        //    mon_tr.io_diffCommits_info_130_rfWen = io_diffCommits_info_130_rfWen;
        //    mon_tr.io_diffCommits_info_130_fpWen = io_diffCommits_info_130_fpWen;
        //    mon_tr.io_diffCommits_info_130_vecWen = io_diffCommits_info_130_vecWen;
        //    mon_tr.io_diffCommits_info_130_v0Wen = io_diffCommits_info_130_v0Wen;
        //    mon_tr.io_diffCommits_info_130_vlWen = io_diffCommits_info_130_vlWen;
        //    mon_tr.io_diffCommits_info_131_ldest = io_diffCommits_info_131_ldest;
        //    mon_tr.io_diffCommits_info_131_pdest = io_diffCommits_info_131_pdest;
        //    mon_tr.io_diffCommits_info_131_rfWen = io_diffCommits_info_131_rfWen;
        //    mon_tr.io_diffCommits_info_131_fpWen = io_diffCommits_info_131_fpWen;
        //    mon_tr.io_diffCommits_info_131_vecWen = io_diffCommits_info_131_vecWen;
        //    mon_tr.io_diffCommits_info_131_v0Wen = io_diffCommits_info_131_v0Wen;
        //    mon_tr.io_diffCommits_info_131_vlWen = io_diffCommits_info_131_vlWen;
        //    mon_tr.io_diffCommits_info_132_ldest = io_diffCommits_info_132_ldest;
        //    mon_tr.io_diffCommits_info_132_pdest = io_diffCommits_info_132_pdest;
        //    mon_tr.io_diffCommits_info_132_rfWen = io_diffCommits_info_132_rfWen;
        //    mon_tr.io_diffCommits_info_132_fpWen = io_diffCommits_info_132_fpWen;
        //    mon_tr.io_diffCommits_info_132_vecWen = io_diffCommits_info_132_vecWen;
        //    mon_tr.io_diffCommits_info_132_v0Wen = io_diffCommits_info_132_v0Wen;
        //    mon_tr.io_diffCommits_info_132_vlWen = io_diffCommits_info_132_vlWen;
        //    mon_tr.io_diffCommits_info_133_ldest = io_diffCommits_info_133_ldest;
        //    mon_tr.io_diffCommits_info_133_pdest = io_diffCommits_info_133_pdest;
        //    mon_tr.io_diffCommits_info_133_rfWen = io_diffCommits_info_133_rfWen;
        //    mon_tr.io_diffCommits_info_133_fpWen = io_diffCommits_info_133_fpWen;
        //    mon_tr.io_diffCommits_info_133_vecWen = io_diffCommits_info_133_vecWen;
        //    mon_tr.io_diffCommits_info_133_v0Wen = io_diffCommits_info_133_v0Wen;
        //    mon_tr.io_diffCommits_info_133_vlWen = io_diffCommits_info_133_vlWen;
        //    mon_tr.io_diffCommits_info_134_ldest = io_diffCommits_info_134_ldest;
        //    mon_tr.io_diffCommits_info_134_pdest = io_diffCommits_info_134_pdest;
        //    mon_tr.io_diffCommits_info_134_rfWen = io_diffCommits_info_134_rfWen;
        //    mon_tr.io_diffCommits_info_134_fpWen = io_diffCommits_info_134_fpWen;
        //    mon_tr.io_diffCommits_info_134_vecWen = io_diffCommits_info_134_vecWen;
        //    mon_tr.io_diffCommits_info_134_v0Wen = io_diffCommits_info_134_v0Wen;
        //    mon_tr.io_diffCommits_info_134_vlWen = io_diffCommits_info_134_vlWen;
        //    mon_tr.io_diffCommits_info_135_ldest = io_diffCommits_info_135_ldest;
        //    mon_tr.io_diffCommits_info_135_pdest = io_diffCommits_info_135_pdest;
        //    mon_tr.io_diffCommits_info_135_rfWen = io_diffCommits_info_135_rfWen;
        //    mon_tr.io_diffCommits_info_135_fpWen = io_diffCommits_info_135_fpWen;
        //    mon_tr.io_diffCommits_info_135_vecWen = io_diffCommits_info_135_vecWen;
        //    mon_tr.io_diffCommits_info_135_v0Wen = io_diffCommits_info_135_v0Wen;
        //    mon_tr.io_diffCommits_info_135_vlWen = io_diffCommits_info_135_vlWen;
        //    mon_tr.io_diffCommits_info_136_ldest = io_diffCommits_info_136_ldest;
        //    mon_tr.io_diffCommits_info_136_pdest = io_diffCommits_info_136_pdest;
        //    mon_tr.io_diffCommits_info_136_rfWen = io_diffCommits_info_136_rfWen;
        //    mon_tr.io_diffCommits_info_136_fpWen = io_diffCommits_info_136_fpWen;
        //    mon_tr.io_diffCommits_info_136_vecWen = io_diffCommits_info_136_vecWen;
        //    mon_tr.io_diffCommits_info_136_v0Wen = io_diffCommits_info_136_v0Wen;
        //    mon_tr.io_diffCommits_info_136_vlWen = io_diffCommits_info_136_vlWen;
        //    mon_tr.io_diffCommits_info_137_ldest = io_diffCommits_info_137_ldest;
        //    mon_tr.io_diffCommits_info_137_pdest = io_diffCommits_info_137_pdest;
        //    mon_tr.io_diffCommits_info_137_rfWen = io_diffCommits_info_137_rfWen;
        //    mon_tr.io_diffCommits_info_137_fpWen = io_diffCommits_info_137_fpWen;
        //    mon_tr.io_diffCommits_info_137_vecWen = io_diffCommits_info_137_vecWen;
        //    mon_tr.io_diffCommits_info_137_v0Wen = io_diffCommits_info_137_v0Wen;
        //    mon_tr.io_diffCommits_info_137_vlWen = io_diffCommits_info_137_vlWen;
        //    mon_tr.io_diffCommits_info_138_ldest = io_diffCommits_info_138_ldest;
        //    mon_tr.io_diffCommits_info_138_pdest = io_diffCommits_info_138_pdest;
        //    mon_tr.io_diffCommits_info_138_rfWen = io_diffCommits_info_138_rfWen;
        //    mon_tr.io_diffCommits_info_138_fpWen = io_diffCommits_info_138_fpWen;
        //    mon_tr.io_diffCommits_info_138_vecWen = io_diffCommits_info_138_vecWen;
        //    mon_tr.io_diffCommits_info_138_v0Wen = io_diffCommits_info_138_v0Wen;
        //    mon_tr.io_diffCommits_info_138_vlWen = io_diffCommits_info_138_vlWen;
        //    mon_tr.io_diffCommits_info_139_ldest = io_diffCommits_info_139_ldest;
        //    mon_tr.io_diffCommits_info_139_pdest = io_diffCommits_info_139_pdest;
        //    mon_tr.io_diffCommits_info_139_rfWen = io_diffCommits_info_139_rfWen;
        //    mon_tr.io_diffCommits_info_139_fpWen = io_diffCommits_info_139_fpWen;
        //    mon_tr.io_diffCommits_info_139_vecWen = io_diffCommits_info_139_vecWen;
        //    mon_tr.io_diffCommits_info_139_v0Wen = io_diffCommits_info_139_v0Wen;
        //    mon_tr.io_diffCommits_info_139_vlWen = io_diffCommits_info_139_vlWen;
        //    mon_tr.io_diffCommits_info_140_ldest = io_diffCommits_info_140_ldest;
        //    mon_tr.io_diffCommits_info_140_pdest = io_diffCommits_info_140_pdest;
        //    mon_tr.io_diffCommits_info_140_rfWen = io_diffCommits_info_140_rfWen;
        //    mon_tr.io_diffCommits_info_140_fpWen = io_diffCommits_info_140_fpWen;
        //    mon_tr.io_diffCommits_info_140_vecWen = io_diffCommits_info_140_vecWen;
        //    mon_tr.io_diffCommits_info_140_v0Wen = io_diffCommits_info_140_v0Wen;
        //    mon_tr.io_diffCommits_info_140_vlWen = io_diffCommits_info_140_vlWen;
        //    mon_tr.io_diffCommits_info_141_ldest = io_diffCommits_info_141_ldest;
        //    mon_tr.io_diffCommits_info_141_pdest = io_diffCommits_info_141_pdest;
        //    mon_tr.io_diffCommits_info_141_rfWen = io_diffCommits_info_141_rfWen;
        //    mon_tr.io_diffCommits_info_141_fpWen = io_diffCommits_info_141_fpWen;
        //    mon_tr.io_diffCommits_info_141_vecWen = io_diffCommits_info_141_vecWen;
        //    mon_tr.io_diffCommits_info_141_v0Wen = io_diffCommits_info_141_v0Wen;
        //    mon_tr.io_diffCommits_info_141_vlWen = io_diffCommits_info_141_vlWen;
        //    mon_tr.io_diffCommits_info_142_ldest = io_diffCommits_info_142_ldest;
        //    mon_tr.io_diffCommits_info_142_pdest = io_diffCommits_info_142_pdest;
        //    mon_tr.io_diffCommits_info_142_rfWen = io_diffCommits_info_142_rfWen;
        //    mon_tr.io_diffCommits_info_142_fpWen = io_diffCommits_info_142_fpWen;
        //    mon_tr.io_diffCommits_info_142_vecWen = io_diffCommits_info_142_vecWen;
        //    mon_tr.io_diffCommits_info_142_v0Wen = io_diffCommits_info_142_v0Wen;
        //    mon_tr.io_diffCommits_info_142_vlWen = io_diffCommits_info_142_vlWen;
        //    mon_tr.io_diffCommits_info_143_ldest = io_diffCommits_info_143_ldest;
        //    mon_tr.io_diffCommits_info_143_pdest = io_diffCommits_info_143_pdest;
        //    mon_tr.io_diffCommits_info_143_rfWen = io_diffCommits_info_143_rfWen;
        //    mon_tr.io_diffCommits_info_143_fpWen = io_diffCommits_info_143_fpWen;
        //    mon_tr.io_diffCommits_info_143_vecWen = io_diffCommits_info_143_vecWen;
        //    mon_tr.io_diffCommits_info_143_v0Wen = io_diffCommits_info_143_v0Wen;
        //    mon_tr.io_diffCommits_info_143_vlWen = io_diffCommits_info_143_vlWen;
        //    mon_tr.io_diffCommits_info_144_ldest = io_diffCommits_info_144_ldest;
        //    mon_tr.io_diffCommits_info_144_pdest = io_diffCommits_info_144_pdest;
        //    mon_tr.io_diffCommits_info_144_rfWen = io_diffCommits_info_144_rfWen;
        //    mon_tr.io_diffCommits_info_144_fpWen = io_diffCommits_info_144_fpWen;
        //    mon_tr.io_diffCommits_info_144_vecWen = io_diffCommits_info_144_vecWen;
        //    mon_tr.io_diffCommits_info_144_v0Wen = io_diffCommits_info_144_v0Wen;
        //    mon_tr.io_diffCommits_info_144_vlWen = io_diffCommits_info_144_vlWen;
        //    mon_tr.io_diffCommits_info_145_ldest = io_diffCommits_info_145_ldest;
        //    mon_tr.io_diffCommits_info_145_pdest = io_diffCommits_info_145_pdest;
        //    mon_tr.io_diffCommits_info_145_rfWen = io_diffCommits_info_145_rfWen;
        //    mon_tr.io_diffCommits_info_145_fpWen = io_diffCommits_info_145_fpWen;
        //    mon_tr.io_diffCommits_info_145_vecWen = io_diffCommits_info_145_vecWen;
        //    mon_tr.io_diffCommits_info_145_v0Wen = io_diffCommits_info_145_v0Wen;
        //    mon_tr.io_diffCommits_info_145_vlWen = io_diffCommits_info_145_vlWen;
        //    mon_tr.io_diffCommits_info_146_ldest = io_diffCommits_info_146_ldest;
        //    mon_tr.io_diffCommits_info_146_pdest = io_diffCommits_info_146_pdest;
        //    mon_tr.io_diffCommits_info_146_rfWen = io_diffCommits_info_146_rfWen;
        //    mon_tr.io_diffCommits_info_146_fpWen = io_diffCommits_info_146_fpWen;
        //    mon_tr.io_diffCommits_info_146_vecWen = io_diffCommits_info_146_vecWen;
        //    mon_tr.io_diffCommits_info_146_v0Wen = io_diffCommits_info_146_v0Wen;
        //    mon_tr.io_diffCommits_info_146_vlWen = io_diffCommits_info_146_vlWen;
        //    mon_tr.io_diffCommits_info_147_ldest = io_diffCommits_info_147_ldest;
        //    mon_tr.io_diffCommits_info_147_pdest = io_diffCommits_info_147_pdest;
        //    mon_tr.io_diffCommits_info_147_rfWen = io_diffCommits_info_147_rfWen;
        //    mon_tr.io_diffCommits_info_147_fpWen = io_diffCommits_info_147_fpWen;
        //    mon_tr.io_diffCommits_info_147_vecWen = io_diffCommits_info_147_vecWen;
        //    mon_tr.io_diffCommits_info_147_v0Wen = io_diffCommits_info_147_v0Wen;
        //    mon_tr.io_diffCommits_info_147_vlWen = io_diffCommits_info_147_vlWen;
        //    mon_tr.io_diffCommits_info_148_ldest = io_diffCommits_info_148_ldest;
        //    mon_tr.io_diffCommits_info_148_pdest = io_diffCommits_info_148_pdest;
        //    mon_tr.io_diffCommits_info_148_rfWen = io_diffCommits_info_148_rfWen;
        //    mon_tr.io_diffCommits_info_148_fpWen = io_diffCommits_info_148_fpWen;
        //    mon_tr.io_diffCommits_info_148_vecWen = io_diffCommits_info_148_vecWen;
        //    mon_tr.io_diffCommits_info_148_v0Wen = io_diffCommits_info_148_v0Wen;
        //    mon_tr.io_diffCommits_info_148_vlWen = io_diffCommits_info_148_vlWen;
        //    mon_tr.io_diffCommits_info_149_ldest = io_diffCommits_info_149_ldest;
        //    mon_tr.io_diffCommits_info_149_pdest = io_diffCommits_info_149_pdest;
        //    mon_tr.io_diffCommits_info_149_rfWen = io_diffCommits_info_149_rfWen;
        //    mon_tr.io_diffCommits_info_149_fpWen = io_diffCommits_info_149_fpWen;
        //    mon_tr.io_diffCommits_info_149_vecWen = io_diffCommits_info_149_vecWen;
        //    mon_tr.io_diffCommits_info_149_v0Wen = io_diffCommits_info_149_v0Wen;
        //    mon_tr.io_diffCommits_info_149_vlWen = io_diffCommits_info_149_vlWen;
        //    mon_tr.io_diffCommits_info_150_ldest = io_diffCommits_info_150_ldest;
        //    mon_tr.io_diffCommits_info_150_pdest = io_diffCommits_info_150_pdest;
        //    mon_tr.io_diffCommits_info_150_rfWen = io_diffCommits_info_150_rfWen;
        //    mon_tr.io_diffCommits_info_150_fpWen = io_diffCommits_info_150_fpWen;
        //    mon_tr.io_diffCommits_info_150_vecWen = io_diffCommits_info_150_vecWen;
        //    mon_tr.io_diffCommits_info_150_v0Wen = io_diffCommits_info_150_v0Wen;
        //    mon_tr.io_diffCommits_info_150_vlWen = io_diffCommits_info_150_vlWen;
        //    mon_tr.io_diffCommits_info_151_ldest = io_diffCommits_info_151_ldest;
        //    mon_tr.io_diffCommits_info_151_pdest = io_diffCommits_info_151_pdest;
        //    mon_tr.io_diffCommits_info_151_rfWen = io_diffCommits_info_151_rfWen;
        //    mon_tr.io_diffCommits_info_151_fpWen = io_diffCommits_info_151_fpWen;
        //    mon_tr.io_diffCommits_info_151_vecWen = io_diffCommits_info_151_vecWen;
        //    mon_tr.io_diffCommits_info_151_v0Wen = io_diffCommits_info_151_v0Wen;
        //    mon_tr.io_diffCommits_info_151_vlWen = io_diffCommits_info_151_vlWen;
        //    mon_tr.io_diffCommits_info_152_ldest = io_diffCommits_info_152_ldest;
        //    mon_tr.io_diffCommits_info_152_pdest = io_diffCommits_info_152_pdest;
        //    mon_tr.io_diffCommits_info_152_rfWen = io_diffCommits_info_152_rfWen;
        //    mon_tr.io_diffCommits_info_152_fpWen = io_diffCommits_info_152_fpWen;
        //    mon_tr.io_diffCommits_info_152_vecWen = io_diffCommits_info_152_vecWen;
        //    mon_tr.io_diffCommits_info_152_v0Wen = io_diffCommits_info_152_v0Wen;
        //    mon_tr.io_diffCommits_info_152_vlWen = io_diffCommits_info_152_vlWen;
        //    mon_tr.io_diffCommits_info_153_ldest = io_diffCommits_info_153_ldest;
        //    mon_tr.io_diffCommits_info_153_pdest = io_diffCommits_info_153_pdest;
        //    mon_tr.io_diffCommits_info_153_rfWen = io_diffCommits_info_153_rfWen;
        //    mon_tr.io_diffCommits_info_153_fpWen = io_diffCommits_info_153_fpWen;
        //    mon_tr.io_diffCommits_info_153_vecWen = io_diffCommits_info_153_vecWen;
        //    mon_tr.io_diffCommits_info_153_v0Wen = io_diffCommits_info_153_v0Wen;
        //    mon_tr.io_diffCommits_info_153_vlWen = io_diffCommits_info_153_vlWen;
        //    mon_tr.io_diffCommits_info_154_ldest = io_diffCommits_info_154_ldest;
        //    mon_tr.io_diffCommits_info_154_pdest = io_diffCommits_info_154_pdest;
        //    mon_tr.io_diffCommits_info_154_rfWen = io_diffCommits_info_154_rfWen;
        //    mon_tr.io_diffCommits_info_154_fpWen = io_diffCommits_info_154_fpWen;
        //    mon_tr.io_diffCommits_info_154_vecWen = io_diffCommits_info_154_vecWen;
        //    mon_tr.io_diffCommits_info_154_v0Wen = io_diffCommits_info_154_v0Wen;
        //    mon_tr.io_diffCommits_info_154_vlWen = io_diffCommits_info_154_vlWen;
        //    mon_tr.io_diffCommits_info_155_ldest = io_diffCommits_info_155_ldest;
        //    mon_tr.io_diffCommits_info_155_pdest = io_diffCommits_info_155_pdest;
        //    mon_tr.io_diffCommits_info_155_rfWen = io_diffCommits_info_155_rfWen;
        //    mon_tr.io_diffCommits_info_155_fpWen = io_diffCommits_info_155_fpWen;
        //    mon_tr.io_diffCommits_info_155_vecWen = io_diffCommits_info_155_vecWen;
        //    mon_tr.io_diffCommits_info_155_v0Wen = io_diffCommits_info_155_v0Wen;
        //    mon_tr.io_diffCommits_info_155_vlWen = io_diffCommits_info_155_vlWen;
        //    mon_tr.io_diffCommits_info_156_ldest = io_diffCommits_info_156_ldest;
        //    mon_tr.io_diffCommits_info_156_pdest = io_diffCommits_info_156_pdest;
        //    mon_tr.io_diffCommits_info_156_rfWen = io_diffCommits_info_156_rfWen;
        //    mon_tr.io_diffCommits_info_156_fpWen = io_diffCommits_info_156_fpWen;
        //    mon_tr.io_diffCommits_info_156_vecWen = io_diffCommits_info_156_vecWen;
        //    mon_tr.io_diffCommits_info_156_v0Wen = io_diffCommits_info_156_v0Wen;
        //    mon_tr.io_diffCommits_info_156_vlWen = io_diffCommits_info_156_vlWen;
        //    mon_tr.io_diffCommits_info_157_ldest = io_diffCommits_info_157_ldest;
        //    mon_tr.io_diffCommits_info_157_pdest = io_diffCommits_info_157_pdest;
        //    mon_tr.io_diffCommits_info_157_rfWen = io_diffCommits_info_157_rfWen;
        //    mon_tr.io_diffCommits_info_157_fpWen = io_diffCommits_info_157_fpWen;
        //    mon_tr.io_diffCommits_info_157_vecWen = io_diffCommits_info_157_vecWen;
        //    mon_tr.io_diffCommits_info_157_v0Wen = io_diffCommits_info_157_v0Wen;
        //    mon_tr.io_diffCommits_info_157_vlWen = io_diffCommits_info_157_vlWen;
        //    mon_tr.io_diffCommits_info_158_ldest = io_diffCommits_info_158_ldest;
        //    mon_tr.io_diffCommits_info_158_pdest = io_diffCommits_info_158_pdest;
        //    mon_tr.io_diffCommits_info_158_rfWen = io_diffCommits_info_158_rfWen;
        //    mon_tr.io_diffCommits_info_158_fpWen = io_diffCommits_info_158_fpWen;
        //    mon_tr.io_diffCommits_info_158_vecWen = io_diffCommits_info_158_vecWen;
        //    mon_tr.io_diffCommits_info_158_v0Wen = io_diffCommits_info_158_v0Wen;
        //    mon_tr.io_diffCommits_info_158_vlWen = io_diffCommits_info_158_vlWen;
        //    mon_tr.io_diffCommits_info_159_ldest = io_diffCommits_info_159_ldest;
        //    mon_tr.io_diffCommits_info_159_pdest = io_diffCommits_info_159_pdest;
        //    mon_tr.io_diffCommits_info_159_rfWen = io_diffCommits_info_159_rfWen;
        //    mon_tr.io_diffCommits_info_159_fpWen = io_diffCommits_info_159_fpWen;
        //    mon_tr.io_diffCommits_info_159_vecWen = io_diffCommits_info_159_vecWen;
        //    mon_tr.io_diffCommits_info_159_v0Wen = io_diffCommits_info_159_v0Wen;
        //    mon_tr.io_diffCommits_info_159_vlWen = io_diffCommits_info_159_vlWen;
        //    mon_tr.io_diffCommits_info_160_ldest = io_diffCommits_info_160_ldest;
        //    mon_tr.io_diffCommits_info_160_pdest = io_diffCommits_info_160_pdest;
        //    mon_tr.io_diffCommits_info_160_rfWen = io_diffCommits_info_160_rfWen;
        //    mon_tr.io_diffCommits_info_160_fpWen = io_diffCommits_info_160_fpWen;
        //    mon_tr.io_diffCommits_info_160_vecWen = io_diffCommits_info_160_vecWen;
        //    mon_tr.io_diffCommits_info_160_v0Wen = io_diffCommits_info_160_v0Wen;
        //    mon_tr.io_diffCommits_info_160_vlWen = io_diffCommits_info_160_vlWen;
        //    mon_tr.io_diffCommits_info_161_ldest = io_diffCommits_info_161_ldest;
        //    mon_tr.io_diffCommits_info_161_pdest = io_diffCommits_info_161_pdest;
        //    mon_tr.io_diffCommits_info_161_rfWen = io_diffCommits_info_161_rfWen;
        //    mon_tr.io_diffCommits_info_161_fpWen = io_diffCommits_info_161_fpWen;
        //    mon_tr.io_diffCommits_info_161_vecWen = io_diffCommits_info_161_vecWen;
        //    mon_tr.io_diffCommits_info_161_v0Wen = io_diffCommits_info_161_v0Wen;
        //    mon_tr.io_diffCommits_info_161_vlWen = io_diffCommits_info_161_vlWen;
        //    mon_tr.io_diffCommits_info_162_ldest = io_diffCommits_info_162_ldest;
        //    mon_tr.io_diffCommits_info_162_pdest = io_diffCommits_info_162_pdest;
        //    mon_tr.io_diffCommits_info_162_rfWen = io_diffCommits_info_162_rfWen;
        //    mon_tr.io_diffCommits_info_162_fpWen = io_diffCommits_info_162_fpWen;
        //    mon_tr.io_diffCommits_info_162_vecWen = io_diffCommits_info_162_vecWen;
        //    mon_tr.io_diffCommits_info_162_v0Wen = io_diffCommits_info_162_v0Wen;
        //    mon_tr.io_diffCommits_info_162_vlWen = io_diffCommits_info_162_vlWen;
        //    mon_tr.io_diffCommits_info_163_ldest = io_diffCommits_info_163_ldest;
        //    mon_tr.io_diffCommits_info_163_pdest = io_diffCommits_info_163_pdest;
        //    mon_tr.io_diffCommits_info_163_rfWen = io_diffCommits_info_163_rfWen;
        //    mon_tr.io_diffCommits_info_163_fpWen = io_diffCommits_info_163_fpWen;
        //    mon_tr.io_diffCommits_info_163_vecWen = io_diffCommits_info_163_vecWen;
        //    mon_tr.io_diffCommits_info_163_v0Wen = io_diffCommits_info_163_v0Wen;
        //    mon_tr.io_diffCommits_info_163_vlWen = io_diffCommits_info_163_vlWen;
        //    mon_tr.io_diffCommits_info_164_ldest = io_diffCommits_info_164_ldest;
        //    mon_tr.io_diffCommits_info_164_pdest = io_diffCommits_info_164_pdest;
        //    mon_tr.io_diffCommits_info_164_rfWen = io_diffCommits_info_164_rfWen;
        //    mon_tr.io_diffCommits_info_164_fpWen = io_diffCommits_info_164_fpWen;
        //    mon_tr.io_diffCommits_info_164_vecWen = io_diffCommits_info_164_vecWen;
        //    mon_tr.io_diffCommits_info_164_v0Wen = io_diffCommits_info_164_v0Wen;
        //    mon_tr.io_diffCommits_info_164_vlWen = io_diffCommits_info_164_vlWen;
        //    mon_tr.io_diffCommits_info_165_ldest = io_diffCommits_info_165_ldest;
        //    mon_tr.io_diffCommits_info_165_pdest = io_diffCommits_info_165_pdest;
        //    mon_tr.io_diffCommits_info_165_rfWen = io_diffCommits_info_165_rfWen;
        //    mon_tr.io_diffCommits_info_165_fpWen = io_diffCommits_info_165_fpWen;
        //    mon_tr.io_diffCommits_info_165_vecWen = io_diffCommits_info_165_vecWen;
        //    mon_tr.io_diffCommits_info_165_v0Wen = io_diffCommits_info_165_v0Wen;
        //    mon_tr.io_diffCommits_info_165_vlWen = io_diffCommits_info_165_vlWen;
        //    mon_tr.io_diffCommits_info_166_ldest = io_diffCommits_info_166_ldest;
        //    mon_tr.io_diffCommits_info_166_pdest = io_diffCommits_info_166_pdest;
        //    mon_tr.io_diffCommits_info_166_rfWen = io_diffCommits_info_166_rfWen;
        //    mon_tr.io_diffCommits_info_166_fpWen = io_diffCommits_info_166_fpWen;
        //    mon_tr.io_diffCommits_info_166_vecWen = io_diffCommits_info_166_vecWen;
        //    mon_tr.io_diffCommits_info_166_v0Wen = io_diffCommits_info_166_v0Wen;
        //    mon_tr.io_diffCommits_info_166_vlWen = io_diffCommits_info_166_vlWen;
        //    mon_tr.io_diffCommits_info_167_ldest = io_diffCommits_info_167_ldest;
        //    mon_tr.io_diffCommits_info_167_pdest = io_diffCommits_info_167_pdest;
        //    mon_tr.io_diffCommits_info_167_rfWen = io_diffCommits_info_167_rfWen;
        //    mon_tr.io_diffCommits_info_167_fpWen = io_diffCommits_info_167_fpWen;
        //    mon_tr.io_diffCommits_info_167_vecWen = io_diffCommits_info_167_vecWen;
        //    mon_tr.io_diffCommits_info_167_v0Wen = io_diffCommits_info_167_v0Wen;
        //    mon_tr.io_diffCommits_info_167_vlWen = io_diffCommits_info_167_vlWen;
        //    mon_tr.io_diffCommits_info_168_ldest = io_diffCommits_info_168_ldest;
        //    mon_tr.io_diffCommits_info_168_pdest = io_diffCommits_info_168_pdest;
        //    mon_tr.io_diffCommits_info_168_rfWen = io_diffCommits_info_168_rfWen;
        //    mon_tr.io_diffCommits_info_168_fpWen = io_diffCommits_info_168_fpWen;
        //    mon_tr.io_diffCommits_info_168_vecWen = io_diffCommits_info_168_vecWen;
        //    mon_tr.io_diffCommits_info_168_v0Wen = io_diffCommits_info_168_v0Wen;
        //    mon_tr.io_diffCommits_info_168_vlWen = io_diffCommits_info_168_vlWen;
        //    mon_tr.io_diffCommits_info_169_ldest = io_diffCommits_info_169_ldest;
        //    mon_tr.io_diffCommits_info_169_pdest = io_diffCommits_info_169_pdest;
        //    mon_tr.io_diffCommits_info_169_rfWen = io_diffCommits_info_169_rfWen;
        //    mon_tr.io_diffCommits_info_169_fpWen = io_diffCommits_info_169_fpWen;
        //    mon_tr.io_diffCommits_info_169_vecWen = io_diffCommits_info_169_vecWen;
        //    mon_tr.io_diffCommits_info_169_v0Wen = io_diffCommits_info_169_v0Wen;
        //    mon_tr.io_diffCommits_info_169_vlWen = io_diffCommits_info_169_vlWen;
        //    mon_tr.io_diffCommits_info_170_ldest = io_diffCommits_info_170_ldest;
        //    mon_tr.io_diffCommits_info_170_pdest = io_diffCommits_info_170_pdest;
        //    mon_tr.io_diffCommits_info_170_rfWen = io_diffCommits_info_170_rfWen;
        //    mon_tr.io_diffCommits_info_170_fpWen = io_diffCommits_info_170_fpWen;
        //    mon_tr.io_diffCommits_info_170_vecWen = io_diffCommits_info_170_vecWen;
        //    mon_tr.io_diffCommits_info_170_v0Wen = io_diffCommits_info_170_v0Wen;
        //    mon_tr.io_diffCommits_info_170_vlWen = io_diffCommits_info_170_vlWen;
        //    mon_tr.io_diffCommits_info_171_ldest = io_diffCommits_info_171_ldest;
        //    mon_tr.io_diffCommits_info_171_pdest = io_diffCommits_info_171_pdest;
        //    mon_tr.io_diffCommits_info_171_rfWen = io_diffCommits_info_171_rfWen;
        //    mon_tr.io_diffCommits_info_171_fpWen = io_diffCommits_info_171_fpWen;
        //    mon_tr.io_diffCommits_info_171_vecWen = io_diffCommits_info_171_vecWen;
        //    mon_tr.io_diffCommits_info_171_v0Wen = io_diffCommits_info_171_v0Wen;
        //    mon_tr.io_diffCommits_info_171_vlWen = io_diffCommits_info_171_vlWen;
        //    mon_tr.io_diffCommits_info_172_ldest = io_diffCommits_info_172_ldest;
        //    mon_tr.io_diffCommits_info_172_pdest = io_diffCommits_info_172_pdest;
        //    mon_tr.io_diffCommits_info_172_rfWen = io_diffCommits_info_172_rfWen;
        //    mon_tr.io_diffCommits_info_172_fpWen = io_diffCommits_info_172_fpWen;
        //    mon_tr.io_diffCommits_info_172_vecWen = io_diffCommits_info_172_vecWen;
        //    mon_tr.io_diffCommits_info_172_v0Wen = io_diffCommits_info_172_v0Wen;
        //    mon_tr.io_diffCommits_info_172_vlWen = io_diffCommits_info_172_vlWen;
        //    mon_tr.io_diffCommits_info_173_ldest = io_diffCommits_info_173_ldest;
        //    mon_tr.io_diffCommits_info_173_pdest = io_diffCommits_info_173_pdest;
        //    mon_tr.io_diffCommits_info_173_rfWen = io_diffCommits_info_173_rfWen;
        //    mon_tr.io_diffCommits_info_173_fpWen = io_diffCommits_info_173_fpWen;
        //    mon_tr.io_diffCommits_info_173_vecWen = io_diffCommits_info_173_vecWen;
        //    mon_tr.io_diffCommits_info_173_v0Wen = io_diffCommits_info_173_v0Wen;
        //    mon_tr.io_diffCommits_info_173_vlWen = io_diffCommits_info_173_vlWen;
        //    mon_tr.io_diffCommits_info_174_ldest = io_diffCommits_info_174_ldest;
        //    mon_tr.io_diffCommits_info_174_pdest = io_diffCommits_info_174_pdest;
        //    mon_tr.io_diffCommits_info_174_rfWen = io_diffCommits_info_174_rfWen;
        //    mon_tr.io_diffCommits_info_174_fpWen = io_diffCommits_info_174_fpWen;
        //    mon_tr.io_diffCommits_info_174_vecWen = io_diffCommits_info_174_vecWen;
        //    mon_tr.io_diffCommits_info_174_v0Wen = io_diffCommits_info_174_v0Wen;
        //    mon_tr.io_diffCommits_info_174_vlWen = io_diffCommits_info_174_vlWen;
        //    mon_tr.io_diffCommits_info_175_ldest = io_diffCommits_info_175_ldest;
        //    mon_tr.io_diffCommits_info_175_pdest = io_diffCommits_info_175_pdest;
        //    mon_tr.io_diffCommits_info_175_rfWen = io_diffCommits_info_175_rfWen;
        //    mon_tr.io_diffCommits_info_175_fpWen = io_diffCommits_info_175_fpWen;
        //    mon_tr.io_diffCommits_info_175_vecWen = io_diffCommits_info_175_vecWen;
        //    mon_tr.io_diffCommits_info_175_v0Wen = io_diffCommits_info_175_v0Wen;
        //    mon_tr.io_diffCommits_info_175_vlWen = io_diffCommits_info_175_vlWen;
        //    mon_tr.io_diffCommits_info_176_ldest = io_diffCommits_info_176_ldest;
        //    mon_tr.io_diffCommits_info_176_pdest = io_diffCommits_info_176_pdest;
        //    mon_tr.io_diffCommits_info_176_rfWen = io_diffCommits_info_176_rfWen;
        //    mon_tr.io_diffCommits_info_176_fpWen = io_diffCommits_info_176_fpWen;
        //    mon_tr.io_diffCommits_info_176_vecWen = io_diffCommits_info_176_vecWen;
        //    mon_tr.io_diffCommits_info_176_v0Wen = io_diffCommits_info_176_v0Wen;
        //    mon_tr.io_diffCommits_info_176_vlWen = io_diffCommits_info_176_vlWen;
        //    mon_tr.io_diffCommits_info_177_ldest = io_diffCommits_info_177_ldest;
        //    mon_tr.io_diffCommits_info_177_pdest = io_diffCommits_info_177_pdest;
        //    mon_tr.io_diffCommits_info_177_rfWen = io_diffCommits_info_177_rfWen;
        //    mon_tr.io_diffCommits_info_177_fpWen = io_diffCommits_info_177_fpWen;
        //    mon_tr.io_diffCommits_info_177_vecWen = io_diffCommits_info_177_vecWen;
        //    mon_tr.io_diffCommits_info_177_v0Wen = io_diffCommits_info_177_v0Wen;
        //    mon_tr.io_diffCommits_info_177_vlWen = io_diffCommits_info_177_vlWen;
        //    mon_tr.io_diffCommits_info_178_ldest = io_diffCommits_info_178_ldest;
        //    mon_tr.io_diffCommits_info_178_pdest = io_diffCommits_info_178_pdest;
        //    mon_tr.io_diffCommits_info_178_rfWen = io_diffCommits_info_178_rfWen;
        //    mon_tr.io_diffCommits_info_178_fpWen = io_diffCommits_info_178_fpWen;
        //    mon_tr.io_diffCommits_info_178_vecWen = io_diffCommits_info_178_vecWen;
        //    mon_tr.io_diffCommits_info_178_v0Wen = io_diffCommits_info_178_v0Wen;
        //    mon_tr.io_diffCommits_info_178_vlWen = io_diffCommits_info_178_vlWen;
        //    mon_tr.io_diffCommits_info_179_ldest = io_diffCommits_info_179_ldest;
        //    mon_tr.io_diffCommits_info_179_pdest = io_diffCommits_info_179_pdest;
        //    mon_tr.io_diffCommits_info_179_rfWen = io_diffCommits_info_179_rfWen;
        //    mon_tr.io_diffCommits_info_179_fpWen = io_diffCommits_info_179_fpWen;
        //    mon_tr.io_diffCommits_info_179_vecWen = io_diffCommits_info_179_vecWen;
        //    mon_tr.io_diffCommits_info_179_v0Wen = io_diffCommits_info_179_v0Wen;
        //    mon_tr.io_diffCommits_info_179_vlWen = io_diffCommits_info_179_vlWen;
        //    mon_tr.io_diffCommits_info_180_ldest = io_diffCommits_info_180_ldest;
        //    mon_tr.io_diffCommits_info_180_pdest = io_diffCommits_info_180_pdest;
        //    mon_tr.io_diffCommits_info_180_rfWen = io_diffCommits_info_180_rfWen;
        //    mon_tr.io_diffCommits_info_180_fpWen = io_diffCommits_info_180_fpWen;
        //    mon_tr.io_diffCommits_info_180_vecWen = io_diffCommits_info_180_vecWen;
        //    mon_tr.io_diffCommits_info_180_v0Wen = io_diffCommits_info_180_v0Wen;
        //    mon_tr.io_diffCommits_info_180_vlWen = io_diffCommits_info_180_vlWen;
        //    mon_tr.io_diffCommits_info_181_ldest = io_diffCommits_info_181_ldest;
        //    mon_tr.io_diffCommits_info_181_pdest = io_diffCommits_info_181_pdest;
        //    mon_tr.io_diffCommits_info_181_rfWen = io_diffCommits_info_181_rfWen;
        //    mon_tr.io_diffCommits_info_181_fpWen = io_diffCommits_info_181_fpWen;
        //    mon_tr.io_diffCommits_info_181_vecWen = io_diffCommits_info_181_vecWen;
        //    mon_tr.io_diffCommits_info_181_v0Wen = io_diffCommits_info_181_v0Wen;
        //    mon_tr.io_diffCommits_info_181_vlWen = io_diffCommits_info_181_vlWen;
        //    mon_tr.io_diffCommits_info_182_ldest = io_diffCommits_info_182_ldest;
        //    mon_tr.io_diffCommits_info_182_pdest = io_diffCommits_info_182_pdest;
        //    mon_tr.io_diffCommits_info_182_rfWen = io_diffCommits_info_182_rfWen;
        //    mon_tr.io_diffCommits_info_182_fpWen = io_diffCommits_info_182_fpWen;
        //    mon_tr.io_diffCommits_info_182_vecWen = io_diffCommits_info_182_vecWen;
        //    mon_tr.io_diffCommits_info_182_v0Wen = io_diffCommits_info_182_v0Wen;
        //    mon_tr.io_diffCommits_info_182_vlWen = io_diffCommits_info_182_vlWen;
        //    mon_tr.io_diffCommits_info_183_ldest = io_diffCommits_info_183_ldest;
        //    mon_tr.io_diffCommits_info_183_pdest = io_diffCommits_info_183_pdest;
        //    mon_tr.io_diffCommits_info_183_rfWen = io_diffCommits_info_183_rfWen;
        //    mon_tr.io_diffCommits_info_183_fpWen = io_diffCommits_info_183_fpWen;
        //    mon_tr.io_diffCommits_info_183_vecWen = io_diffCommits_info_183_vecWen;
        //    mon_tr.io_diffCommits_info_183_v0Wen = io_diffCommits_info_183_v0Wen;
        //    mon_tr.io_diffCommits_info_183_vlWen = io_diffCommits_info_183_vlWen;
        //    mon_tr.io_diffCommits_info_184_ldest = io_diffCommits_info_184_ldest;
        //    mon_tr.io_diffCommits_info_184_pdest = io_diffCommits_info_184_pdest;
        //    mon_tr.io_diffCommits_info_184_rfWen = io_diffCommits_info_184_rfWen;
        //    mon_tr.io_diffCommits_info_184_fpWen = io_diffCommits_info_184_fpWen;
        //    mon_tr.io_diffCommits_info_184_vecWen = io_diffCommits_info_184_vecWen;
        //    mon_tr.io_diffCommits_info_184_v0Wen = io_diffCommits_info_184_v0Wen;
        //    mon_tr.io_diffCommits_info_184_vlWen = io_diffCommits_info_184_vlWen;
        //    mon_tr.io_diffCommits_info_185_ldest = io_diffCommits_info_185_ldest;
        //    mon_tr.io_diffCommits_info_185_pdest = io_diffCommits_info_185_pdest;
        //    mon_tr.io_diffCommits_info_185_rfWen = io_diffCommits_info_185_rfWen;
        //    mon_tr.io_diffCommits_info_185_fpWen = io_diffCommits_info_185_fpWen;
        //    mon_tr.io_diffCommits_info_185_vecWen = io_diffCommits_info_185_vecWen;
        //    mon_tr.io_diffCommits_info_185_v0Wen = io_diffCommits_info_185_v0Wen;
        //    mon_tr.io_diffCommits_info_185_vlWen = io_diffCommits_info_185_vlWen;
        //    mon_tr.io_diffCommits_info_186_ldest = io_diffCommits_info_186_ldest;
        //    mon_tr.io_diffCommits_info_186_pdest = io_diffCommits_info_186_pdest;
        //    mon_tr.io_diffCommits_info_186_rfWen = io_diffCommits_info_186_rfWen;
        //    mon_tr.io_diffCommits_info_186_fpWen = io_diffCommits_info_186_fpWen;
        //    mon_tr.io_diffCommits_info_186_vecWen = io_diffCommits_info_186_vecWen;
        //    mon_tr.io_diffCommits_info_186_v0Wen = io_diffCommits_info_186_v0Wen;
        //    mon_tr.io_diffCommits_info_186_vlWen = io_diffCommits_info_186_vlWen;
        //    mon_tr.io_diffCommits_info_187_ldest = io_diffCommits_info_187_ldest;
        //    mon_tr.io_diffCommits_info_187_pdest = io_diffCommits_info_187_pdest;
        //    mon_tr.io_diffCommits_info_187_rfWen = io_diffCommits_info_187_rfWen;
        //    mon_tr.io_diffCommits_info_187_fpWen = io_diffCommits_info_187_fpWen;
        //    mon_tr.io_diffCommits_info_187_vecWen = io_diffCommits_info_187_vecWen;
        //    mon_tr.io_diffCommits_info_187_v0Wen = io_diffCommits_info_187_v0Wen;
        //    mon_tr.io_diffCommits_info_187_vlWen = io_diffCommits_info_187_vlWen;
        //    mon_tr.io_diffCommits_info_188_ldest = io_diffCommits_info_188_ldest;
        //    mon_tr.io_diffCommits_info_188_pdest = io_diffCommits_info_188_pdest;
        //    mon_tr.io_diffCommits_info_188_rfWen = io_diffCommits_info_188_rfWen;
        //    mon_tr.io_diffCommits_info_188_fpWen = io_diffCommits_info_188_fpWen;
        //    mon_tr.io_diffCommits_info_188_vecWen = io_diffCommits_info_188_vecWen;
        //    mon_tr.io_diffCommits_info_188_v0Wen = io_diffCommits_info_188_v0Wen;
        //    mon_tr.io_diffCommits_info_188_vlWen = io_diffCommits_info_188_vlWen;
        //    mon_tr.io_diffCommits_info_189_ldest = io_diffCommits_info_189_ldest;
        //    mon_tr.io_diffCommits_info_189_pdest = io_diffCommits_info_189_pdest;
        //    mon_tr.io_diffCommits_info_189_rfWen = io_diffCommits_info_189_rfWen;
        //    mon_tr.io_diffCommits_info_189_fpWen = io_diffCommits_info_189_fpWen;
        //    mon_tr.io_diffCommits_info_189_vecWen = io_diffCommits_info_189_vecWen;
        //    mon_tr.io_diffCommits_info_189_v0Wen = io_diffCommits_info_189_v0Wen;
        //    mon_tr.io_diffCommits_info_189_vlWen = io_diffCommits_info_189_vlWen;
        //    mon_tr.io_diffCommits_info_190_ldest = io_diffCommits_info_190_ldest;
        //    mon_tr.io_diffCommits_info_190_pdest = io_diffCommits_info_190_pdest;
        //    mon_tr.io_diffCommits_info_190_rfWen = io_diffCommits_info_190_rfWen;
        //    mon_tr.io_diffCommits_info_190_fpWen = io_diffCommits_info_190_fpWen;
        //    mon_tr.io_diffCommits_info_190_vecWen = io_diffCommits_info_190_vecWen;
        //    mon_tr.io_diffCommits_info_190_v0Wen = io_diffCommits_info_190_v0Wen;
        //    mon_tr.io_diffCommits_info_190_vlWen = io_diffCommits_info_190_vlWen;
        //    mon_tr.io_diffCommits_info_191_ldest = io_diffCommits_info_191_ldest;
        //    mon_tr.io_diffCommits_info_191_pdest = io_diffCommits_info_191_pdest;
        //    mon_tr.io_diffCommits_info_191_rfWen = io_diffCommits_info_191_rfWen;
        //    mon_tr.io_diffCommits_info_191_fpWen = io_diffCommits_info_191_fpWen;
        //    mon_tr.io_diffCommits_info_191_vecWen = io_diffCommits_info_191_vecWen;
        //    mon_tr.io_diffCommits_info_191_v0Wen = io_diffCommits_info_191_v0Wen;
        //    mon_tr.io_diffCommits_info_191_vlWen = io_diffCommits_info_191_vlWen;
        //    mon_tr.io_diffCommits_info_192_ldest = io_diffCommits_info_192_ldest;
        //    mon_tr.io_diffCommits_info_192_pdest = io_diffCommits_info_192_pdest;
        //    mon_tr.io_diffCommits_info_192_rfWen = io_diffCommits_info_192_rfWen;
        //    mon_tr.io_diffCommits_info_192_fpWen = io_diffCommits_info_192_fpWen;
        //    mon_tr.io_diffCommits_info_192_vecWen = io_diffCommits_info_192_vecWen;
        //    mon_tr.io_diffCommits_info_192_v0Wen = io_diffCommits_info_192_v0Wen;
        //    mon_tr.io_diffCommits_info_192_vlWen = io_diffCommits_info_192_vlWen;
        //    mon_tr.io_diffCommits_info_193_ldest = io_diffCommits_info_193_ldest;
        //    mon_tr.io_diffCommits_info_193_pdest = io_diffCommits_info_193_pdest;
        //    mon_tr.io_diffCommits_info_193_rfWen = io_diffCommits_info_193_rfWen;
        //    mon_tr.io_diffCommits_info_193_fpWen = io_diffCommits_info_193_fpWen;
        //    mon_tr.io_diffCommits_info_193_vecWen = io_diffCommits_info_193_vecWen;
        //    mon_tr.io_diffCommits_info_193_v0Wen = io_diffCommits_info_193_v0Wen;
        //    mon_tr.io_diffCommits_info_193_vlWen = io_diffCommits_info_193_vlWen;
        //    mon_tr.io_diffCommits_info_194_ldest = io_diffCommits_info_194_ldest;
        //    mon_tr.io_diffCommits_info_194_pdest = io_diffCommits_info_194_pdest;
        //    mon_tr.io_diffCommits_info_194_rfWen = io_diffCommits_info_194_rfWen;
        //    mon_tr.io_diffCommits_info_194_fpWen = io_diffCommits_info_194_fpWen;
        //    mon_tr.io_diffCommits_info_194_vecWen = io_diffCommits_info_194_vecWen;
        //    mon_tr.io_diffCommits_info_194_v0Wen = io_diffCommits_info_194_v0Wen;
        //    mon_tr.io_diffCommits_info_194_vlWen = io_diffCommits_info_194_vlWen;
        //    mon_tr.io_diffCommits_info_195_ldest = io_diffCommits_info_195_ldest;
        //    mon_tr.io_diffCommits_info_195_pdest = io_diffCommits_info_195_pdest;
        //    mon_tr.io_diffCommits_info_195_rfWen = io_diffCommits_info_195_rfWen;
        //    mon_tr.io_diffCommits_info_195_fpWen = io_diffCommits_info_195_fpWen;
        //    mon_tr.io_diffCommits_info_195_vecWen = io_diffCommits_info_195_vecWen;
        //    mon_tr.io_diffCommits_info_195_v0Wen = io_diffCommits_info_195_v0Wen;
        //    mon_tr.io_diffCommits_info_195_vlWen = io_diffCommits_info_195_vlWen;
        //    mon_tr.io_diffCommits_info_196_ldest = io_diffCommits_info_196_ldest;
        //    mon_tr.io_diffCommits_info_196_pdest = io_diffCommits_info_196_pdest;
        //    mon_tr.io_diffCommits_info_196_rfWen = io_diffCommits_info_196_rfWen;
        //    mon_tr.io_diffCommits_info_196_fpWen = io_diffCommits_info_196_fpWen;
        //    mon_tr.io_diffCommits_info_196_vecWen = io_diffCommits_info_196_vecWen;
        //    mon_tr.io_diffCommits_info_196_v0Wen = io_diffCommits_info_196_v0Wen;
        //    mon_tr.io_diffCommits_info_196_vlWen = io_diffCommits_info_196_vlWen;
        //    mon_tr.io_diffCommits_info_197_ldest = io_diffCommits_info_197_ldest;
        //    mon_tr.io_diffCommits_info_197_pdest = io_diffCommits_info_197_pdest;
        //    mon_tr.io_diffCommits_info_197_rfWen = io_diffCommits_info_197_rfWen;
        //    mon_tr.io_diffCommits_info_197_fpWen = io_diffCommits_info_197_fpWen;
        //    mon_tr.io_diffCommits_info_197_vecWen = io_diffCommits_info_197_vecWen;
        //    mon_tr.io_diffCommits_info_197_v0Wen = io_diffCommits_info_197_v0Wen;
        //    mon_tr.io_diffCommits_info_197_vlWen = io_diffCommits_info_197_vlWen;
        //    mon_tr.io_diffCommits_info_198_ldest = io_diffCommits_info_198_ldest;
        //    mon_tr.io_diffCommits_info_198_pdest = io_diffCommits_info_198_pdest;
        //    mon_tr.io_diffCommits_info_198_rfWen = io_diffCommits_info_198_rfWen;
        //    mon_tr.io_diffCommits_info_198_fpWen = io_diffCommits_info_198_fpWen;
        //    mon_tr.io_diffCommits_info_198_vecWen = io_diffCommits_info_198_vecWen;
        //    mon_tr.io_diffCommits_info_198_v0Wen = io_diffCommits_info_198_v0Wen;
        //    mon_tr.io_diffCommits_info_198_vlWen = io_diffCommits_info_198_vlWen;
        //    mon_tr.io_diffCommits_info_199_ldest = io_diffCommits_info_199_ldest;
        //    mon_tr.io_diffCommits_info_199_pdest = io_diffCommits_info_199_pdest;
        //    mon_tr.io_diffCommits_info_199_rfWen = io_diffCommits_info_199_rfWen;
        //    mon_tr.io_diffCommits_info_199_fpWen = io_diffCommits_info_199_fpWen;
        //    mon_tr.io_diffCommits_info_199_vecWen = io_diffCommits_info_199_vecWen;
        //    mon_tr.io_diffCommits_info_199_v0Wen = io_diffCommits_info_199_v0Wen;
        //    mon_tr.io_diffCommits_info_199_vlWen = io_diffCommits_info_199_vlWen;
        //    mon_tr.io_diffCommits_info_200_ldest = io_diffCommits_info_200_ldest;
        //    mon_tr.io_diffCommits_info_200_pdest = io_diffCommits_info_200_pdest;
        //    mon_tr.io_diffCommits_info_200_rfWen = io_diffCommits_info_200_rfWen;
        //    mon_tr.io_diffCommits_info_200_fpWen = io_diffCommits_info_200_fpWen;
        //    mon_tr.io_diffCommits_info_200_vecWen = io_diffCommits_info_200_vecWen;
        //    mon_tr.io_diffCommits_info_200_v0Wen = io_diffCommits_info_200_v0Wen;
        //    mon_tr.io_diffCommits_info_200_vlWen = io_diffCommits_info_200_vlWen;
        //    mon_tr.io_diffCommits_info_201_ldest = io_diffCommits_info_201_ldest;
        //    mon_tr.io_diffCommits_info_201_pdest = io_diffCommits_info_201_pdest;
        //    mon_tr.io_diffCommits_info_201_rfWen = io_diffCommits_info_201_rfWen;
        //    mon_tr.io_diffCommits_info_201_fpWen = io_diffCommits_info_201_fpWen;
        //    mon_tr.io_diffCommits_info_201_vecWen = io_diffCommits_info_201_vecWen;
        //    mon_tr.io_diffCommits_info_201_v0Wen = io_diffCommits_info_201_v0Wen;
        //    mon_tr.io_diffCommits_info_201_vlWen = io_diffCommits_info_201_vlWen;
        //    mon_tr.io_diffCommits_info_202_ldest = io_diffCommits_info_202_ldest;
        //    mon_tr.io_diffCommits_info_202_pdest = io_diffCommits_info_202_pdest;
        //    mon_tr.io_diffCommits_info_202_rfWen = io_diffCommits_info_202_rfWen;
        //    mon_tr.io_diffCommits_info_202_fpWen = io_diffCommits_info_202_fpWen;
        //    mon_tr.io_diffCommits_info_202_vecWen = io_diffCommits_info_202_vecWen;
        //    mon_tr.io_diffCommits_info_202_v0Wen = io_diffCommits_info_202_v0Wen;
        //    mon_tr.io_diffCommits_info_202_vlWen = io_diffCommits_info_202_vlWen;
        //    mon_tr.io_diffCommits_info_203_ldest = io_diffCommits_info_203_ldest;
        //    mon_tr.io_diffCommits_info_203_pdest = io_diffCommits_info_203_pdest;
        //    mon_tr.io_diffCommits_info_203_rfWen = io_diffCommits_info_203_rfWen;
        //    mon_tr.io_diffCommits_info_203_fpWen = io_diffCommits_info_203_fpWen;
        //    mon_tr.io_diffCommits_info_203_vecWen = io_diffCommits_info_203_vecWen;
        //    mon_tr.io_diffCommits_info_203_v0Wen = io_diffCommits_info_203_v0Wen;
        //    mon_tr.io_diffCommits_info_203_vlWen = io_diffCommits_info_203_vlWen;
        //    mon_tr.io_diffCommits_info_204_ldest = io_diffCommits_info_204_ldest;
        //    mon_tr.io_diffCommits_info_204_pdest = io_diffCommits_info_204_pdest;
        //    mon_tr.io_diffCommits_info_204_rfWen = io_diffCommits_info_204_rfWen;
        //    mon_tr.io_diffCommits_info_204_fpWen = io_diffCommits_info_204_fpWen;
        //    mon_tr.io_diffCommits_info_204_vecWen = io_diffCommits_info_204_vecWen;
        //    mon_tr.io_diffCommits_info_204_v0Wen = io_diffCommits_info_204_v0Wen;
        //    mon_tr.io_diffCommits_info_204_vlWen = io_diffCommits_info_204_vlWen;
        //    mon_tr.io_diffCommits_info_205_ldest = io_diffCommits_info_205_ldest;
        //    mon_tr.io_diffCommits_info_205_pdest = io_diffCommits_info_205_pdest;
        //    mon_tr.io_diffCommits_info_205_rfWen = io_diffCommits_info_205_rfWen;
        //    mon_tr.io_diffCommits_info_205_fpWen = io_diffCommits_info_205_fpWen;
        //    mon_tr.io_diffCommits_info_205_vecWen = io_diffCommits_info_205_vecWen;
        //    mon_tr.io_diffCommits_info_205_v0Wen = io_diffCommits_info_205_v0Wen;
        //    mon_tr.io_diffCommits_info_205_vlWen = io_diffCommits_info_205_vlWen;
        //    mon_tr.io_diffCommits_info_206_ldest = io_diffCommits_info_206_ldest;
        //    mon_tr.io_diffCommits_info_206_pdest = io_diffCommits_info_206_pdest;
        //    mon_tr.io_diffCommits_info_206_rfWen = io_diffCommits_info_206_rfWen;
        //    mon_tr.io_diffCommits_info_206_fpWen = io_diffCommits_info_206_fpWen;
        //    mon_tr.io_diffCommits_info_206_vecWen = io_diffCommits_info_206_vecWen;
        //    mon_tr.io_diffCommits_info_206_v0Wen = io_diffCommits_info_206_v0Wen;
        //    mon_tr.io_diffCommits_info_206_vlWen = io_diffCommits_info_206_vlWen;
        //    mon_tr.io_diffCommits_info_207_ldest = io_diffCommits_info_207_ldest;
        //    mon_tr.io_diffCommits_info_207_pdest = io_diffCommits_info_207_pdest;
        //    mon_tr.io_diffCommits_info_207_rfWen = io_diffCommits_info_207_rfWen;
        //    mon_tr.io_diffCommits_info_207_fpWen = io_diffCommits_info_207_fpWen;
        //    mon_tr.io_diffCommits_info_207_vecWen = io_diffCommits_info_207_vecWen;
        //    mon_tr.io_diffCommits_info_207_v0Wen = io_diffCommits_info_207_v0Wen;
        //    mon_tr.io_diffCommits_info_207_vlWen = io_diffCommits_info_207_vlWen;
        //    mon_tr.io_diffCommits_info_208_ldest = io_diffCommits_info_208_ldest;
        //    mon_tr.io_diffCommits_info_208_pdest = io_diffCommits_info_208_pdest;
        //    mon_tr.io_diffCommits_info_208_rfWen = io_diffCommits_info_208_rfWen;
        //    mon_tr.io_diffCommits_info_208_fpWen = io_diffCommits_info_208_fpWen;
        //    mon_tr.io_diffCommits_info_208_vecWen = io_diffCommits_info_208_vecWen;
        //    mon_tr.io_diffCommits_info_208_v0Wen = io_diffCommits_info_208_v0Wen;
        //    mon_tr.io_diffCommits_info_208_vlWen = io_diffCommits_info_208_vlWen;
        //    mon_tr.io_diffCommits_info_209_ldest = io_diffCommits_info_209_ldest;
        //    mon_tr.io_diffCommits_info_209_pdest = io_diffCommits_info_209_pdest;
        //    mon_tr.io_diffCommits_info_209_rfWen = io_diffCommits_info_209_rfWen;
        //    mon_tr.io_diffCommits_info_209_fpWen = io_diffCommits_info_209_fpWen;
        //    mon_tr.io_diffCommits_info_209_vecWen = io_diffCommits_info_209_vecWen;
        //    mon_tr.io_diffCommits_info_209_v0Wen = io_diffCommits_info_209_v0Wen;
        //    mon_tr.io_diffCommits_info_209_vlWen = io_diffCommits_info_209_vlWen;
        //    mon_tr.io_diffCommits_info_210_ldest = io_diffCommits_info_210_ldest;
        //    mon_tr.io_diffCommits_info_210_pdest = io_diffCommits_info_210_pdest;
        //    mon_tr.io_diffCommits_info_210_rfWen = io_diffCommits_info_210_rfWen;
        //    mon_tr.io_diffCommits_info_210_fpWen = io_diffCommits_info_210_fpWen;
        //    mon_tr.io_diffCommits_info_210_vecWen = io_diffCommits_info_210_vecWen;
        //    mon_tr.io_diffCommits_info_210_v0Wen = io_diffCommits_info_210_v0Wen;
        //    mon_tr.io_diffCommits_info_210_vlWen = io_diffCommits_info_210_vlWen;
        //    mon_tr.io_diffCommits_info_211_ldest = io_diffCommits_info_211_ldest;
        //    mon_tr.io_diffCommits_info_211_pdest = io_diffCommits_info_211_pdest;
        //    mon_tr.io_diffCommits_info_211_rfWen = io_diffCommits_info_211_rfWen;
        //    mon_tr.io_diffCommits_info_211_fpWen = io_diffCommits_info_211_fpWen;
        //    mon_tr.io_diffCommits_info_211_vecWen = io_diffCommits_info_211_vecWen;
        //    mon_tr.io_diffCommits_info_211_v0Wen = io_diffCommits_info_211_v0Wen;
        //    mon_tr.io_diffCommits_info_211_vlWen = io_diffCommits_info_211_vlWen;
        //    mon_tr.io_diffCommits_info_212_ldest = io_diffCommits_info_212_ldest;
        //    mon_tr.io_diffCommits_info_212_pdest = io_diffCommits_info_212_pdest;
        //    mon_tr.io_diffCommits_info_212_rfWen = io_diffCommits_info_212_rfWen;
        //    mon_tr.io_diffCommits_info_212_fpWen = io_diffCommits_info_212_fpWen;
        //    mon_tr.io_diffCommits_info_212_vecWen = io_diffCommits_info_212_vecWen;
        //    mon_tr.io_diffCommits_info_212_v0Wen = io_diffCommits_info_212_v0Wen;
        //    mon_tr.io_diffCommits_info_212_vlWen = io_diffCommits_info_212_vlWen;
        //    mon_tr.io_diffCommits_info_213_ldest = io_diffCommits_info_213_ldest;
        //    mon_tr.io_diffCommits_info_213_pdest = io_diffCommits_info_213_pdest;
        //    mon_tr.io_diffCommits_info_213_rfWen = io_diffCommits_info_213_rfWen;
        //    mon_tr.io_diffCommits_info_213_fpWen = io_diffCommits_info_213_fpWen;
        //    mon_tr.io_diffCommits_info_213_vecWen = io_diffCommits_info_213_vecWen;
        //    mon_tr.io_diffCommits_info_213_v0Wen = io_diffCommits_info_213_v0Wen;
        //    mon_tr.io_diffCommits_info_213_vlWen = io_diffCommits_info_213_vlWen;
        //    mon_tr.io_diffCommits_info_214_ldest = io_diffCommits_info_214_ldest;
        //    mon_tr.io_diffCommits_info_214_pdest = io_diffCommits_info_214_pdest;
        //    mon_tr.io_diffCommits_info_214_rfWen = io_diffCommits_info_214_rfWen;
        //    mon_tr.io_diffCommits_info_214_fpWen = io_diffCommits_info_214_fpWen;
        //    mon_tr.io_diffCommits_info_214_vecWen = io_diffCommits_info_214_vecWen;
        //    mon_tr.io_diffCommits_info_214_v0Wen = io_diffCommits_info_214_v0Wen;
        //    mon_tr.io_diffCommits_info_214_vlWen = io_diffCommits_info_214_vlWen;
        //    mon_tr.io_diffCommits_info_215_ldest = io_diffCommits_info_215_ldest;
        //    mon_tr.io_diffCommits_info_215_pdest = io_diffCommits_info_215_pdest;
        //    mon_tr.io_diffCommits_info_215_rfWen = io_diffCommits_info_215_rfWen;
        //    mon_tr.io_diffCommits_info_215_fpWen = io_diffCommits_info_215_fpWen;
        //    mon_tr.io_diffCommits_info_215_vecWen = io_diffCommits_info_215_vecWen;
        //    mon_tr.io_diffCommits_info_215_v0Wen = io_diffCommits_info_215_v0Wen;
        //    mon_tr.io_diffCommits_info_215_vlWen = io_diffCommits_info_215_vlWen;
        //    mon_tr.io_diffCommits_info_216_ldest = io_diffCommits_info_216_ldest;
        //    mon_tr.io_diffCommits_info_216_pdest = io_diffCommits_info_216_pdest;
        //    mon_tr.io_diffCommits_info_216_rfWen = io_diffCommits_info_216_rfWen;
        //    mon_tr.io_diffCommits_info_216_fpWen = io_diffCommits_info_216_fpWen;
        //    mon_tr.io_diffCommits_info_216_vecWen = io_diffCommits_info_216_vecWen;
        //    mon_tr.io_diffCommits_info_216_v0Wen = io_diffCommits_info_216_v0Wen;
        //    mon_tr.io_diffCommits_info_216_vlWen = io_diffCommits_info_216_vlWen;
        //    mon_tr.io_diffCommits_info_217_ldest = io_diffCommits_info_217_ldest;
        //    mon_tr.io_diffCommits_info_217_pdest = io_diffCommits_info_217_pdest;
        //    mon_tr.io_diffCommits_info_217_rfWen = io_diffCommits_info_217_rfWen;
        //    mon_tr.io_diffCommits_info_217_fpWen = io_diffCommits_info_217_fpWen;
        //    mon_tr.io_diffCommits_info_217_vecWen = io_diffCommits_info_217_vecWen;
        //    mon_tr.io_diffCommits_info_217_v0Wen = io_diffCommits_info_217_v0Wen;
        //    mon_tr.io_diffCommits_info_217_vlWen = io_diffCommits_info_217_vlWen;
        //    mon_tr.io_diffCommits_info_218_ldest = io_diffCommits_info_218_ldest;
        //    mon_tr.io_diffCommits_info_218_pdest = io_diffCommits_info_218_pdest;
        //    mon_tr.io_diffCommits_info_218_rfWen = io_diffCommits_info_218_rfWen;
        //    mon_tr.io_diffCommits_info_218_fpWen = io_diffCommits_info_218_fpWen;
        //    mon_tr.io_diffCommits_info_218_vecWen = io_diffCommits_info_218_vecWen;
        //    mon_tr.io_diffCommits_info_218_v0Wen = io_diffCommits_info_218_v0Wen;
        //    mon_tr.io_diffCommits_info_218_vlWen = io_diffCommits_info_218_vlWen;
        //    mon_tr.io_diffCommits_info_219_ldest = io_diffCommits_info_219_ldest;
        //    mon_tr.io_diffCommits_info_219_pdest = io_diffCommits_info_219_pdest;
        //    mon_tr.io_diffCommits_info_219_rfWen = io_diffCommits_info_219_rfWen;
        //    mon_tr.io_diffCommits_info_219_fpWen = io_diffCommits_info_219_fpWen;
        //    mon_tr.io_diffCommits_info_219_vecWen = io_diffCommits_info_219_vecWen;
        //    mon_tr.io_diffCommits_info_219_v0Wen = io_diffCommits_info_219_v0Wen;
        //    mon_tr.io_diffCommits_info_219_vlWen = io_diffCommits_info_219_vlWen;
        //    mon_tr.io_diffCommits_info_220_ldest = io_diffCommits_info_220_ldest;
        //    mon_tr.io_diffCommits_info_220_pdest = io_diffCommits_info_220_pdest;
        //    mon_tr.io_diffCommits_info_220_rfWen = io_diffCommits_info_220_rfWen;
        //    mon_tr.io_diffCommits_info_220_fpWen = io_diffCommits_info_220_fpWen;
        //    mon_tr.io_diffCommits_info_220_vecWen = io_diffCommits_info_220_vecWen;
        //    mon_tr.io_diffCommits_info_220_v0Wen = io_diffCommits_info_220_v0Wen;
        //    mon_tr.io_diffCommits_info_220_vlWen = io_diffCommits_info_220_vlWen;
        //    mon_tr.io_diffCommits_info_221_ldest = io_diffCommits_info_221_ldest;
        //    mon_tr.io_diffCommits_info_221_pdest = io_diffCommits_info_221_pdest;
        //    mon_tr.io_diffCommits_info_221_rfWen = io_diffCommits_info_221_rfWen;
        //    mon_tr.io_diffCommits_info_221_fpWen = io_diffCommits_info_221_fpWen;
        //    mon_tr.io_diffCommits_info_221_vecWen = io_diffCommits_info_221_vecWen;
        //    mon_tr.io_diffCommits_info_221_v0Wen = io_diffCommits_info_221_v0Wen;
        //    mon_tr.io_diffCommits_info_221_vlWen = io_diffCommits_info_221_vlWen;
        //    mon_tr.io_diffCommits_info_222_ldest = io_diffCommits_info_222_ldest;
        //    mon_tr.io_diffCommits_info_222_pdest = io_diffCommits_info_222_pdest;
        //    mon_tr.io_diffCommits_info_222_rfWen = io_diffCommits_info_222_rfWen;
        //    mon_tr.io_diffCommits_info_222_fpWen = io_diffCommits_info_222_fpWen;
        //    mon_tr.io_diffCommits_info_222_vecWen = io_diffCommits_info_222_vecWen;
        //    mon_tr.io_diffCommits_info_222_v0Wen = io_diffCommits_info_222_v0Wen;
        //    mon_tr.io_diffCommits_info_222_vlWen = io_diffCommits_info_222_vlWen;
        //    mon_tr.io_diffCommits_info_223_ldest = io_diffCommits_info_223_ldest;
        //    mon_tr.io_diffCommits_info_223_pdest = io_diffCommits_info_223_pdest;
        //    mon_tr.io_diffCommits_info_223_rfWen = io_diffCommits_info_223_rfWen;
        //    mon_tr.io_diffCommits_info_223_fpWen = io_diffCommits_info_223_fpWen;
        //    mon_tr.io_diffCommits_info_223_vecWen = io_diffCommits_info_223_vecWen;
        //    mon_tr.io_diffCommits_info_223_v0Wen = io_diffCommits_info_223_v0Wen;
        //    mon_tr.io_diffCommits_info_223_vlWen = io_diffCommits_info_223_vlWen;
        //    mon_tr.io_diffCommits_info_224_ldest = io_diffCommits_info_224_ldest;
        //    mon_tr.io_diffCommits_info_224_pdest = io_diffCommits_info_224_pdest;
        //    mon_tr.io_diffCommits_info_224_rfWen = io_diffCommits_info_224_rfWen;
        //    mon_tr.io_diffCommits_info_224_fpWen = io_diffCommits_info_224_fpWen;
        //    mon_tr.io_diffCommits_info_224_vecWen = io_diffCommits_info_224_vecWen;
        //    mon_tr.io_diffCommits_info_224_v0Wen = io_diffCommits_info_224_v0Wen;
        //    mon_tr.io_diffCommits_info_224_vlWen = io_diffCommits_info_224_vlWen;
        //    mon_tr.io_diffCommits_info_225_ldest = io_diffCommits_info_225_ldest;
        //    mon_tr.io_diffCommits_info_225_pdest = io_diffCommits_info_225_pdest;
        //    mon_tr.io_diffCommits_info_225_rfWen = io_diffCommits_info_225_rfWen;
        //    mon_tr.io_diffCommits_info_225_fpWen = io_diffCommits_info_225_fpWen;
        //    mon_tr.io_diffCommits_info_225_vecWen = io_diffCommits_info_225_vecWen;
        //    mon_tr.io_diffCommits_info_225_v0Wen = io_diffCommits_info_225_v0Wen;
        //    mon_tr.io_diffCommits_info_225_vlWen = io_diffCommits_info_225_vlWen;
        //    mon_tr.io_diffCommits_info_226_ldest = io_diffCommits_info_226_ldest;
        //    mon_tr.io_diffCommits_info_226_pdest = io_diffCommits_info_226_pdest;
        //    mon_tr.io_diffCommits_info_226_rfWen = io_diffCommits_info_226_rfWen;
        //    mon_tr.io_diffCommits_info_226_fpWen = io_diffCommits_info_226_fpWen;
        //    mon_tr.io_diffCommits_info_226_vecWen = io_diffCommits_info_226_vecWen;
        //    mon_tr.io_diffCommits_info_226_v0Wen = io_diffCommits_info_226_v0Wen;
        //    mon_tr.io_diffCommits_info_226_vlWen = io_diffCommits_info_226_vlWen;
        //    mon_tr.io_diffCommits_info_227_ldest = io_diffCommits_info_227_ldest;
        //    mon_tr.io_diffCommits_info_227_pdest = io_diffCommits_info_227_pdest;
        //    mon_tr.io_diffCommits_info_227_rfWen = io_diffCommits_info_227_rfWen;
        //    mon_tr.io_diffCommits_info_227_fpWen = io_diffCommits_info_227_fpWen;
        //    mon_tr.io_diffCommits_info_227_vecWen = io_diffCommits_info_227_vecWen;
        //    mon_tr.io_diffCommits_info_227_v0Wen = io_diffCommits_info_227_v0Wen;
        //    mon_tr.io_diffCommits_info_227_vlWen = io_diffCommits_info_227_vlWen;
        //    mon_tr.io_diffCommits_info_228_ldest = io_diffCommits_info_228_ldest;
        //    mon_tr.io_diffCommits_info_228_pdest = io_diffCommits_info_228_pdest;
        //    mon_tr.io_diffCommits_info_228_rfWen = io_diffCommits_info_228_rfWen;
        //    mon_tr.io_diffCommits_info_228_fpWen = io_diffCommits_info_228_fpWen;
        //    mon_tr.io_diffCommits_info_228_vecWen = io_diffCommits_info_228_vecWen;
        //    mon_tr.io_diffCommits_info_228_v0Wen = io_diffCommits_info_228_v0Wen;
        //    mon_tr.io_diffCommits_info_228_vlWen = io_diffCommits_info_228_vlWen;
        //    mon_tr.io_diffCommits_info_229_ldest = io_diffCommits_info_229_ldest;
        //    mon_tr.io_diffCommits_info_229_pdest = io_diffCommits_info_229_pdest;
        //    mon_tr.io_diffCommits_info_229_rfWen = io_diffCommits_info_229_rfWen;
        //    mon_tr.io_diffCommits_info_229_fpWen = io_diffCommits_info_229_fpWen;
        //    mon_tr.io_diffCommits_info_229_vecWen = io_diffCommits_info_229_vecWen;
        //    mon_tr.io_diffCommits_info_229_v0Wen = io_diffCommits_info_229_v0Wen;
        //    mon_tr.io_diffCommits_info_229_vlWen = io_diffCommits_info_229_vlWen;
        //    mon_tr.io_diffCommits_info_230_ldest = io_diffCommits_info_230_ldest;
        //    mon_tr.io_diffCommits_info_230_pdest = io_diffCommits_info_230_pdest;
        //    mon_tr.io_diffCommits_info_230_rfWen = io_diffCommits_info_230_rfWen;
        //    mon_tr.io_diffCommits_info_230_fpWen = io_diffCommits_info_230_fpWen;
        //    mon_tr.io_diffCommits_info_230_vecWen = io_diffCommits_info_230_vecWen;
        //    mon_tr.io_diffCommits_info_230_v0Wen = io_diffCommits_info_230_v0Wen;
        //    mon_tr.io_diffCommits_info_230_vlWen = io_diffCommits_info_230_vlWen;
        //    mon_tr.io_diffCommits_info_231_ldest = io_diffCommits_info_231_ldest;
        //    mon_tr.io_diffCommits_info_231_pdest = io_diffCommits_info_231_pdest;
        //    mon_tr.io_diffCommits_info_231_rfWen = io_diffCommits_info_231_rfWen;
        //    mon_tr.io_diffCommits_info_231_fpWen = io_diffCommits_info_231_fpWen;
        //    mon_tr.io_diffCommits_info_231_vecWen = io_diffCommits_info_231_vecWen;
        //    mon_tr.io_diffCommits_info_231_v0Wen = io_diffCommits_info_231_v0Wen;
        //    mon_tr.io_diffCommits_info_231_vlWen = io_diffCommits_info_231_vlWen;
        //    mon_tr.io_diffCommits_info_232_ldest = io_diffCommits_info_232_ldest;
        //    mon_tr.io_diffCommits_info_232_pdest = io_diffCommits_info_232_pdest;
        //    mon_tr.io_diffCommits_info_232_rfWen = io_diffCommits_info_232_rfWen;
        //    mon_tr.io_diffCommits_info_232_fpWen = io_diffCommits_info_232_fpWen;
        //    mon_tr.io_diffCommits_info_232_vecWen = io_diffCommits_info_232_vecWen;
        //    mon_tr.io_diffCommits_info_232_v0Wen = io_diffCommits_info_232_v0Wen;
        //    mon_tr.io_diffCommits_info_232_vlWen = io_diffCommits_info_232_vlWen;
        //    mon_tr.io_diffCommits_info_233_ldest = io_diffCommits_info_233_ldest;
        //    mon_tr.io_diffCommits_info_233_pdest = io_diffCommits_info_233_pdest;
        //    mon_tr.io_diffCommits_info_233_rfWen = io_diffCommits_info_233_rfWen;
        //    mon_tr.io_diffCommits_info_233_fpWen = io_diffCommits_info_233_fpWen;
        //    mon_tr.io_diffCommits_info_233_vecWen = io_diffCommits_info_233_vecWen;
        //    mon_tr.io_diffCommits_info_233_v0Wen = io_diffCommits_info_233_v0Wen;
        //    mon_tr.io_diffCommits_info_233_vlWen = io_diffCommits_info_233_vlWen;
        //    mon_tr.io_diffCommits_info_234_ldest = io_diffCommits_info_234_ldest;
        //    mon_tr.io_diffCommits_info_234_pdest = io_diffCommits_info_234_pdest;
        //    mon_tr.io_diffCommits_info_234_rfWen = io_diffCommits_info_234_rfWen;
        //    mon_tr.io_diffCommits_info_234_fpWen = io_diffCommits_info_234_fpWen;
        //    mon_tr.io_diffCommits_info_234_vecWen = io_diffCommits_info_234_vecWen;
        //    mon_tr.io_diffCommits_info_234_v0Wen = io_diffCommits_info_234_v0Wen;
        //    mon_tr.io_diffCommits_info_234_vlWen = io_diffCommits_info_234_vlWen;
        //    mon_tr.io_diffCommits_info_235_ldest = io_diffCommits_info_235_ldest;
        //    mon_tr.io_diffCommits_info_235_pdest = io_diffCommits_info_235_pdest;
        //    mon_tr.io_diffCommits_info_235_rfWen = io_diffCommits_info_235_rfWen;
        //    mon_tr.io_diffCommits_info_235_fpWen = io_diffCommits_info_235_fpWen;
        //    mon_tr.io_diffCommits_info_235_vecWen = io_diffCommits_info_235_vecWen;
        //    mon_tr.io_diffCommits_info_235_v0Wen = io_diffCommits_info_235_v0Wen;
        //    mon_tr.io_diffCommits_info_235_vlWen = io_diffCommits_info_235_vlWen;
        //    mon_tr.io_diffCommits_info_236_ldest = io_diffCommits_info_236_ldest;
        //    mon_tr.io_diffCommits_info_236_pdest = io_diffCommits_info_236_pdest;
        //    mon_tr.io_diffCommits_info_236_rfWen = io_diffCommits_info_236_rfWen;
        //    mon_tr.io_diffCommits_info_236_fpWen = io_diffCommits_info_236_fpWen;
        //    mon_tr.io_diffCommits_info_236_vecWen = io_diffCommits_info_236_vecWen;
        //    mon_tr.io_diffCommits_info_236_v0Wen = io_diffCommits_info_236_v0Wen;
        //    mon_tr.io_diffCommits_info_236_vlWen = io_diffCommits_info_236_vlWen;
        //    mon_tr.io_diffCommits_info_237_ldest = io_diffCommits_info_237_ldest;
        //    mon_tr.io_diffCommits_info_237_pdest = io_diffCommits_info_237_pdest;
        //    mon_tr.io_diffCommits_info_237_rfWen = io_diffCommits_info_237_rfWen;
        //    mon_tr.io_diffCommits_info_237_fpWen = io_diffCommits_info_237_fpWen;
        //    mon_tr.io_diffCommits_info_237_vecWen = io_diffCommits_info_237_vecWen;
        //    mon_tr.io_diffCommits_info_237_v0Wen = io_diffCommits_info_237_v0Wen;
        //    mon_tr.io_diffCommits_info_237_vlWen = io_diffCommits_info_237_vlWen;
        //    mon_tr.io_diffCommits_info_238_ldest = io_diffCommits_info_238_ldest;
        //    mon_tr.io_diffCommits_info_238_pdest = io_diffCommits_info_238_pdest;
        //    mon_tr.io_diffCommits_info_238_rfWen = io_diffCommits_info_238_rfWen;
        //    mon_tr.io_diffCommits_info_238_fpWen = io_diffCommits_info_238_fpWen;
        //    mon_tr.io_diffCommits_info_238_vecWen = io_diffCommits_info_238_vecWen;
        //    mon_tr.io_diffCommits_info_238_v0Wen = io_diffCommits_info_238_v0Wen;
        //    mon_tr.io_diffCommits_info_238_vlWen = io_diffCommits_info_238_vlWen;
        //    mon_tr.io_diffCommits_info_239_ldest = io_diffCommits_info_239_ldest;
        //    mon_tr.io_diffCommits_info_239_pdest = io_diffCommits_info_239_pdest;
        //    mon_tr.io_diffCommits_info_239_rfWen = io_diffCommits_info_239_rfWen;
        //    mon_tr.io_diffCommits_info_239_fpWen = io_diffCommits_info_239_fpWen;
        //    mon_tr.io_diffCommits_info_239_vecWen = io_diffCommits_info_239_vecWen;
        //    mon_tr.io_diffCommits_info_239_v0Wen = io_diffCommits_info_239_v0Wen;
        //    mon_tr.io_diffCommits_info_239_vlWen = io_diffCommits_info_239_vlWen;
        //    mon_tr.io_diffCommits_info_240_ldest = io_diffCommits_info_240_ldest;
        //    mon_tr.io_diffCommits_info_240_pdest = io_diffCommits_info_240_pdest;
        //    mon_tr.io_diffCommits_info_240_rfWen = io_diffCommits_info_240_rfWen;
        //    mon_tr.io_diffCommits_info_240_fpWen = io_diffCommits_info_240_fpWen;
        //    mon_tr.io_diffCommits_info_240_vecWen = io_diffCommits_info_240_vecWen;
        //    mon_tr.io_diffCommits_info_240_v0Wen = io_diffCommits_info_240_v0Wen;
        //    mon_tr.io_diffCommits_info_240_vlWen = io_diffCommits_info_240_vlWen;
        //    mon_tr.io_diffCommits_info_241_ldest = io_diffCommits_info_241_ldest;
        //    mon_tr.io_diffCommits_info_241_pdest = io_diffCommits_info_241_pdest;
        //    mon_tr.io_diffCommits_info_241_rfWen = io_diffCommits_info_241_rfWen;
        //    mon_tr.io_diffCommits_info_241_fpWen = io_diffCommits_info_241_fpWen;
        //    mon_tr.io_diffCommits_info_241_vecWen = io_diffCommits_info_241_vecWen;
        //    mon_tr.io_diffCommits_info_241_v0Wen = io_diffCommits_info_241_v0Wen;
        //    mon_tr.io_diffCommits_info_241_vlWen = io_diffCommits_info_241_vlWen;
        //    mon_tr.io_diffCommits_info_242_ldest = io_diffCommits_info_242_ldest;
        //    mon_tr.io_diffCommits_info_242_pdest = io_diffCommits_info_242_pdest;
        //    mon_tr.io_diffCommits_info_242_rfWen = io_diffCommits_info_242_rfWen;
        //    mon_tr.io_diffCommits_info_242_fpWen = io_diffCommits_info_242_fpWen;
        //    mon_tr.io_diffCommits_info_242_vecWen = io_diffCommits_info_242_vecWen;
        //    mon_tr.io_diffCommits_info_242_v0Wen = io_diffCommits_info_242_v0Wen;
        //    mon_tr.io_diffCommits_info_242_vlWen = io_diffCommits_info_242_vlWen;
        //    mon_tr.io_diffCommits_info_243_ldest = io_diffCommits_info_243_ldest;
        //    mon_tr.io_diffCommits_info_243_pdest = io_diffCommits_info_243_pdest;
        //    mon_tr.io_diffCommits_info_243_rfWen = io_diffCommits_info_243_rfWen;
        //    mon_tr.io_diffCommits_info_243_fpWen = io_diffCommits_info_243_fpWen;
        //    mon_tr.io_diffCommits_info_243_vecWen = io_diffCommits_info_243_vecWen;
        //    mon_tr.io_diffCommits_info_243_v0Wen = io_diffCommits_info_243_v0Wen;
        //    mon_tr.io_diffCommits_info_243_vlWen = io_diffCommits_info_243_vlWen;
        //    mon_tr.io_diffCommits_info_244_ldest = io_diffCommits_info_244_ldest;
        //    mon_tr.io_diffCommits_info_244_pdest = io_diffCommits_info_244_pdest;
        //    mon_tr.io_diffCommits_info_244_rfWen = io_diffCommits_info_244_rfWen;
        //    mon_tr.io_diffCommits_info_244_fpWen = io_diffCommits_info_244_fpWen;
        //    mon_tr.io_diffCommits_info_244_vecWen = io_diffCommits_info_244_vecWen;
        //    mon_tr.io_diffCommits_info_244_v0Wen = io_diffCommits_info_244_v0Wen;
        //    mon_tr.io_diffCommits_info_244_vlWen = io_diffCommits_info_244_vlWen;
        //    mon_tr.io_diffCommits_info_245_ldest = io_diffCommits_info_245_ldest;
        //    mon_tr.io_diffCommits_info_245_pdest = io_diffCommits_info_245_pdest;
        //    mon_tr.io_diffCommits_info_245_rfWen = io_diffCommits_info_245_rfWen;
        //    mon_tr.io_diffCommits_info_245_fpWen = io_diffCommits_info_245_fpWen;
        //    mon_tr.io_diffCommits_info_245_vecWen = io_diffCommits_info_245_vecWen;
        //    mon_tr.io_diffCommits_info_245_v0Wen = io_diffCommits_info_245_v0Wen;
        //    mon_tr.io_diffCommits_info_245_vlWen = io_diffCommits_info_245_vlWen;
        //    mon_tr.io_diffCommits_info_246_ldest = io_diffCommits_info_246_ldest;
        //    mon_tr.io_diffCommits_info_246_pdest = io_diffCommits_info_246_pdest;
        //    mon_tr.io_diffCommits_info_246_rfWen = io_diffCommits_info_246_rfWen;
        //    mon_tr.io_diffCommits_info_246_fpWen = io_diffCommits_info_246_fpWen;
        //    mon_tr.io_diffCommits_info_246_vecWen = io_diffCommits_info_246_vecWen;
        //    mon_tr.io_diffCommits_info_246_v0Wen = io_diffCommits_info_246_v0Wen;
        //    mon_tr.io_diffCommits_info_246_vlWen = io_diffCommits_info_246_vlWen;
        //    mon_tr.io_diffCommits_info_247_ldest = io_diffCommits_info_247_ldest;
        //    mon_tr.io_diffCommits_info_247_pdest = io_diffCommits_info_247_pdest;
        //    mon_tr.io_diffCommits_info_247_rfWen = io_diffCommits_info_247_rfWen;
        //    mon_tr.io_diffCommits_info_247_fpWen = io_diffCommits_info_247_fpWen;
        //    mon_tr.io_diffCommits_info_247_vecWen = io_diffCommits_info_247_vecWen;
        //    mon_tr.io_diffCommits_info_247_v0Wen = io_diffCommits_info_247_v0Wen;
        //    mon_tr.io_diffCommits_info_247_vlWen = io_diffCommits_info_247_vlWen;
        //    mon_tr.io_diffCommits_info_248_ldest = io_diffCommits_info_248_ldest;
        //    mon_tr.io_diffCommits_info_248_pdest = io_diffCommits_info_248_pdest;
        //    mon_tr.io_diffCommits_info_248_rfWen = io_diffCommits_info_248_rfWen;
        //    mon_tr.io_diffCommits_info_248_fpWen = io_diffCommits_info_248_fpWen;
        //    mon_tr.io_diffCommits_info_248_vecWen = io_diffCommits_info_248_vecWen;
        //    mon_tr.io_diffCommits_info_248_v0Wen = io_diffCommits_info_248_v0Wen;
        //    mon_tr.io_diffCommits_info_248_vlWen = io_diffCommits_info_248_vlWen;
        //    mon_tr.io_diffCommits_info_249_ldest = io_diffCommits_info_249_ldest;
        //    mon_tr.io_diffCommits_info_249_pdest = io_diffCommits_info_249_pdest;
        //    mon_tr.io_diffCommits_info_249_rfWen = io_diffCommits_info_249_rfWen;
        //    mon_tr.io_diffCommits_info_249_fpWen = io_diffCommits_info_249_fpWen;
        //    mon_tr.io_diffCommits_info_249_vecWen = io_diffCommits_info_249_vecWen;
        //    mon_tr.io_diffCommits_info_249_v0Wen = io_diffCommits_info_249_v0Wen;
        //    mon_tr.io_diffCommits_info_249_vlWen = io_diffCommits_info_249_vlWen;
        //    mon_tr.io_diffCommits_info_250_ldest = io_diffCommits_info_250_ldest;
        //    mon_tr.io_diffCommits_info_250_pdest = io_diffCommits_info_250_pdest;
        //    mon_tr.io_diffCommits_info_250_rfWen = io_diffCommits_info_250_rfWen;
        //    mon_tr.io_diffCommits_info_250_fpWen = io_diffCommits_info_250_fpWen;
        //    mon_tr.io_diffCommits_info_250_vecWen = io_diffCommits_info_250_vecWen;
        //    mon_tr.io_diffCommits_info_250_v0Wen = io_diffCommits_info_250_v0Wen;
        //    mon_tr.io_diffCommits_info_250_vlWen = io_diffCommits_info_250_vlWen;
        //    mon_tr.io_diffCommits_info_251_ldest = io_diffCommits_info_251_ldest;
        //    mon_tr.io_diffCommits_info_251_pdest = io_diffCommits_info_251_pdest;
        //    mon_tr.io_diffCommits_info_251_rfWen = io_diffCommits_info_251_rfWen;
        //    mon_tr.io_diffCommits_info_251_fpWen = io_diffCommits_info_251_fpWen;
        //    mon_tr.io_diffCommits_info_251_vecWen = io_diffCommits_info_251_vecWen;
        //    mon_tr.io_diffCommits_info_251_v0Wen = io_diffCommits_info_251_v0Wen;
        //    mon_tr.io_diffCommits_info_251_vlWen = io_diffCommits_info_251_vlWen;
        //    mon_tr.io_diffCommits_info_252_ldest = io_diffCommits_info_252_ldest;
        //    mon_tr.io_diffCommits_info_252_pdest = io_diffCommits_info_252_pdest;
        //    mon_tr.io_diffCommits_info_252_rfWen = io_diffCommits_info_252_rfWen;
        //    mon_tr.io_diffCommits_info_252_fpWen = io_diffCommits_info_252_fpWen;
        //    mon_tr.io_diffCommits_info_252_vecWen = io_diffCommits_info_252_vecWen;
        //    mon_tr.io_diffCommits_info_252_v0Wen = io_diffCommits_info_252_v0Wen;
        //    mon_tr.io_diffCommits_info_252_vlWen = io_diffCommits_info_252_vlWen;
        //    mon_tr.io_diffCommits_info_253_ldest = io_diffCommits_info_253_ldest;
        //    mon_tr.io_diffCommits_info_253_pdest = io_diffCommits_info_253_pdest;
        //    mon_tr.io_diffCommits_info_253_rfWen = io_diffCommits_info_253_rfWen;
        //    mon_tr.io_diffCommits_info_253_fpWen = io_diffCommits_info_253_fpWen;
        //    mon_tr.io_diffCommits_info_253_vecWen = io_diffCommits_info_253_vecWen;
        //    mon_tr.io_diffCommits_info_253_v0Wen = io_diffCommits_info_253_v0Wen;
        //    mon_tr.io_diffCommits_info_253_vlWen = io_diffCommits_info_253_vlWen;
        //    mon_tr.io_diffCommits_info_254_ldest = io_diffCommits_info_254_ldest;
        //    mon_tr.io_diffCommits_info_254_pdest = io_diffCommits_info_254_pdest;
        //    mon_tr.io_diffCommits_info_254_rfWen = io_diffCommits_info_254_rfWen;
        //    mon_tr.io_diffCommits_info_254_fpWen = io_diffCommits_info_254_fpWen;
        //    mon_tr.io_diffCommits_info_254_vecWen = io_diffCommits_info_254_vecWen;
        //    mon_tr.io_diffCommits_info_254_v0Wen = io_diffCommits_info_254_v0Wen;
        //    mon_tr.io_diffCommits_info_254_vlWen = io_diffCommits_info_254_vlWen;
        //    mon_tr.io_diffCommits_info_255_ldest = io_diffCommits_info_255_ldest;
        //    mon_tr.io_diffCommits_info_255_pdest = io_diffCommits_info_255_pdest;
        //    mon_tr.io_diffCommits_info_256_ldest = io_diffCommits_info_256_ldest;
        //    mon_tr.io_diffCommits_info_256_pdest = io_diffCommits_info_256_pdest;
        //    mon_tr.io_diffCommits_info_257_ldest = io_diffCommits_info_257_ldest;
        //    mon_tr.io_diffCommits_info_257_pdest = io_diffCommits_info_257_pdest;
        //    mon_tr.io_diffCommits_info_258_ldest = io_diffCommits_info_258_ldest;
        //    mon_tr.io_diffCommits_info_258_pdest = io_diffCommits_info_258_pdest;
        //    mon_tr.io_diffCommits_info_259_ldest = io_diffCommits_info_259_ldest;
        //    mon_tr.io_diffCommits_info_259_pdest = io_diffCommits_info_259_pdest;
        //    mon_tr.io_diffCommits_info_260_ldest = io_diffCommits_info_260_ldest;
        //    mon_tr.io_diffCommits_info_260_pdest = io_diffCommits_info_260_pdest;
        //    mon_tr.io_diffCommits_info_261_ldest = io_diffCommits_info_261_ldest;
        //    mon_tr.io_diffCommits_info_261_pdest = io_diffCommits_info_261_pdest;
        //    mon_tr.io_diffCommits_info_262_ldest = io_diffCommits_info_262_ldest;
        //    mon_tr.io_diffCommits_info_262_pdest = io_diffCommits_info_262_pdest;
        //    mon_tr.io_diffCommits_info_263_ldest = io_diffCommits_info_263_ldest;
        //    mon_tr.io_diffCommits_info_263_pdest = io_diffCommits_info_263_pdest;
        //    mon_tr.io_diffCommits_info_264_ldest = io_diffCommits_info_264_ldest;
        //    mon_tr.io_diffCommits_info_264_pdest = io_diffCommits_info_264_pdest;
        //    mon_tr.io_diffCommits_info_265_ldest = io_diffCommits_info_265_ldest;
        //    mon_tr.io_diffCommits_info_265_pdest = io_diffCommits_info_265_pdest;
        //    mon_tr.io_diffCommits_info_266_ldest = io_diffCommits_info_266_ldest;
        //    mon_tr.io_diffCommits_info_266_pdest = io_diffCommits_info_266_pdest;
        //    mon_tr.io_diffCommits_info_267_ldest = io_diffCommits_info_267_ldest;
        //    mon_tr.io_diffCommits_info_267_pdest = io_diffCommits_info_267_pdest;
        //    mon_tr.io_diffCommits_info_268_ldest = io_diffCommits_info_268_ldest;
        //    mon_tr.io_diffCommits_info_268_pdest = io_diffCommits_info_268_pdest;
        //    mon_tr.io_diffCommits_info_269_ldest = io_diffCommits_info_269_ldest;
        //    mon_tr.io_diffCommits_info_269_pdest = io_diffCommits_info_269_pdest;
        //    mon_tr.io_diffCommits_info_270_ldest = io_diffCommits_info_270_ldest;
        //    mon_tr.io_diffCommits_info_270_pdest = io_diffCommits_info_270_pdest;
        //    mon_tr.io_diffCommits_info_271_ldest = io_diffCommits_info_271_ldest;
        //    mon_tr.io_diffCommits_info_271_pdest = io_diffCommits_info_271_pdest;
        //    mon_tr.io_diffCommits_info_272_ldest = io_diffCommits_info_272_ldest;
        //    mon_tr.io_diffCommits_info_272_pdest = io_diffCommits_info_272_pdest;
        //    mon_tr.io_diffCommits_info_273_ldest = io_diffCommits_info_273_ldest;
        //    mon_tr.io_diffCommits_info_273_pdest = io_diffCommits_info_273_pdest;
        //    mon_tr.io_diffCommits_info_274_ldest = io_diffCommits_info_274_ldest;
        //    mon_tr.io_diffCommits_info_274_pdest = io_diffCommits_info_274_pdest;
        //    mon_tr.io_diffCommits_info_275_ldest = io_diffCommits_info_275_ldest;
        //    mon_tr.io_diffCommits_info_275_pdest = io_diffCommits_info_275_pdest;
        //    mon_tr.io_diffCommits_info_276_ldest = io_diffCommits_info_276_ldest;
        //    mon_tr.io_diffCommits_info_276_pdest = io_diffCommits_info_276_pdest;
        //    mon_tr.io_diffCommits_info_277_ldest = io_diffCommits_info_277_ldest;
        //    mon_tr.io_diffCommits_info_277_pdest = io_diffCommits_info_277_pdest;
        //    mon_tr.io_diffCommits_info_278_ldest = io_diffCommits_info_278_ldest;
        //    mon_tr.io_diffCommits_info_278_pdest = io_diffCommits_info_278_pdest;
        //    mon_tr.io_diffCommits_info_279_ldest = io_diffCommits_info_279_ldest;
        //    mon_tr.io_diffCommits_info_279_pdest = io_diffCommits_info_279_pdest;
        //    mon_tr.io_diffCommits_info_280_ldest = io_diffCommits_info_280_ldest;
        //    mon_tr.io_diffCommits_info_280_pdest = io_diffCommits_info_280_pdest;
        //    mon_tr.io_diffCommits_info_281_ldest = io_diffCommits_info_281_ldest;
        //    mon_tr.io_diffCommits_info_281_pdest = io_diffCommits_info_281_pdest;
        //    mon_tr.io_diffCommits_info_282_ldest = io_diffCommits_info_282_ldest;
        //    mon_tr.io_diffCommits_info_282_pdest = io_diffCommits_info_282_pdest;
        //    mon_tr.io_diffCommits_info_283_ldest = io_diffCommits_info_283_ldest;
        //    mon_tr.io_diffCommits_info_283_pdest = io_diffCommits_info_283_pdest;
        //    mon_tr.io_diffCommits_info_284_ldest = io_diffCommits_info_284_ldest;
        //    mon_tr.io_diffCommits_info_284_pdest = io_diffCommits_info_284_pdest;
        //    mon_tr.io_diffCommits_info_285_ldest = io_diffCommits_info_285_ldest;
        //    mon_tr.io_diffCommits_info_285_pdest = io_diffCommits_info_285_pdest;
        //    mon_tr.io_diffCommits_info_286_ldest = io_diffCommits_info_286_ldest;
        //    mon_tr.io_diffCommits_info_286_pdest = io_diffCommits_info_286_pdest;
        //    mon_tr.io_diffCommits_info_287_ldest = io_diffCommits_info_287_ldest;
        //    mon_tr.io_diffCommits_info_287_pdest = io_diffCommits_info_287_pdest;
        //    mon_tr.io_diffCommits_info_288_ldest = io_diffCommits_info_288_ldest;
        //    mon_tr.io_diffCommits_info_288_pdest = io_diffCommits_info_288_pdest;
        //    mon_tr.io_diffCommits_info_289_ldest = io_diffCommits_info_289_ldest;
        //    mon_tr.io_diffCommits_info_289_pdest = io_diffCommits_info_289_pdest;
        //    mon_tr.io_diffCommits_info_290_ldest = io_diffCommits_info_290_ldest;
        //    mon_tr.io_diffCommits_info_290_pdest = io_diffCommits_info_290_pdest;
        //    mon_tr.io_diffCommits_info_291_ldest = io_diffCommits_info_291_ldest;
        //    mon_tr.io_diffCommits_info_291_pdest = io_diffCommits_info_291_pdest;
        //    mon_tr.io_diffCommits_info_292_ldest = io_diffCommits_info_292_ldest;
        //    mon_tr.io_diffCommits_info_292_pdest = io_diffCommits_info_292_pdest;
        //    mon_tr.io_diffCommits_info_293_ldest = io_diffCommits_info_293_ldest;
        //    mon_tr.io_diffCommits_info_293_pdest = io_diffCommits_info_293_pdest;
        //    mon_tr.io_diffCommits_info_294_ldest = io_diffCommits_info_294_ldest;
        //    mon_tr.io_diffCommits_info_294_pdest = io_diffCommits_info_294_pdest;
        //    mon_tr.io_diffCommits_info_295_ldest = io_diffCommits_info_295_ldest;
        //    mon_tr.io_diffCommits_info_295_pdest = io_diffCommits_info_295_pdest;
        //    mon_tr.io_diffCommits_info_296_ldest = io_diffCommits_info_296_ldest;
        //    mon_tr.io_diffCommits_info_296_pdest = io_diffCommits_info_296_pdest;
        //    mon_tr.io_diffCommits_info_297_ldest = io_diffCommits_info_297_ldest;
        //    mon_tr.io_diffCommits_info_297_pdest = io_diffCommits_info_297_pdest;
        //    mon_tr.io_diffCommits_info_298_ldest = io_diffCommits_info_298_ldest;
        //    mon_tr.io_diffCommits_info_298_pdest = io_diffCommits_info_298_pdest;
        //    mon_tr.io_diffCommits_info_299_ldest = io_diffCommits_info_299_ldest;
        //    mon_tr.io_diffCommits_info_299_pdest = io_diffCommits_info_299_pdest;
        //    mon_tr.io_diffCommits_info_300_ldest = io_diffCommits_info_300_ldest;
        //    mon_tr.io_diffCommits_info_300_pdest = io_diffCommits_info_300_pdest;
        //    mon_tr.io_diffCommits_info_301_ldest = io_diffCommits_info_301_ldest;
        //    mon_tr.io_diffCommits_info_301_pdest = io_diffCommits_info_301_pdest;
        //    mon_tr.io_diffCommits_info_302_ldest = io_diffCommits_info_302_ldest;
        //    mon_tr.io_diffCommits_info_302_pdest = io_diffCommits_info_302_pdest;
        //    mon_tr.io_diffCommits_info_303_ldest = io_diffCommits_info_303_ldest;
        //    mon_tr.io_diffCommits_info_303_pdest = io_diffCommits_info_303_pdest;
        //    mon_tr.io_diffCommits_info_304_ldest = io_diffCommits_info_304_ldest;
        //    mon_tr.io_diffCommits_info_304_pdest = io_diffCommits_info_304_pdest;
        //    mon_tr.io_diffCommits_info_305_ldest = io_diffCommits_info_305_ldest;
        //    mon_tr.io_diffCommits_info_305_pdest = io_diffCommits_info_305_pdest;
        //    mon_tr.io_diffCommits_info_306_ldest = io_diffCommits_info_306_ldest;
        //    mon_tr.io_diffCommits_info_306_pdest = io_diffCommits_info_306_pdest;
        //    mon_tr.io_diffCommits_info_307_ldest = io_diffCommits_info_307_ldest;
        //    mon_tr.io_diffCommits_info_307_pdest = io_diffCommits_info_307_pdest;
        //    mon_tr.io_diffCommits_info_308_ldest = io_diffCommits_info_308_ldest;
        //    mon_tr.io_diffCommits_info_308_pdest = io_diffCommits_info_308_pdest;
        //    mon_tr.io_diffCommits_info_309_ldest = io_diffCommits_info_309_ldest;
        //    mon_tr.io_diffCommits_info_309_pdest = io_diffCommits_info_309_pdest;
        //    mon_tr.io_diffCommits_info_310_ldest = io_diffCommits_info_310_ldest;
        //    mon_tr.io_diffCommits_info_310_pdest = io_diffCommits_info_310_pdest;
        //    mon_tr.io_diffCommits_info_311_ldest = io_diffCommits_info_311_ldest;
        //    mon_tr.io_diffCommits_info_311_pdest = io_diffCommits_info_311_pdest;
        //    mon_tr.io_diffCommits_info_312_ldest = io_diffCommits_info_312_ldest;
        //    mon_tr.io_diffCommits_info_312_pdest = io_diffCommits_info_312_pdest;
        //    mon_tr.io_diffCommits_info_313_ldest = io_diffCommits_info_313_ldest;
        //    mon_tr.io_diffCommits_info_313_pdest = io_diffCommits_info_313_pdest;
        //    mon_tr.io_diffCommits_info_314_ldest = io_diffCommits_info_314_ldest;
        //    mon_tr.io_diffCommits_info_314_pdest = io_diffCommits_info_314_pdest;
        //    mon_tr.io_diffCommits_info_315_ldest = io_diffCommits_info_315_ldest;
        //    mon_tr.io_diffCommits_info_315_pdest = io_diffCommits_info_315_pdest;
        //    mon_tr.io_diffCommits_info_316_ldest = io_diffCommits_info_316_ldest;
        //    mon_tr.io_diffCommits_info_316_pdest = io_diffCommits_info_316_pdest;
        //    mon_tr.io_diffCommits_info_317_ldest = io_diffCommits_info_317_ldest;
        //    mon_tr.io_diffCommits_info_317_pdest = io_diffCommits_info_317_pdest;
        //    mon_tr.io_diffCommits_info_318_ldest = io_diffCommits_info_318_ldest;
        //    mon_tr.io_diffCommits_info_318_pdest = io_diffCommits_info_318_pdest;
        //    mon_tr.io_diffCommits_info_319_ldest = io_diffCommits_info_319_ldest;
        //    mon_tr.io_diffCommits_info_319_pdest = io_diffCommits_info_319_pdest;
        //    mon_tr.io_diffCommits_info_320_ldest = io_diffCommits_info_320_ldest;
        //    mon_tr.io_diffCommits_info_320_pdest = io_diffCommits_info_320_pdest;
        //    mon_tr.io_diffCommits_info_321_ldest = io_diffCommits_info_321_ldest;
        //    mon_tr.io_diffCommits_info_321_pdest = io_diffCommits_info_321_pdest;
        //    mon_tr.io_diffCommits_info_322_ldest = io_diffCommits_info_322_ldest;
        //    mon_tr.io_diffCommits_info_322_pdest = io_diffCommits_info_322_pdest;
        //    mon_tr.io_diffCommits_info_323_ldest = io_diffCommits_info_323_ldest;
        //    mon_tr.io_diffCommits_info_323_pdest = io_diffCommits_info_323_pdest;
        //    mon_tr.io_diffCommits_info_324_ldest = io_diffCommits_info_324_ldest;
        //    mon_tr.io_diffCommits_info_324_pdest = io_diffCommits_info_324_pdest;
        //    mon_tr.io_diffCommits_info_325_ldest = io_diffCommits_info_325_ldest;
        //    mon_tr.io_diffCommits_info_325_pdest = io_diffCommits_info_325_pdest;
        //    mon_tr.io_diffCommits_info_326_ldest = io_diffCommits_info_326_ldest;
        //    mon_tr.io_diffCommits_info_326_pdest = io_diffCommits_info_326_pdest;
        //    mon_tr.io_diffCommits_info_327_ldest = io_diffCommits_info_327_ldest;
        //    mon_tr.io_diffCommits_info_327_pdest = io_diffCommits_info_327_pdest;
        //    mon_tr.io_diffCommits_info_328_ldest = io_diffCommits_info_328_ldest;
        //    mon_tr.io_diffCommits_info_328_pdest = io_diffCommits_info_328_pdest;
        //    mon_tr.io_diffCommits_info_329_ldest = io_diffCommits_info_329_ldest;
        //    mon_tr.io_diffCommits_info_329_pdest = io_diffCommits_info_329_pdest;
        //    mon_tr.io_diffCommits_info_330_ldest = io_diffCommits_info_330_ldest;
        //    mon_tr.io_diffCommits_info_330_pdest = io_diffCommits_info_330_pdest;
        //    mon_tr.io_diffCommits_info_331_ldest = io_diffCommits_info_331_ldest;
        //    mon_tr.io_diffCommits_info_331_pdest = io_diffCommits_info_331_pdest;
        //    mon_tr.io_diffCommits_info_332_ldest = io_diffCommits_info_332_ldest;
        //    mon_tr.io_diffCommits_info_332_pdest = io_diffCommits_info_332_pdest;
        //    mon_tr.io_diffCommits_info_333_ldest = io_diffCommits_info_333_ldest;
        //    mon_tr.io_diffCommits_info_333_pdest = io_diffCommits_info_333_pdest;
        //    mon_tr.io_diffCommits_info_334_ldest = io_diffCommits_info_334_ldest;
        //    mon_tr.io_diffCommits_info_334_pdest = io_diffCommits_info_334_pdest;
        //    mon_tr.io_diffCommits_info_335_ldest = io_diffCommits_info_335_ldest;
        //    mon_tr.io_diffCommits_info_335_pdest = io_diffCommits_info_335_pdest;
        //    mon_tr.io_diffCommits_info_336_ldest = io_diffCommits_info_336_ldest;
        //    mon_tr.io_diffCommits_info_336_pdest = io_diffCommits_info_336_pdest;
        //    mon_tr.io_diffCommits_info_337_ldest = io_diffCommits_info_337_ldest;
        //    mon_tr.io_diffCommits_info_337_pdest = io_diffCommits_info_337_pdest;
        //    mon_tr.io_diffCommits_info_338_ldest = io_diffCommits_info_338_ldest;
        //    mon_tr.io_diffCommits_info_338_pdest = io_diffCommits_info_338_pdest;
        //    mon_tr.io_diffCommits_info_339_ldest = io_diffCommits_info_339_ldest;
        //    mon_tr.io_diffCommits_info_339_pdest = io_diffCommits_info_339_pdest;
        //    mon_tr.io_diffCommits_info_340_ldest = io_diffCommits_info_340_ldest;
        //    mon_tr.io_diffCommits_info_340_pdest = io_diffCommits_info_340_pdest;
        //    mon_tr.io_diffCommits_info_341_ldest = io_diffCommits_info_341_ldest;
        //    mon_tr.io_diffCommits_info_341_pdest = io_diffCommits_info_341_pdest;
        //    mon_tr.io_diffCommits_info_342_ldest = io_diffCommits_info_342_ldest;
        //    mon_tr.io_diffCommits_info_342_pdest = io_diffCommits_info_342_pdest;
        //    mon_tr.io_diffCommits_info_343_ldest = io_diffCommits_info_343_ldest;
        //    mon_tr.io_diffCommits_info_343_pdest = io_diffCommits_info_343_pdest;
        //    mon_tr.io_diffCommits_info_344_ldest = io_diffCommits_info_344_ldest;
        //    mon_tr.io_diffCommits_info_344_pdest = io_diffCommits_info_344_pdest;
        //    mon_tr.io_diffCommits_info_345_ldest = io_diffCommits_info_345_ldest;
        //    mon_tr.io_diffCommits_info_345_pdest = io_diffCommits_info_345_pdest;
        //    mon_tr.io_diffCommits_info_346_ldest = io_diffCommits_info_346_ldest;
        //    mon_tr.io_diffCommits_info_346_pdest = io_diffCommits_info_346_pdest;
        //    mon_tr.io_diffCommits_info_347_ldest = io_diffCommits_info_347_ldest;
        //    mon_tr.io_diffCommits_info_347_pdest = io_diffCommits_info_347_pdest;
        //    mon_tr.io_diffCommits_info_348_ldest = io_diffCommits_info_348_ldest;
        //    mon_tr.io_diffCommits_info_348_pdest = io_diffCommits_info_348_pdest;
        //    mon_tr.io_diffCommits_info_349_ldest = io_diffCommits_info_349_ldest;
        //    mon_tr.io_diffCommits_info_349_pdest = io_diffCommits_info_349_pdest;
        //    mon_tr.io_diffCommits_info_350_ldest = io_diffCommits_info_350_ldest;
        //    mon_tr.io_diffCommits_info_350_pdest = io_diffCommits_info_350_pdest;
        //    mon_tr.io_diffCommits_info_351_ldest = io_diffCommits_info_351_ldest;
        //    mon_tr.io_diffCommits_info_351_pdest = io_diffCommits_info_351_pdest;
        //    mon_tr.io_diffCommits_info_352_ldest = io_diffCommits_info_352_ldest;
        //    mon_tr.io_diffCommits_info_352_pdest = io_diffCommits_info_352_pdest;
        //    mon_tr.io_diffCommits_info_353_ldest = io_diffCommits_info_353_ldest;
        //    mon_tr.io_diffCommits_info_353_pdest = io_diffCommits_info_353_pdest;
        //    mon_tr.io_diffCommits_info_354_ldest = io_diffCommits_info_354_ldest;
        //    mon_tr.io_diffCommits_info_354_pdest = io_diffCommits_info_354_pdest;
        //    mon_tr.io_diffCommits_info_355_ldest = io_diffCommits_info_355_ldest;
        //    mon_tr.io_diffCommits_info_355_pdest = io_diffCommits_info_355_pdest;
        //    mon_tr.io_diffCommits_info_356_ldest = io_diffCommits_info_356_ldest;
        //    mon_tr.io_diffCommits_info_356_pdest = io_diffCommits_info_356_pdest;
        //    mon_tr.io_diffCommits_info_357_ldest = io_diffCommits_info_357_ldest;
        //    mon_tr.io_diffCommits_info_357_pdest = io_diffCommits_info_357_pdest;
        //    mon_tr.io_diffCommits_info_358_ldest = io_diffCommits_info_358_ldest;
        //    mon_tr.io_diffCommits_info_358_pdest = io_diffCommits_info_358_pdest;
        //    mon_tr.io_diffCommits_info_359_ldest = io_diffCommits_info_359_ldest;
        //    mon_tr.io_diffCommits_info_359_pdest = io_diffCommits_info_359_pdest;
        //    mon_tr.io_diffCommits_info_360_ldest = io_diffCommits_info_360_ldest;
        //    mon_tr.io_diffCommits_info_360_pdest = io_diffCommits_info_360_pdest;
        //    mon_tr.io_diffCommits_info_361_ldest = io_diffCommits_info_361_ldest;
        //    mon_tr.io_diffCommits_info_361_pdest = io_diffCommits_info_361_pdest;
        //    mon_tr.io_diffCommits_info_362_ldest = io_diffCommits_info_362_ldest;
        //    mon_tr.io_diffCommits_info_362_pdest = io_diffCommits_info_362_pdest;
        //    mon_tr.io_diffCommits_info_363_ldest = io_diffCommits_info_363_ldest;
        //    mon_tr.io_diffCommits_info_363_pdest = io_diffCommits_info_363_pdest;
        //    mon_tr.io_diffCommits_info_364_ldest = io_diffCommits_info_364_ldest;
        //    mon_tr.io_diffCommits_info_364_pdest = io_diffCommits_info_364_pdest;
        //    mon_tr.io_diffCommits_info_365_ldest = io_diffCommits_info_365_ldest;
        //    mon_tr.io_diffCommits_info_365_pdest = io_diffCommits_info_365_pdest;
        //    mon_tr.io_diffCommits_info_366_ldest = io_diffCommits_info_366_ldest;
        //    mon_tr.io_diffCommits_info_366_pdest = io_diffCommits_info_366_pdest;
        //    mon_tr.io_diffCommits_info_367_ldest = io_diffCommits_info_367_ldest;
        //    mon_tr.io_diffCommits_info_367_pdest = io_diffCommits_info_367_pdest;
        //    mon_tr.io_diffCommits_info_368_ldest = io_diffCommits_info_368_ldest;
        //    mon_tr.io_diffCommits_info_368_pdest = io_diffCommits_info_368_pdest;
        //    mon_tr.io_diffCommits_info_369_ldest = io_diffCommits_info_369_ldest;
        //    mon_tr.io_diffCommits_info_369_pdest = io_diffCommits_info_369_pdest;
        //    mon_tr.io_diffCommits_info_370_ldest = io_diffCommits_info_370_ldest;
        //    mon_tr.io_diffCommits_info_370_pdest = io_diffCommits_info_370_pdest;
        //    mon_tr.io_diffCommits_info_371_ldest = io_diffCommits_info_371_ldest;
        //    mon_tr.io_diffCommits_info_371_pdest = io_diffCommits_info_371_pdest;
        //    mon_tr.io_diffCommits_info_372_ldest = io_diffCommits_info_372_ldest;
        //    mon_tr.io_diffCommits_info_372_pdest = io_diffCommits_info_372_pdest;
        //    mon_tr.io_diffCommits_info_373_ldest = io_diffCommits_info_373_ldest;
        //    mon_tr.io_diffCommits_info_373_pdest = io_diffCommits_info_373_pdest;
        //    mon_tr.io_diffCommits_info_374_ldest = io_diffCommits_info_374_ldest;
        //    mon_tr.io_diffCommits_info_374_pdest = io_diffCommits_info_374_pdest;
        //    mon_tr.io_diffCommits_info_375_ldest = io_diffCommits_info_375_ldest;
        //    mon_tr.io_diffCommits_info_375_pdest = io_diffCommits_info_375_pdest;
        //    mon_tr.io_diffCommits_info_376_ldest = io_diffCommits_info_376_ldest;
        //    mon_tr.io_diffCommits_info_376_pdest = io_diffCommits_info_376_pdest;
        //    mon_tr.io_diffCommits_info_377_ldest = io_diffCommits_info_377_ldest;
        //    mon_tr.io_diffCommits_info_377_pdest = io_diffCommits_info_377_pdest;
        //    mon_tr.io_diffCommits_info_378_ldest = io_diffCommits_info_378_ldest;
        //    mon_tr.io_diffCommits_info_378_pdest = io_diffCommits_info_378_pdest;
        //    mon_tr.io_diffCommits_info_379_ldest = io_diffCommits_info_379_ldest;
        //    mon_tr.io_diffCommits_info_379_pdest = io_diffCommits_info_379_pdest;
        //    mon_tr.io_diffCommits_info_380_ldest = io_diffCommits_info_380_ldest;
        //    mon_tr.io_diffCommits_info_380_pdest = io_diffCommits_info_380_pdest;
        //    mon_tr.io_diffCommits_info_381_ldest = io_diffCommits_info_381_ldest;
        //    mon_tr.io_diffCommits_info_381_pdest = io_diffCommits_info_381_pdest;
        //    mon_tr.io_diffCommits_info_382_ldest = io_diffCommits_info_382_ldest;
        //    mon_tr.io_diffCommits_info_382_pdest = io_diffCommits_info_382_pdest;
        //    mon_tr.io_diffCommits_info_383_ldest = io_diffCommits_info_383_ldest;
        //    mon_tr.io_diffCommits_info_383_pdest = io_diffCommits_info_383_pdest;
        //    mon_tr.io_diffCommits_info_384_ldest = io_diffCommits_info_384_ldest;
        //    mon_tr.io_diffCommits_info_384_pdest = io_diffCommits_info_384_pdest;
        //    mon_tr.io_diffCommits_info_385_ldest = io_diffCommits_info_385_ldest;
        //    mon_tr.io_diffCommits_info_385_pdest = io_diffCommits_info_385_pdest;
        //    mon_tr.io_diffCommits_info_386_ldest = io_diffCommits_info_386_ldest;
        //    mon_tr.io_diffCommits_info_386_pdest = io_diffCommits_info_386_pdest;
        //    mon_tr.io_diffCommits_info_387_ldest = io_diffCommits_info_387_ldest;
        //    mon_tr.io_diffCommits_info_387_pdest = io_diffCommits_info_387_pdest;
        //    mon_tr.io_diffCommits_info_388_ldest = io_diffCommits_info_388_ldest;
        //    mon_tr.io_diffCommits_info_388_pdest = io_diffCommits_info_388_pdest;
        //    mon_tr.io_diffCommits_info_389_ldest = io_diffCommits_info_389_ldest;
        //    mon_tr.io_diffCommits_info_389_pdest = io_diffCommits_info_389_pdest;
        //    mon_tr.io_lsq_scommit = io_lsq_scommit;
        //    mon_tr.io_lsq_pendingMMIOld = io_lsq_pendingMMIOld;
        //    mon_tr.io_lsq_pendingst = io_lsq_pendingst;
        //    mon_tr.io_lsq_pendingPtr_flag = io_lsq_pendingPtr_flag;
        //    mon_tr.io_lsq_pendingPtr_value = io_lsq_pendingPtr_value;
        //    mon_tr.io_robDeqPtr_flag = io_robDeqPtr_flag;
        //    mon_tr.io_robDeqPtr_value = io_robDeqPtr_value;
        //    mon_tr.io_csr_fflags_valid = io_csr_fflags_valid;
        //    mon_tr.io_csr_fflags_bits = io_csr_fflags_bits;
        //    mon_tr.io_csr_vxsat_valid = io_csr_vxsat_valid;
        //    mon_tr.io_csr_vxsat_bits = io_csr_vxsat_bits;
        //    mon_tr.io_csr_vstart_valid = io_csr_vstart_valid;
        //    mon_tr.io_csr_vstart_bits = io_csr_vstart_bits;
        //    mon_tr.io_csr_dirty_fs = io_csr_dirty_fs;
        //    mon_tr.io_csr_dirty_vs = io_csr_dirty_vs;
        //    mon_tr.io_csr_perfinfo_retiredInstr = io_csr_perfinfo_retiredInstr;
        //    mon_tr.io_cpu_halt = io_cpu_halt;
        //    mon_tr.io_wfi_wfiReq = io_wfi_wfiReq;
        //    mon_tr.io_toDecode_isResumeVType = io_toDecode_isResumeVType;
        //    mon_tr.io_toDecode_walkToArchVType = io_toDecode_walkToArchVType;
        //    mon_tr.io_toDecode_walkVType_valid = io_toDecode_walkVType_valid;
        //    mon_tr.io_toDecode_walkVType_bits_illegal = io_toDecode_walkVType_bits_illegal;
        //    mon_tr.io_toDecode_walkVType_bits_vma = io_toDecode_walkVType_bits_vma;
        //    mon_tr.io_toDecode_walkVType_bits_vta = io_toDecode_walkVType_bits_vta;
        //    mon_tr.io_toDecode_walkVType_bits_vsew = io_toDecode_walkVType_bits_vsew;
        //    mon_tr.io_toDecode_walkVType_bits_vlmul = io_toDecode_walkVType_bits_vlmul;
        //    mon_tr.io_toDecode_commitVType_vtype_valid = io_toDecode_commitVType_vtype_valid;
        //    mon_tr.io_toDecode_commitVType_vtype_bits_illegal = io_toDecode_commitVType_vtype_bits_illegal;
        //    mon_tr.io_toDecode_commitVType_vtype_bits_vma = io_toDecode_commitVType_vtype_bits_vma;
        //    mon_tr.io_toDecode_commitVType_vtype_bits_vta = io_toDecode_commitVType_vtype_bits_vta;
        //    mon_tr.io_toDecode_commitVType_vtype_bits_vsew = io_toDecode_commitVType_vtype_bits_vsew;
        //    mon_tr.io_toDecode_commitVType_vtype_bits_vlmul = io_toDecode_commitVType_vtype_bits_vlmul;
        //    mon_tr.io_toDecode_commitVType_hasVsetvl = io_toDecode_commitVType_hasVsetvl;
        //    mon_tr.io_readGPAMemAddr_valid = io_readGPAMemAddr_valid;
        //    mon_tr.io_readGPAMemAddr_bits_ftqPtr_value = io_readGPAMemAddr_bits_ftqPtr_value;
        //    mon_tr.io_readGPAMemAddr_bits_ftqOffset = io_readGPAMemAddr_bits_ftqOffset;
        //    mon_tr.io_toVecExcpMod_logicPhyRegMap_0_valid = io_toVecExcpMod_logicPhyRegMap_0_valid;
        //    mon_tr.io_toVecExcpMod_logicPhyRegMap_0_bits_lreg = io_toVecExcpMod_logicPhyRegMap_0_bits_lreg;
        //    mon_tr.io_toVecExcpMod_logicPhyRegMap_0_bits_preg = io_toVecExcpMod_logicPhyRegMap_0_bits_preg;
        //    mon_tr.io_toVecExcpMod_logicPhyRegMap_1_valid = io_toVecExcpMod_logicPhyRegMap_1_valid;
        //    mon_tr.io_toVecExcpMod_logicPhyRegMap_1_bits_lreg = io_toVecExcpMod_logicPhyRegMap_1_bits_lreg;
        //    mon_tr.io_toVecExcpMod_logicPhyRegMap_1_bits_preg = io_toVecExcpMod_logicPhyRegMap_1_bits_preg;
        //    mon_tr.io_toVecExcpMod_logicPhyRegMap_2_valid = io_toVecExcpMod_logicPhyRegMap_2_valid;
        //    mon_tr.io_toVecExcpMod_logicPhyRegMap_2_bits_lreg = io_toVecExcpMod_logicPhyRegMap_2_bits_lreg;
        //    mon_tr.io_toVecExcpMod_logicPhyRegMap_2_bits_preg = io_toVecExcpMod_logicPhyRegMap_2_bits_preg;
        //    mon_tr.io_toVecExcpMod_logicPhyRegMap_3_valid = io_toVecExcpMod_logicPhyRegMap_3_valid;
        //    mon_tr.io_toVecExcpMod_logicPhyRegMap_3_bits_lreg = io_toVecExcpMod_logicPhyRegMap_3_bits_lreg;
        //    mon_tr.io_toVecExcpMod_logicPhyRegMap_3_bits_preg = io_toVecExcpMod_logicPhyRegMap_3_bits_preg;
        //    mon_tr.io_toVecExcpMod_logicPhyRegMap_4_valid = io_toVecExcpMod_logicPhyRegMap_4_valid;
        //    mon_tr.io_toVecExcpMod_logicPhyRegMap_4_bits_lreg = io_toVecExcpMod_logicPhyRegMap_4_bits_lreg;
        //    mon_tr.io_toVecExcpMod_logicPhyRegMap_4_bits_preg = io_toVecExcpMod_logicPhyRegMap_4_bits_preg;
        //    mon_tr.io_toVecExcpMod_logicPhyRegMap_5_valid = io_toVecExcpMod_logicPhyRegMap_5_valid;
        //    mon_tr.io_toVecExcpMod_logicPhyRegMap_5_bits_lreg = io_toVecExcpMod_logicPhyRegMap_5_bits_lreg;
        //    mon_tr.io_toVecExcpMod_logicPhyRegMap_5_bits_preg = io_toVecExcpMod_logicPhyRegMap_5_bits_preg;
        //    mon_tr.io_toVecExcpMod_excpInfo_valid = io_toVecExcpMod_excpInfo_valid;
        //    mon_tr.io_toVecExcpMod_excpInfo_bits_vstart = io_toVecExcpMod_excpInfo_bits_vstart;
        //    mon_tr.io_toVecExcpMod_excpInfo_bits_vsew = io_toVecExcpMod_excpInfo_bits_vsew;
        //    mon_tr.io_toVecExcpMod_excpInfo_bits_veew = io_toVecExcpMod_excpInfo_bits_veew;
        //    mon_tr.io_toVecExcpMod_excpInfo_bits_vlmul = io_toVecExcpMod_excpInfo_bits_vlmul;
        //    mon_tr.io_toVecExcpMod_excpInfo_bits_nf = io_toVecExcpMod_excpInfo_bits_nf;
        //    mon_tr.io_toVecExcpMod_excpInfo_bits_isStride = io_toVecExcpMod_excpInfo_bits_isStride;
        //    mon_tr.io_toVecExcpMod_excpInfo_bits_isIndexed = io_toVecExcpMod_excpInfo_bits_isIndexed;
        //    mon_tr.io_toVecExcpMod_excpInfo_bits_isWhole = io_toVecExcpMod_excpInfo_bits_isWhole;
        //    mon_tr.io_toVecExcpMod_excpInfo_bits_isVlm = io_toVecExcpMod_excpInfo_bits_isVlm;
        //    mon_tr.io_storeDebugInfo_1_pc = io_storeDebugInfo_1_pc;
        //    mon_tr.io_perf_0_value = io_perf_0_value;
        //    mon_tr.io_perf_1_value = io_perf_1_value;
        //    mon_tr.io_perf_2_value = io_perf_2_value;
        //    mon_tr.io_perf_3_value = io_perf_3_value;
        //    mon_tr.io_perf_4_value = io_perf_4_value;
        //    mon_tr.io_perf_5_value = io_perf_5_value;
        //    mon_tr.io_perf_6_value = io_perf_6_value;
        //    mon_tr.io_perf_7_value = io_perf_7_value;
        //    mon_tr.io_perf_8_value = io_perf_8_value;
        //    mon_tr.io_perf_9_value = io_perf_9_value;
        //    mon_tr.io_perf_10_value = io_perf_10_value;
        //    mon_tr.io_perf_11_value = io_perf_11_value;
        //    mon_tr.io_perf_12_value = io_perf_12_value;
        //    mon_tr.io_perf_13_value = io_perf_13_value;
        //    mon_tr.io_perf_14_value = io_perf_14_value;
        //    mon_tr.io_perf_15_value = io_perf_15_value;
        //    mon_tr.io_perf_16_value = io_perf_16_value;
        //    mon_tr.io_perf_17_value = io_perf_17_value;
        //    mon_tr.io_error_0 = io_error_0;

        //    mon_tr.channel_id = this.cfg.channel_id;
        //    mon_tr.unpack();
        //    this.mon_item_port.write(mon_tr);
        //end
    end
endtask:mon_data

`endif


//=========================================================
//File name    : Rob_output_agent_dec.sv
//Author       : nanyunhao
//Module name  : Rob_output_agent_dec
//Discribution : Rob_output_agent_dec : parameter
//Date         : 2026-01-22
//=========================================================
`ifndef ROB_OUTPUT_AGENT_DEC__SV
`define ROB_OUTPUT_AGENT_DEC__SV

package Rob_output_agent_dec;

endpackage:Rob_output_agent_dec

import Rob_output_agent_dec::*;

`endif


//=========================================================
//File name    : Rob_output_agent_xaction.sv
//Author       : nanyunhao
//Module name  : Rob_output_agent_xaction
//Discribution : Rob_output_agent_xaction : agent transaction
//Date         : 2026-01-22
//=========================================================
`ifndef ROB_OUTPUT_AGENT_XACTION__SV
`define ROB_OUTPUT_AGENT_XACTION__SV

class Rob_output_agent_xaction  extends tcnt_data_base;
    rand bit         io_enq_canAccept  ;
    rand bit         io_enq_canAcceptForDispatch;
    rand bit         io_enq_isEmpty    ;
    rand bit         io_flushOut_valid ;
    rand bit         io_flushOut_bits_isRVC;
    rand bit         io_flushOut_bits_robIdx_flag;
    rand bit [7:0]   io_flushOut_bits_robIdx_value;
    rand bit         io_flushOut_bits_ftqIdx_flag;
    rand bit [5:0]   io_flushOut_bits_ftqIdx_value;
    rand bit [3:0]   io_flushOut_bits_ftqOffset;
    rand bit         io_flushOut_bits_level;
    rand bit         io_exception_valid;
    rand bit [31:0]  io_exception_bits_instr;
    rand bit [2:0]   io_exception_bits_commitType;
    rand bit         io_exception_bits_exceptionVec_0;
    rand bit         io_exception_bits_exceptionVec_1;
    rand bit         io_exception_bits_exceptionVec_2;
    rand bit         io_exception_bits_exceptionVec_3;
    rand bit         io_exception_bits_exceptionVec_4;
    rand bit         io_exception_bits_exceptionVec_5;
    rand bit         io_exception_bits_exceptionVec_6;
    rand bit         io_exception_bits_exceptionVec_7;
    rand bit         io_exception_bits_exceptionVec_8;
    rand bit         io_exception_bits_exceptionVec_9;
    rand bit         io_exception_bits_exceptionVec_10;
    rand bit         io_exception_bits_exceptionVec_11;
    rand bit         io_exception_bits_exceptionVec_12;
    rand bit         io_exception_bits_exceptionVec_13;
    rand bit         io_exception_bits_exceptionVec_14;
    rand bit         io_exception_bits_exceptionVec_15;
    rand bit         io_exception_bits_exceptionVec_16;
    rand bit         io_exception_bits_exceptionVec_17;
    rand bit         io_exception_bits_exceptionVec_18;
    rand bit         io_exception_bits_exceptionVec_19;
    rand bit         io_exception_bits_exceptionVec_20;
    rand bit         io_exception_bits_exceptionVec_21;
    rand bit         io_exception_bits_exceptionVec_22;
    rand bit         io_exception_bits_exceptionVec_23;
    rand bit         io_exception_bits_isPcBkpt;
    rand bit         io_exception_bits_isFetchMalAddr;
    rand bit [63:0]  io_exception_bits_gpaddr;
    rand bit         io_exception_bits_singleStep;
    rand bit         io_exception_bits_crossPageIPFFix;
    rand bit         io_exception_bits_isInterrupt;
    rand bit         io_exception_bits_isHls;
    rand bit [3:0]   io_exception_bits_trigger;
    rand bit         io_exception_bits_isForVSnonLeafPTE;
    rand bit         io_commits_isCommit;
    rand bit         io_commits_commitValid_0;
    rand bit         io_commits_commitValid_1;
    rand bit         io_commits_commitValid_2;
    rand bit         io_commits_commitValid_3;
    rand bit         io_commits_commitValid_4;
    rand bit         io_commits_commitValid_5;
    rand bit         io_commits_commitValid_6;
    rand bit         io_commits_commitValid_7;
    rand bit         io_commits_isWalk ;
    rand bit         io_commits_walkValid_0;
    rand bit         io_commits_walkValid_1;
    rand bit         io_commits_walkValid_2;
    rand bit         io_commits_walkValid_3;
    rand bit         io_commits_walkValid_4;
    rand bit         io_commits_walkValid_5;
    rand bit         io_commits_walkValid_6;
    rand bit         io_commits_walkValid_7;
    rand bit         io_commits_info_0_walk_v;
    rand bit         io_commits_info_0_commit_v;
    rand bit         io_commits_info_0_commit_w;
    rand bit [6:0]   io_commits_info_0_realDestSize;
    rand bit         io_commits_info_0_interrupt_safe;
    rand bit         io_commits_info_0_wflags;
    rand bit [4:0]   io_commits_info_0_fflags;
    rand bit         io_commits_info_0_vxsat;
    rand bit         io_commits_info_0_isRVC;
    rand bit         io_commits_info_0_isVset;
    rand bit         io_commits_info_0_isHls;
    rand bit         io_commits_info_0_isVls;
    rand bit         io_commits_info_0_vls;
    rand bit         io_commits_info_0_mmio;
    rand bit [2:0]   io_commits_info_0_commitType;
    rand bit         io_commits_info_0_ftqIdx_flag;
    rand bit [5:0]   io_commits_info_0_ftqIdx_value;
    rand bit [3:0]   io_commits_info_0_ftqOffset;
    rand bit [2:0]   io_commits_info_0_instrSize;
    rand bit         io_commits_info_0_fpWen;
    rand bit         io_commits_info_0_rfWen;
    rand bit         io_commits_info_0_needFlush;
    rand bit [3:0]   io_commits_info_0_traceBlockInPipe_itype;
    rand bit [3:0]   io_commits_info_0_traceBlockInPipe_iretire;
    rand bit         io_commits_info_0_traceBlockInPipe_ilastsize;
    rand bit [49:0]  io_commits_info_0_debug_pc;
    rand bit [31:0]  io_commits_info_0_debug_instr;
    rand bit [5:0]   io_commits_info_0_debug_ldest;
    rand bit [7:0]   io_commits_info_0_debug_pdest;
    rand bit [7:0]   io_commits_info_0_debug_otherPdest_0;
    rand bit [7:0]   io_commits_info_0_debug_otherPdest_1;
    rand bit [7:0]   io_commits_info_0_debug_otherPdest_2;
    rand bit [7:0]   io_commits_info_0_debug_otherPdest_3;
    rand bit [7:0]   io_commits_info_0_debug_otherPdest_4;
    rand bit [7:0]   io_commits_info_0_debug_otherPdest_5;
    rand bit [7:0]   io_commits_info_0_debug_otherPdest_6;
    rand bit [34:0]  io_commits_info_0_debug_fuType;
    rand bit         io_commits_info_0_dirtyFs;
    rand bit         io_commits_info_0_dirtyVs;
    rand bit         io_commits_info_1_walk_v;
    rand bit         io_commits_info_1_commit_v;
    rand bit         io_commits_info_1_commit_w;
    rand bit [6:0]   io_commits_info_1_realDestSize;
    rand bit         io_commits_info_1_interrupt_safe;
    rand bit         io_commits_info_1_wflags;
    rand bit [4:0]   io_commits_info_1_fflags;
    rand bit         io_commits_info_1_vxsat;
    rand bit         io_commits_info_1_isRVC;
    rand bit         io_commits_info_1_isVset;
    rand bit         io_commits_info_1_isHls;
    rand bit         io_commits_info_1_isVls;
    rand bit         io_commits_info_1_vls;
    rand bit         io_commits_info_1_mmio;
    rand bit [2:0]   io_commits_info_1_commitType;
    rand bit         io_commits_info_1_ftqIdx_flag;
    rand bit [5:0]   io_commits_info_1_ftqIdx_value;
    rand bit [3:0]   io_commits_info_1_ftqOffset;
    rand bit [2:0]   io_commits_info_1_instrSize;
    rand bit         io_commits_info_1_fpWen;
    rand bit         io_commits_info_1_rfWen;
    rand bit         io_commits_info_1_needFlush;
    rand bit [3:0]   io_commits_info_1_traceBlockInPipe_itype;
    rand bit [3:0]   io_commits_info_1_traceBlockInPipe_iretire;
    rand bit         io_commits_info_1_traceBlockInPipe_ilastsize;
    rand bit [49:0]  io_commits_info_1_debug_pc;
    rand bit [31:0]  io_commits_info_1_debug_instr;
    rand bit [5:0]   io_commits_info_1_debug_ldest;
    rand bit [7:0]   io_commits_info_1_debug_pdest;
    rand bit [7:0]   io_commits_info_1_debug_otherPdest_0;
    rand bit [7:0]   io_commits_info_1_debug_otherPdest_1;
    rand bit [7:0]   io_commits_info_1_debug_otherPdest_2;
    rand bit [7:0]   io_commits_info_1_debug_otherPdest_3;
    rand bit [7:0]   io_commits_info_1_debug_otherPdest_4;
    rand bit [7:0]   io_commits_info_1_debug_otherPdest_5;
    rand bit [7:0]   io_commits_info_1_debug_otherPdest_6;
    rand bit [34:0]  io_commits_info_1_debug_fuType;
    rand bit         io_commits_info_1_dirtyFs;
    rand bit         io_commits_info_1_dirtyVs;
    rand bit         io_commits_info_2_walk_v;
    rand bit         io_commits_info_2_commit_v;
    rand bit         io_commits_info_2_commit_w;
    rand bit [6:0]   io_commits_info_2_realDestSize;
    rand bit         io_commits_info_2_interrupt_safe;
    rand bit         io_commits_info_2_wflags;
    rand bit [4:0]   io_commits_info_2_fflags;
    rand bit         io_commits_info_2_vxsat;
    rand bit         io_commits_info_2_isRVC;
    rand bit         io_commits_info_2_isVset;
    rand bit         io_commits_info_2_isHls;
    rand bit         io_commits_info_2_isVls;
    rand bit         io_commits_info_2_vls;
    rand bit         io_commits_info_2_mmio;
    rand bit [2:0]   io_commits_info_2_commitType;
    rand bit         io_commits_info_2_ftqIdx_flag;
    rand bit [5:0]   io_commits_info_2_ftqIdx_value;
    rand bit [3:0]   io_commits_info_2_ftqOffset;
    rand bit [2:0]   io_commits_info_2_instrSize;
    rand bit         io_commits_info_2_fpWen;
    rand bit         io_commits_info_2_rfWen;
    rand bit         io_commits_info_2_needFlush;
    rand bit [3:0]   io_commits_info_2_traceBlockInPipe_itype;
    rand bit [3:0]   io_commits_info_2_traceBlockInPipe_iretire;
    rand bit         io_commits_info_2_traceBlockInPipe_ilastsize;
    rand bit [49:0]  io_commits_info_2_debug_pc;
    rand bit [31:0]  io_commits_info_2_debug_instr;
    rand bit [5:0]   io_commits_info_2_debug_ldest;
    rand bit [7:0]   io_commits_info_2_debug_pdest;
    rand bit [7:0]   io_commits_info_2_debug_otherPdest_0;
    rand bit [7:0]   io_commits_info_2_debug_otherPdest_1;
    rand bit [7:0]   io_commits_info_2_debug_otherPdest_2;
    rand bit [7:0]   io_commits_info_2_debug_otherPdest_3;
    rand bit [7:0]   io_commits_info_2_debug_otherPdest_4;
    rand bit [7:0]   io_commits_info_2_debug_otherPdest_5;
    rand bit [7:0]   io_commits_info_2_debug_otherPdest_6;
    rand bit [34:0]  io_commits_info_2_debug_fuType;
    rand bit         io_commits_info_2_dirtyFs;
    rand bit         io_commits_info_2_dirtyVs;
    rand bit         io_commits_info_3_walk_v;
    rand bit         io_commits_info_3_commit_v;
    rand bit         io_commits_info_3_commit_w;
    rand bit [6:0]   io_commits_info_3_realDestSize;
    rand bit         io_commits_info_3_interrupt_safe;
    rand bit         io_commits_info_3_wflags;
    rand bit [4:0]   io_commits_info_3_fflags;
    rand bit         io_commits_info_3_vxsat;
    rand bit         io_commits_info_3_isRVC;
    rand bit         io_commits_info_3_isVset;
    rand bit         io_commits_info_3_isHls;
    rand bit         io_commits_info_3_isVls;
    rand bit         io_commits_info_3_vls;
    rand bit         io_commits_info_3_mmio;
    rand bit [2:0]   io_commits_info_3_commitType;
    rand bit         io_commits_info_3_ftqIdx_flag;
    rand bit [5:0]   io_commits_info_3_ftqIdx_value;
    rand bit [3:0]   io_commits_info_3_ftqOffset;
    rand bit [2:0]   io_commits_info_3_instrSize;
    rand bit         io_commits_info_3_fpWen;
    rand bit         io_commits_info_3_rfWen;
    rand bit         io_commits_info_3_needFlush;
    rand bit [3:0]   io_commits_info_3_traceBlockInPipe_itype;
    rand bit [3:0]   io_commits_info_3_traceBlockInPipe_iretire;
    rand bit         io_commits_info_3_traceBlockInPipe_ilastsize;
    rand bit [49:0]  io_commits_info_3_debug_pc;
    rand bit [31:0]  io_commits_info_3_debug_instr;
    rand bit [5:0]   io_commits_info_3_debug_ldest;
    rand bit [7:0]   io_commits_info_3_debug_pdest;
    rand bit [7:0]   io_commits_info_3_debug_otherPdest_0;
    rand bit [7:0]   io_commits_info_3_debug_otherPdest_1;
    rand bit [7:0]   io_commits_info_3_debug_otherPdest_2;
    rand bit [7:0]   io_commits_info_3_debug_otherPdest_3;
    rand bit [7:0]   io_commits_info_3_debug_otherPdest_4;
    rand bit [7:0]   io_commits_info_3_debug_otherPdest_5;
    rand bit [7:0]   io_commits_info_3_debug_otherPdest_6;
    rand bit [34:0]  io_commits_info_3_debug_fuType;
    rand bit         io_commits_info_3_dirtyFs;
    rand bit         io_commits_info_3_dirtyVs;
    rand bit         io_commits_info_4_walk_v;
    rand bit         io_commits_info_4_commit_v;
    rand bit         io_commits_info_4_commit_w;
    rand bit [6:0]   io_commits_info_4_realDestSize;
    rand bit         io_commits_info_4_interrupt_safe;
    rand bit         io_commits_info_4_wflags;
    rand bit [4:0]   io_commits_info_4_fflags;
    rand bit         io_commits_info_4_vxsat;
    rand bit         io_commits_info_4_isRVC;
    rand bit         io_commits_info_4_isVset;
    rand bit         io_commits_info_4_isHls;
    rand bit         io_commits_info_4_isVls;
    rand bit         io_commits_info_4_vls;
    rand bit         io_commits_info_4_mmio;
    rand bit [2:0]   io_commits_info_4_commitType;
    rand bit         io_commits_info_4_ftqIdx_flag;
    rand bit [5:0]   io_commits_info_4_ftqIdx_value;
    rand bit [3:0]   io_commits_info_4_ftqOffset;
    rand bit [2:0]   io_commits_info_4_instrSize;
    rand bit         io_commits_info_4_fpWen;
    rand bit         io_commits_info_4_rfWen;
    rand bit         io_commits_info_4_needFlush;
    rand bit [3:0]   io_commits_info_4_traceBlockInPipe_itype;
    rand bit [3:0]   io_commits_info_4_traceBlockInPipe_iretire;
    rand bit         io_commits_info_4_traceBlockInPipe_ilastsize;
    rand bit [49:0]  io_commits_info_4_debug_pc;
    rand bit [31:0]  io_commits_info_4_debug_instr;
    rand bit [5:0]   io_commits_info_4_debug_ldest;
    rand bit [7:0]   io_commits_info_4_debug_pdest;
    rand bit [7:0]   io_commits_info_4_debug_otherPdest_0;
    rand bit [7:0]   io_commits_info_4_debug_otherPdest_1;
    rand bit [7:0]   io_commits_info_4_debug_otherPdest_2;
    rand bit [7:0]   io_commits_info_4_debug_otherPdest_3;
    rand bit [7:0]   io_commits_info_4_debug_otherPdest_4;
    rand bit [7:0]   io_commits_info_4_debug_otherPdest_5;
    rand bit [7:0]   io_commits_info_4_debug_otherPdest_6;
    rand bit [34:0]  io_commits_info_4_debug_fuType;
    rand bit         io_commits_info_4_dirtyFs;
    rand bit         io_commits_info_4_dirtyVs;
    rand bit         io_commits_info_5_walk_v;
    rand bit         io_commits_info_5_commit_v;
    rand bit         io_commits_info_5_commit_w;
    rand bit [6:0]   io_commits_info_5_realDestSize;
    rand bit         io_commits_info_5_interrupt_safe;
    rand bit         io_commits_info_5_wflags;
    rand bit [4:0]   io_commits_info_5_fflags;
    rand bit         io_commits_info_5_vxsat;
    rand bit         io_commits_info_5_isRVC;
    rand bit         io_commits_info_5_isVset;
    rand bit         io_commits_info_5_isHls;
    rand bit         io_commits_info_5_isVls;
    rand bit         io_commits_info_5_vls;
    rand bit         io_commits_info_5_mmio;
    rand bit [2:0]   io_commits_info_5_commitType;
    rand bit         io_commits_info_5_ftqIdx_flag;
    rand bit [5:0]   io_commits_info_5_ftqIdx_value;
    rand bit [3:0]   io_commits_info_5_ftqOffset;
    rand bit [2:0]   io_commits_info_5_instrSize;
    rand bit         io_commits_info_5_fpWen;
    rand bit         io_commits_info_5_rfWen;
    rand bit         io_commits_info_5_needFlush;
    rand bit [3:0]   io_commits_info_5_traceBlockInPipe_itype;
    rand bit [3:0]   io_commits_info_5_traceBlockInPipe_iretire;
    rand bit         io_commits_info_5_traceBlockInPipe_ilastsize;
    rand bit [49:0]  io_commits_info_5_debug_pc;
    rand bit [31:0]  io_commits_info_5_debug_instr;
    rand bit [5:0]   io_commits_info_5_debug_ldest;
    rand bit [7:0]   io_commits_info_5_debug_pdest;
    rand bit [7:0]   io_commits_info_5_debug_otherPdest_0;
    rand bit [7:0]   io_commits_info_5_debug_otherPdest_1;
    rand bit [7:0]   io_commits_info_5_debug_otherPdest_2;
    rand bit [7:0]   io_commits_info_5_debug_otherPdest_3;
    rand bit [7:0]   io_commits_info_5_debug_otherPdest_4;
    rand bit [7:0]   io_commits_info_5_debug_otherPdest_5;
    rand bit [7:0]   io_commits_info_5_debug_otherPdest_6;
    rand bit [34:0]  io_commits_info_5_debug_fuType;
    rand bit         io_commits_info_5_dirtyFs;
    rand bit         io_commits_info_5_dirtyVs;
    rand bit         io_commits_info_6_walk_v;
    rand bit         io_commits_info_6_commit_v;
    rand bit         io_commits_info_6_commit_w;
    rand bit [6:0]   io_commits_info_6_realDestSize;
    rand bit         io_commits_info_6_interrupt_safe;
    rand bit         io_commits_info_6_wflags;
    rand bit [4:0]   io_commits_info_6_fflags;
    rand bit         io_commits_info_6_vxsat;
    rand bit         io_commits_info_6_isRVC;
    rand bit         io_commits_info_6_isVset;
    rand bit         io_commits_info_6_isHls;
    rand bit         io_commits_info_6_isVls;
    rand bit         io_commits_info_6_vls;
    rand bit         io_commits_info_6_mmio;
    rand bit [2:0]   io_commits_info_6_commitType;
    rand bit         io_commits_info_6_ftqIdx_flag;
    rand bit [5:0]   io_commits_info_6_ftqIdx_value;
    rand bit [3:0]   io_commits_info_6_ftqOffset;
    rand bit [2:0]   io_commits_info_6_instrSize;
    rand bit         io_commits_info_6_fpWen;
    rand bit         io_commits_info_6_rfWen;
    rand bit         io_commits_info_6_needFlush;
    rand bit [3:0]   io_commits_info_6_traceBlockInPipe_itype;
    rand bit [3:0]   io_commits_info_6_traceBlockInPipe_iretire;
    rand bit         io_commits_info_6_traceBlockInPipe_ilastsize;
    rand bit [49:0]  io_commits_info_6_debug_pc;
    rand bit [31:0]  io_commits_info_6_debug_instr;
    rand bit [5:0]   io_commits_info_6_debug_ldest;
    rand bit [7:0]   io_commits_info_6_debug_pdest;
    rand bit [7:0]   io_commits_info_6_debug_otherPdest_0;
    rand bit [7:0]   io_commits_info_6_debug_otherPdest_1;
    rand bit [7:0]   io_commits_info_6_debug_otherPdest_2;
    rand bit [7:0]   io_commits_info_6_debug_otherPdest_3;
    rand bit [7:0]   io_commits_info_6_debug_otherPdest_4;
    rand bit [7:0]   io_commits_info_6_debug_otherPdest_5;
    rand bit [7:0]   io_commits_info_6_debug_otherPdest_6;
    rand bit [34:0]  io_commits_info_6_debug_fuType;
    rand bit         io_commits_info_6_dirtyFs;
    rand bit         io_commits_info_6_dirtyVs;
    rand bit         io_commits_info_7_walk_v;
    rand bit         io_commits_info_7_commit_v;
    rand bit         io_commits_info_7_commit_w;
    rand bit [6:0]   io_commits_info_7_realDestSize;
    rand bit         io_commits_info_7_interrupt_safe;
    rand bit         io_commits_info_7_wflags;
    rand bit [4:0]   io_commits_info_7_fflags;
    rand bit         io_commits_info_7_vxsat;
    rand bit         io_commits_info_7_isRVC;
    rand bit         io_commits_info_7_isVset;
    rand bit         io_commits_info_7_isHls;
    rand bit         io_commits_info_7_isVls;
    rand bit         io_commits_info_7_vls;
    rand bit         io_commits_info_7_mmio;
    rand bit [2:0]   io_commits_info_7_commitType;
    rand bit         io_commits_info_7_ftqIdx_flag;
    rand bit [5:0]   io_commits_info_7_ftqIdx_value;
    rand bit [3:0]   io_commits_info_7_ftqOffset;
    rand bit [2:0]   io_commits_info_7_instrSize;
    rand bit         io_commits_info_7_fpWen;
    rand bit         io_commits_info_7_rfWen;
    rand bit         io_commits_info_7_needFlush;
    rand bit [3:0]   io_commits_info_7_traceBlockInPipe_itype;
    rand bit [3:0]   io_commits_info_7_traceBlockInPipe_iretire;
    rand bit         io_commits_info_7_traceBlockInPipe_ilastsize;
    rand bit [49:0]  io_commits_info_7_debug_pc;
    rand bit [31:0]  io_commits_info_7_debug_instr;
    rand bit [5:0]   io_commits_info_7_debug_ldest;
    rand bit [7:0]   io_commits_info_7_debug_pdest;
    rand bit [7:0]   io_commits_info_7_debug_otherPdest_0;
    rand bit [7:0]   io_commits_info_7_debug_otherPdest_1;
    rand bit [7:0]   io_commits_info_7_debug_otherPdest_2;
    rand bit [7:0]   io_commits_info_7_debug_otherPdest_3;
    rand bit [7:0]   io_commits_info_7_debug_otherPdest_4;
    rand bit [7:0]   io_commits_info_7_debug_otherPdest_5;
    rand bit [7:0]   io_commits_info_7_debug_otherPdest_6;
    rand bit [34:0]  io_commits_info_7_debug_fuType;
    rand bit         io_commits_info_7_dirtyFs;
    rand bit         io_commits_info_7_dirtyVs;
    rand bit         io_commits_robIdx_0_flag;
    rand bit [7:0]   io_commits_robIdx_0_value;
    rand bit         io_commits_robIdx_1_flag;
    rand bit [7:0]   io_commits_robIdx_1_value;
    rand bit         io_commits_robIdx_2_flag;
    rand bit [7:0]   io_commits_robIdx_2_value;
    rand bit         io_commits_robIdx_3_flag;
    rand bit [7:0]   io_commits_robIdx_3_value;
    rand bit         io_commits_robIdx_4_flag;
    rand bit [7:0]   io_commits_robIdx_4_value;
    rand bit         io_commits_robIdx_5_flag;
    rand bit [7:0]   io_commits_robIdx_5_value;
    rand bit         io_commits_robIdx_6_flag;
    rand bit [7:0]   io_commits_robIdx_6_value;
    rand bit         io_commits_robIdx_7_flag;
    rand bit [7:0]   io_commits_robIdx_7_value;
    rand bit         io_trace_blockCommit;
    rand bit         io_trace_traceCommitInfo_blocks_0_valid;
    rand bit [5:0]   io_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value;
    rand bit [3:0]   io_trace_traceCommitInfo_blocks_0_bits_ftqOffset;
    rand bit [3:0]   io_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype;
    rand bit [3:0]   io_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire;
    rand bit         io_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize;
    rand bit         io_trace_traceCommitInfo_blocks_1_valid;
    rand bit [5:0]   io_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value;
    rand bit [3:0]   io_trace_traceCommitInfo_blocks_1_bits_ftqOffset;
    rand bit [3:0]   io_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype;
    rand bit [3:0]   io_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire;
    rand bit         io_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize;
    rand bit         io_trace_traceCommitInfo_blocks_2_valid;
    rand bit [5:0]   io_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value;
    rand bit [3:0]   io_trace_traceCommitInfo_blocks_2_bits_ftqOffset;
    rand bit [3:0]   io_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype;
    rand bit [3:0]   io_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire;
    rand bit         io_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize;
    rand bit         io_trace_traceCommitInfo_blocks_3_valid;
    rand bit [5:0]   io_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value;
    rand bit [3:0]   io_trace_traceCommitInfo_blocks_3_bits_ftqOffset;
    rand bit [3:0]   io_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype;
    rand bit [3:0]   io_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire;
    rand bit         io_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize;
    rand bit         io_trace_traceCommitInfo_blocks_4_valid;
    rand bit [5:0]   io_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value;
    rand bit [3:0]   io_trace_traceCommitInfo_blocks_4_bits_ftqOffset;
    rand bit [3:0]   io_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype;
    rand bit [3:0]   io_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire;
    rand bit         io_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize;
    rand bit         io_trace_traceCommitInfo_blocks_5_valid;
    rand bit [5:0]   io_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value;
    rand bit [3:0]   io_trace_traceCommitInfo_blocks_5_bits_ftqOffset;
    rand bit [3:0]   io_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype;
    rand bit [3:0]   io_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire;
    rand bit         io_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize;
    rand bit         io_trace_traceCommitInfo_blocks_6_valid;
    rand bit [5:0]   io_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value;
    rand bit [3:0]   io_trace_traceCommitInfo_blocks_6_bits_ftqOffset;
    rand bit [3:0]   io_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype;
    rand bit [3:0]   io_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire;
    rand bit         io_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize;
    rand bit         io_trace_traceCommitInfo_blocks_7_valid;
    rand bit [5:0]   io_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value;
    rand bit [3:0]   io_trace_traceCommitInfo_blocks_7_bits_ftqOffset;
    rand bit [3:0]   io_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype;
    rand bit [3:0]   io_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire;
    rand bit         io_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize;
    rand bit         io_rabCommits_isCommit;
    rand bit         io_rabCommits_commitValid_0;
    rand bit         io_rabCommits_commitValid_1;
    rand bit         io_rabCommits_commitValid_2;
    rand bit         io_rabCommits_commitValid_3;
    rand bit         io_rabCommits_commitValid_4;
    rand bit         io_rabCommits_commitValid_5;
    rand bit         io_rabCommits_isWalk;
    rand bit         io_rabCommits_walkValid_0;
    rand bit         io_rabCommits_walkValid_1;
    rand bit         io_rabCommits_walkValid_2;
    rand bit         io_rabCommits_walkValid_3;
    rand bit         io_rabCommits_walkValid_4;
    rand bit         io_rabCommits_walkValid_5;
    rand bit [5:0]   io_rabCommits_info_0_ldest;
    rand bit [7:0]   io_rabCommits_info_0_pdest;
    rand bit         io_rabCommits_info_0_rfWen;
    rand bit         io_rabCommits_info_0_fpWen;
    rand bit         io_rabCommits_info_0_vecWen;
    rand bit         io_rabCommits_info_0_v0Wen;
    rand bit         io_rabCommits_info_0_vlWen;
    rand bit         io_rabCommits_info_0_isMove;
    rand bit [5:0]   io_rabCommits_info_1_ldest;
    rand bit [7:0]   io_rabCommits_info_1_pdest;
    rand bit         io_rabCommits_info_1_rfWen;
    rand bit         io_rabCommits_info_1_fpWen;
    rand bit         io_rabCommits_info_1_vecWen;
    rand bit         io_rabCommits_info_1_v0Wen;
    rand bit         io_rabCommits_info_1_vlWen;
    rand bit         io_rabCommits_info_1_isMove;
    rand bit [5:0]   io_rabCommits_info_2_ldest;
    rand bit [7:0]   io_rabCommits_info_2_pdest;
    rand bit         io_rabCommits_info_2_rfWen;
    rand bit         io_rabCommits_info_2_fpWen;
    rand bit         io_rabCommits_info_2_vecWen;
    rand bit         io_rabCommits_info_2_v0Wen;
    rand bit         io_rabCommits_info_2_vlWen;
    rand bit         io_rabCommits_info_2_isMove;
    rand bit [5:0]   io_rabCommits_info_3_ldest;
    rand bit [7:0]   io_rabCommits_info_3_pdest;
    rand bit         io_rabCommits_info_3_rfWen;
    rand bit         io_rabCommits_info_3_fpWen;
    rand bit         io_rabCommits_info_3_vecWen;
    rand bit         io_rabCommits_info_3_v0Wen;
    rand bit         io_rabCommits_info_3_vlWen;
    rand bit         io_rabCommits_info_3_isMove;
    rand bit [5:0]   io_rabCommits_info_4_ldest;
    rand bit [7:0]   io_rabCommits_info_4_pdest;
    rand bit         io_rabCommits_info_4_rfWen;
    rand bit         io_rabCommits_info_4_fpWen;
    rand bit         io_rabCommits_info_4_vecWen;
    rand bit         io_rabCommits_info_4_v0Wen;
    rand bit         io_rabCommits_info_4_vlWen;
    rand bit         io_rabCommits_info_4_isMove;
    rand bit [5:0]   io_rabCommits_info_5_ldest;
    rand bit [7:0]   io_rabCommits_info_5_pdest;
    rand bit         io_rabCommits_info_5_rfWen;
    rand bit         io_rabCommits_info_5_fpWen;
    rand bit         io_rabCommits_info_5_vecWen;
    rand bit         io_rabCommits_info_5_v0Wen;
    rand bit         io_rabCommits_info_5_vlWen;
    rand bit         io_rabCommits_info_5_isMove;
    rand bit         io_diffCommits_commitValid_0;
    rand bit         io_diffCommits_commitValid_1;
    rand bit         io_diffCommits_commitValid_2;
    rand bit         io_diffCommits_commitValid_3;
    rand bit         io_diffCommits_commitValid_4;
    rand bit         io_diffCommits_commitValid_5;
    rand bit         io_diffCommits_commitValid_6;
    rand bit         io_diffCommits_commitValid_7;
    rand bit         io_diffCommits_commitValid_8;
    rand bit         io_diffCommits_commitValid_9;
    rand bit         io_diffCommits_commitValid_10;
    rand bit         io_diffCommits_commitValid_11;
    rand bit         io_diffCommits_commitValid_12;
    rand bit         io_diffCommits_commitValid_13;
    rand bit         io_diffCommits_commitValid_14;
    rand bit         io_diffCommits_commitValid_15;
    rand bit         io_diffCommits_commitValid_16;
    rand bit         io_diffCommits_commitValid_17;
    rand bit         io_diffCommits_commitValid_18;
    rand bit         io_diffCommits_commitValid_19;
    rand bit         io_diffCommits_commitValid_20;
    rand bit         io_diffCommits_commitValid_21;
    rand bit         io_diffCommits_commitValid_22;
    rand bit         io_diffCommits_commitValid_23;
    rand bit         io_diffCommits_commitValid_24;
    rand bit         io_diffCommits_commitValid_25;
    rand bit         io_diffCommits_commitValid_26;
    rand bit         io_diffCommits_commitValid_27;
    rand bit         io_diffCommits_commitValid_28;
    rand bit         io_diffCommits_commitValid_29;
    rand bit         io_diffCommits_commitValid_30;
    rand bit         io_diffCommits_commitValid_31;
    rand bit         io_diffCommits_commitValid_32;
    rand bit         io_diffCommits_commitValid_33;
    rand bit         io_diffCommits_commitValid_34;
    rand bit         io_diffCommits_commitValid_35;
    rand bit         io_diffCommits_commitValid_36;
    rand bit         io_diffCommits_commitValid_37;
    rand bit         io_diffCommits_commitValid_38;
    rand bit         io_diffCommits_commitValid_39;
    rand bit         io_diffCommits_commitValid_40;
    rand bit         io_diffCommits_commitValid_41;
    rand bit         io_diffCommits_commitValid_42;
    rand bit         io_diffCommits_commitValid_43;
    rand bit         io_diffCommits_commitValid_44;
    rand bit         io_diffCommits_commitValid_45;
    rand bit         io_diffCommits_commitValid_46;
    rand bit         io_diffCommits_commitValid_47;
    rand bit         io_diffCommits_commitValid_48;
    rand bit         io_diffCommits_commitValid_49;
    rand bit         io_diffCommits_commitValid_50;
    rand bit         io_diffCommits_commitValid_51;
    rand bit         io_diffCommits_commitValid_52;
    rand bit         io_diffCommits_commitValid_53;
    rand bit         io_diffCommits_commitValid_54;
    rand bit         io_diffCommits_commitValid_55;
    rand bit         io_diffCommits_commitValid_56;
    rand bit         io_diffCommits_commitValid_57;
    rand bit         io_diffCommits_commitValid_58;
    rand bit         io_diffCommits_commitValid_59;
    rand bit         io_diffCommits_commitValid_60;
    rand bit         io_diffCommits_commitValid_61;
    rand bit         io_diffCommits_commitValid_62;
    rand bit         io_diffCommits_commitValid_63;
    rand bit         io_diffCommits_commitValid_64;
    rand bit         io_diffCommits_commitValid_65;
    rand bit         io_diffCommits_commitValid_66;
    rand bit         io_diffCommits_commitValid_67;
    rand bit         io_diffCommits_commitValid_68;
    rand bit         io_diffCommits_commitValid_69;
    rand bit         io_diffCommits_commitValid_70;
    rand bit         io_diffCommits_commitValid_71;
    rand bit         io_diffCommits_commitValid_72;
    rand bit         io_diffCommits_commitValid_73;
    rand bit         io_diffCommits_commitValid_74;
    rand bit         io_diffCommits_commitValid_75;
    rand bit         io_diffCommits_commitValid_76;
    rand bit         io_diffCommits_commitValid_77;
    rand bit         io_diffCommits_commitValid_78;
    rand bit         io_diffCommits_commitValid_79;
    rand bit         io_diffCommits_commitValid_80;
    rand bit         io_diffCommits_commitValid_81;
    rand bit         io_diffCommits_commitValid_82;
    rand bit         io_diffCommits_commitValid_83;
    rand bit         io_diffCommits_commitValid_84;
    rand bit         io_diffCommits_commitValid_85;
    rand bit         io_diffCommits_commitValid_86;
    rand bit         io_diffCommits_commitValid_87;
    rand bit         io_diffCommits_commitValid_88;
    rand bit         io_diffCommits_commitValid_89;
    rand bit         io_diffCommits_commitValid_90;
    rand bit         io_diffCommits_commitValid_91;
    rand bit         io_diffCommits_commitValid_92;
    rand bit         io_diffCommits_commitValid_93;
    rand bit         io_diffCommits_commitValid_94;
    rand bit         io_diffCommits_commitValid_95;
    rand bit         io_diffCommits_commitValid_96;
    rand bit         io_diffCommits_commitValid_97;
    rand bit         io_diffCommits_commitValid_98;
    rand bit         io_diffCommits_commitValid_99;
    rand bit         io_diffCommits_commitValid_100;
    rand bit         io_diffCommits_commitValid_101;
    rand bit         io_diffCommits_commitValid_102;
    rand bit         io_diffCommits_commitValid_103;
    rand bit         io_diffCommits_commitValid_104;
    rand bit         io_diffCommits_commitValid_105;
    rand bit         io_diffCommits_commitValid_106;
    rand bit         io_diffCommits_commitValid_107;
    rand bit         io_diffCommits_commitValid_108;
    rand bit         io_diffCommits_commitValid_109;
    rand bit         io_diffCommits_commitValid_110;
    rand bit         io_diffCommits_commitValid_111;
    rand bit         io_diffCommits_commitValid_112;
    rand bit         io_diffCommits_commitValid_113;
    rand bit         io_diffCommits_commitValid_114;
    rand bit         io_diffCommits_commitValid_115;
    rand bit         io_diffCommits_commitValid_116;
    rand bit         io_diffCommits_commitValid_117;
    rand bit         io_diffCommits_commitValid_118;
    rand bit         io_diffCommits_commitValid_119;
    rand bit         io_diffCommits_commitValid_120;
    rand bit         io_diffCommits_commitValid_121;
    rand bit         io_diffCommits_commitValid_122;
    rand bit         io_diffCommits_commitValid_123;
    rand bit         io_diffCommits_commitValid_124;
    rand bit         io_diffCommits_commitValid_125;
    rand bit         io_diffCommits_commitValid_126;
    rand bit         io_diffCommits_commitValid_127;
    rand bit         io_diffCommits_commitValid_128;
    rand bit         io_diffCommits_commitValid_129;
    rand bit         io_diffCommits_commitValid_130;
    rand bit         io_diffCommits_commitValid_131;
    rand bit         io_diffCommits_commitValid_132;
    rand bit         io_diffCommits_commitValid_133;
    rand bit         io_diffCommits_commitValid_134;
    rand bit         io_diffCommits_commitValid_135;
    rand bit         io_diffCommits_commitValid_136;
    rand bit         io_diffCommits_commitValid_137;
    rand bit         io_diffCommits_commitValid_138;
    rand bit         io_diffCommits_commitValid_139;
    rand bit         io_diffCommits_commitValid_140;
    rand bit         io_diffCommits_commitValid_141;
    rand bit         io_diffCommits_commitValid_142;
    rand bit         io_diffCommits_commitValid_143;
    rand bit         io_diffCommits_commitValid_144;
    rand bit         io_diffCommits_commitValid_145;
    rand bit         io_diffCommits_commitValid_146;
    rand bit         io_diffCommits_commitValid_147;
    rand bit         io_diffCommits_commitValid_148;
    rand bit         io_diffCommits_commitValid_149;
    rand bit         io_diffCommits_commitValid_150;
    rand bit         io_diffCommits_commitValid_151;
    rand bit         io_diffCommits_commitValid_152;
    rand bit         io_diffCommits_commitValid_153;
    rand bit         io_diffCommits_commitValid_154;
    rand bit         io_diffCommits_commitValid_155;
    rand bit         io_diffCommits_commitValid_156;
    rand bit         io_diffCommits_commitValid_157;
    rand bit         io_diffCommits_commitValid_158;
    rand bit         io_diffCommits_commitValid_159;
    rand bit         io_diffCommits_commitValid_160;
    rand bit         io_diffCommits_commitValid_161;
    rand bit         io_diffCommits_commitValid_162;
    rand bit         io_diffCommits_commitValid_163;
    rand bit         io_diffCommits_commitValid_164;
    rand bit         io_diffCommits_commitValid_165;
    rand bit         io_diffCommits_commitValid_166;
    rand bit         io_diffCommits_commitValid_167;
    rand bit         io_diffCommits_commitValid_168;
    rand bit         io_diffCommits_commitValid_169;
    rand bit         io_diffCommits_commitValid_170;
    rand bit         io_diffCommits_commitValid_171;
    rand bit         io_diffCommits_commitValid_172;
    rand bit         io_diffCommits_commitValid_173;
    rand bit         io_diffCommits_commitValid_174;
    rand bit         io_diffCommits_commitValid_175;
    rand bit         io_diffCommits_commitValid_176;
    rand bit         io_diffCommits_commitValid_177;
    rand bit         io_diffCommits_commitValid_178;
    rand bit         io_diffCommits_commitValid_179;
    rand bit         io_diffCommits_commitValid_180;
    rand bit         io_diffCommits_commitValid_181;
    rand bit         io_diffCommits_commitValid_182;
    rand bit         io_diffCommits_commitValid_183;
    rand bit         io_diffCommits_commitValid_184;
    rand bit         io_diffCommits_commitValid_185;
    rand bit         io_diffCommits_commitValid_186;
    rand bit         io_diffCommits_commitValid_187;
    rand bit         io_diffCommits_commitValid_188;
    rand bit         io_diffCommits_commitValid_189;
    rand bit         io_diffCommits_commitValid_190;
    rand bit         io_diffCommits_commitValid_191;
    rand bit         io_diffCommits_commitValid_192;
    rand bit         io_diffCommits_commitValid_193;
    rand bit         io_diffCommits_commitValid_194;
    rand bit         io_diffCommits_commitValid_195;
    rand bit         io_diffCommits_commitValid_196;
    rand bit         io_diffCommits_commitValid_197;
    rand bit         io_diffCommits_commitValid_198;
    rand bit         io_diffCommits_commitValid_199;
    rand bit         io_diffCommits_commitValid_200;
    rand bit         io_diffCommits_commitValid_201;
    rand bit         io_diffCommits_commitValid_202;
    rand bit         io_diffCommits_commitValid_203;
    rand bit         io_diffCommits_commitValid_204;
    rand bit         io_diffCommits_commitValid_205;
    rand bit         io_diffCommits_commitValid_206;
    rand bit         io_diffCommits_commitValid_207;
    rand bit         io_diffCommits_commitValid_208;
    rand bit         io_diffCommits_commitValid_209;
    rand bit         io_diffCommits_commitValid_210;
    rand bit         io_diffCommits_commitValid_211;
    rand bit         io_diffCommits_commitValid_212;
    rand bit         io_diffCommits_commitValid_213;
    rand bit         io_diffCommits_commitValid_214;
    rand bit         io_diffCommits_commitValid_215;
    rand bit         io_diffCommits_commitValid_216;
    rand bit         io_diffCommits_commitValid_217;
    rand bit         io_diffCommits_commitValid_218;
    rand bit         io_diffCommits_commitValid_219;
    rand bit         io_diffCommits_commitValid_220;
    rand bit         io_diffCommits_commitValid_221;
    rand bit         io_diffCommits_commitValid_222;
    rand bit         io_diffCommits_commitValid_223;
    rand bit         io_diffCommits_commitValid_224;
    rand bit         io_diffCommits_commitValid_225;
    rand bit         io_diffCommits_commitValid_226;
    rand bit         io_diffCommits_commitValid_227;
    rand bit         io_diffCommits_commitValid_228;
    rand bit         io_diffCommits_commitValid_229;
    rand bit         io_diffCommits_commitValid_230;
    rand bit         io_diffCommits_commitValid_231;
    rand bit         io_diffCommits_commitValid_232;
    rand bit         io_diffCommits_commitValid_233;
    rand bit         io_diffCommits_commitValid_234;
    rand bit         io_diffCommits_commitValid_235;
    rand bit         io_diffCommits_commitValid_236;
    rand bit         io_diffCommits_commitValid_237;
    rand bit         io_diffCommits_commitValid_238;
    rand bit         io_diffCommits_commitValid_239;
    rand bit         io_diffCommits_commitValid_240;
    rand bit         io_diffCommits_commitValid_241;
    rand bit         io_diffCommits_commitValid_242;
    rand bit         io_diffCommits_commitValid_243;
    rand bit         io_diffCommits_commitValid_244;
    rand bit         io_diffCommits_commitValid_245;
    rand bit         io_diffCommits_commitValid_246;
    rand bit         io_diffCommits_commitValid_247;
    rand bit         io_diffCommits_commitValid_248;
    rand bit         io_diffCommits_commitValid_249;
    rand bit         io_diffCommits_commitValid_250;
    rand bit         io_diffCommits_commitValid_251;
    rand bit         io_diffCommits_commitValid_252;
    rand bit         io_diffCommits_commitValid_253;
    rand bit         io_diffCommits_commitValid_254;
    rand bit [5:0]   io_diffCommits_info_0_ldest;
    rand bit [7:0]   io_diffCommits_info_0_pdest;
    rand bit         io_diffCommits_info_0_rfWen;
    rand bit         io_diffCommits_info_0_fpWen;
    rand bit         io_diffCommits_info_0_vecWen;
    rand bit         io_diffCommits_info_0_v0Wen;
    rand bit         io_diffCommits_info_0_vlWen;
    rand bit [5:0]   io_diffCommits_info_1_ldest;
    rand bit [7:0]   io_diffCommits_info_1_pdest;
    rand bit         io_diffCommits_info_1_rfWen;
    rand bit         io_diffCommits_info_1_fpWen;
    rand bit         io_diffCommits_info_1_vecWen;
    rand bit         io_diffCommits_info_1_v0Wen;
    rand bit         io_diffCommits_info_1_vlWen;
    rand bit [5:0]   io_diffCommits_info_2_ldest;
    rand bit [7:0]   io_diffCommits_info_2_pdest;
    rand bit         io_diffCommits_info_2_rfWen;
    rand bit         io_diffCommits_info_2_fpWen;
    rand bit         io_diffCommits_info_2_vecWen;
    rand bit         io_diffCommits_info_2_v0Wen;
    rand bit         io_diffCommits_info_2_vlWen;
    rand bit [5:0]   io_diffCommits_info_3_ldest;
    rand bit [7:0]   io_diffCommits_info_3_pdest;
    rand bit         io_diffCommits_info_3_rfWen;
    rand bit         io_diffCommits_info_3_fpWen;
    rand bit         io_diffCommits_info_3_vecWen;
    rand bit         io_diffCommits_info_3_v0Wen;
    rand bit         io_diffCommits_info_3_vlWen;
    rand bit [5:0]   io_diffCommits_info_4_ldest;
    rand bit [7:0]   io_diffCommits_info_4_pdest;
    rand bit         io_diffCommits_info_4_rfWen;
    rand bit         io_diffCommits_info_4_fpWen;
    rand bit         io_diffCommits_info_4_vecWen;
    rand bit         io_diffCommits_info_4_v0Wen;
    rand bit         io_diffCommits_info_4_vlWen;
    rand bit [5:0]   io_diffCommits_info_5_ldest;
    rand bit [7:0]   io_diffCommits_info_5_pdest;
    rand bit         io_diffCommits_info_5_rfWen;
    rand bit         io_diffCommits_info_5_fpWen;
    rand bit         io_diffCommits_info_5_vecWen;
    rand bit         io_diffCommits_info_5_v0Wen;
    rand bit         io_diffCommits_info_5_vlWen;
    rand bit [5:0]   io_diffCommits_info_6_ldest;
    rand bit [7:0]   io_diffCommits_info_6_pdest;
    rand bit         io_diffCommits_info_6_rfWen;
    rand bit         io_diffCommits_info_6_fpWen;
    rand bit         io_diffCommits_info_6_vecWen;
    rand bit         io_diffCommits_info_6_v0Wen;
    rand bit         io_diffCommits_info_6_vlWen;
    rand bit [5:0]   io_diffCommits_info_7_ldest;
    rand bit [7:0]   io_diffCommits_info_7_pdest;
    rand bit         io_diffCommits_info_7_rfWen;
    rand bit         io_diffCommits_info_7_fpWen;
    rand bit         io_diffCommits_info_7_vecWen;
    rand bit         io_diffCommits_info_7_v0Wen;
    rand bit         io_diffCommits_info_7_vlWen;
    rand bit [5:0]   io_diffCommits_info_8_ldest;
    rand bit [7:0]   io_diffCommits_info_8_pdest;
    rand bit         io_diffCommits_info_8_rfWen;
    rand bit         io_diffCommits_info_8_fpWen;
    rand bit         io_diffCommits_info_8_vecWen;
    rand bit         io_diffCommits_info_8_v0Wen;
    rand bit         io_diffCommits_info_8_vlWen;
    rand bit [5:0]   io_diffCommits_info_9_ldest;
    rand bit [7:0]   io_diffCommits_info_9_pdest;
    rand bit         io_diffCommits_info_9_rfWen;
    rand bit         io_diffCommits_info_9_fpWen;
    rand bit         io_diffCommits_info_9_vecWen;
    rand bit         io_diffCommits_info_9_v0Wen;
    rand bit         io_diffCommits_info_9_vlWen;
    rand bit [5:0]   io_diffCommits_info_10_ldest;
    rand bit [7:0]   io_diffCommits_info_10_pdest;
    rand bit         io_diffCommits_info_10_rfWen;
    rand bit         io_diffCommits_info_10_fpWen;
    rand bit         io_diffCommits_info_10_vecWen;
    rand bit         io_diffCommits_info_10_v0Wen;
    rand bit         io_diffCommits_info_10_vlWen;
    rand bit [5:0]   io_diffCommits_info_11_ldest;
    rand bit [7:0]   io_diffCommits_info_11_pdest;
    rand bit         io_diffCommits_info_11_rfWen;
    rand bit         io_diffCommits_info_11_fpWen;
    rand bit         io_diffCommits_info_11_vecWen;
    rand bit         io_diffCommits_info_11_v0Wen;
    rand bit         io_diffCommits_info_11_vlWen;
    rand bit [5:0]   io_diffCommits_info_12_ldest;
    rand bit [7:0]   io_diffCommits_info_12_pdest;
    rand bit         io_diffCommits_info_12_rfWen;
    rand bit         io_diffCommits_info_12_fpWen;
    rand bit         io_diffCommits_info_12_vecWen;
    rand bit         io_diffCommits_info_12_v0Wen;
    rand bit         io_diffCommits_info_12_vlWen;
    rand bit [5:0]   io_diffCommits_info_13_ldest;
    rand bit [7:0]   io_diffCommits_info_13_pdest;
    rand bit         io_diffCommits_info_13_rfWen;
    rand bit         io_diffCommits_info_13_fpWen;
    rand bit         io_diffCommits_info_13_vecWen;
    rand bit         io_diffCommits_info_13_v0Wen;
    rand bit         io_diffCommits_info_13_vlWen;
    rand bit [5:0]   io_diffCommits_info_14_ldest;
    rand bit [7:0]   io_diffCommits_info_14_pdest;
    rand bit         io_diffCommits_info_14_rfWen;
    rand bit         io_diffCommits_info_14_fpWen;
    rand bit         io_diffCommits_info_14_vecWen;
    rand bit         io_diffCommits_info_14_v0Wen;
    rand bit         io_diffCommits_info_14_vlWen;
    rand bit [5:0]   io_diffCommits_info_15_ldest;
    rand bit [7:0]   io_diffCommits_info_15_pdest;
    rand bit         io_diffCommits_info_15_rfWen;
    rand bit         io_diffCommits_info_15_fpWen;
    rand bit         io_diffCommits_info_15_vecWen;
    rand bit         io_diffCommits_info_15_v0Wen;
    rand bit         io_diffCommits_info_15_vlWen;
    rand bit [5:0]   io_diffCommits_info_16_ldest;
    rand bit [7:0]   io_diffCommits_info_16_pdest;
    rand bit         io_diffCommits_info_16_rfWen;
    rand bit         io_diffCommits_info_16_fpWen;
    rand bit         io_diffCommits_info_16_vecWen;
    rand bit         io_diffCommits_info_16_v0Wen;
    rand bit         io_diffCommits_info_16_vlWen;
    rand bit [5:0]   io_diffCommits_info_17_ldest;
    rand bit [7:0]   io_diffCommits_info_17_pdest;
    rand bit         io_diffCommits_info_17_rfWen;
    rand bit         io_diffCommits_info_17_fpWen;
    rand bit         io_diffCommits_info_17_vecWen;
    rand bit         io_diffCommits_info_17_v0Wen;
    rand bit         io_diffCommits_info_17_vlWen;
    rand bit [5:0]   io_diffCommits_info_18_ldest;
    rand bit [7:0]   io_diffCommits_info_18_pdest;
    rand bit         io_diffCommits_info_18_rfWen;
    rand bit         io_diffCommits_info_18_fpWen;
    rand bit         io_diffCommits_info_18_vecWen;
    rand bit         io_diffCommits_info_18_v0Wen;
    rand bit         io_diffCommits_info_18_vlWen;
    rand bit [5:0]   io_diffCommits_info_19_ldest;
    rand bit [7:0]   io_diffCommits_info_19_pdest;
    rand bit         io_diffCommits_info_19_rfWen;
    rand bit         io_diffCommits_info_19_fpWen;
    rand bit         io_diffCommits_info_19_vecWen;
    rand bit         io_diffCommits_info_19_v0Wen;
    rand bit         io_diffCommits_info_19_vlWen;
    rand bit [5:0]   io_diffCommits_info_20_ldest;
    rand bit [7:0]   io_diffCommits_info_20_pdest;
    rand bit         io_diffCommits_info_20_rfWen;
    rand bit         io_diffCommits_info_20_fpWen;
    rand bit         io_diffCommits_info_20_vecWen;
    rand bit         io_diffCommits_info_20_v0Wen;
    rand bit         io_diffCommits_info_20_vlWen;
    rand bit [5:0]   io_diffCommits_info_21_ldest;
    rand bit [7:0]   io_diffCommits_info_21_pdest;
    rand bit         io_diffCommits_info_21_rfWen;
    rand bit         io_diffCommits_info_21_fpWen;
    rand bit         io_diffCommits_info_21_vecWen;
    rand bit         io_diffCommits_info_21_v0Wen;
    rand bit         io_diffCommits_info_21_vlWen;
    rand bit [5:0]   io_diffCommits_info_22_ldest;
    rand bit [7:0]   io_diffCommits_info_22_pdest;
    rand bit         io_diffCommits_info_22_rfWen;
    rand bit         io_diffCommits_info_22_fpWen;
    rand bit         io_diffCommits_info_22_vecWen;
    rand bit         io_diffCommits_info_22_v0Wen;
    rand bit         io_diffCommits_info_22_vlWen;
    rand bit [5:0]   io_diffCommits_info_23_ldest;
    rand bit [7:0]   io_diffCommits_info_23_pdest;
    rand bit         io_diffCommits_info_23_rfWen;
    rand bit         io_diffCommits_info_23_fpWen;
    rand bit         io_diffCommits_info_23_vecWen;
    rand bit         io_diffCommits_info_23_v0Wen;
    rand bit         io_diffCommits_info_23_vlWen;
    rand bit [5:0]   io_diffCommits_info_24_ldest;
    rand bit [7:0]   io_diffCommits_info_24_pdest;
    rand bit         io_diffCommits_info_24_rfWen;
    rand bit         io_diffCommits_info_24_fpWen;
    rand bit         io_diffCommits_info_24_vecWen;
    rand bit         io_diffCommits_info_24_v0Wen;
    rand bit         io_diffCommits_info_24_vlWen;
    rand bit [5:0]   io_diffCommits_info_25_ldest;
    rand bit [7:0]   io_diffCommits_info_25_pdest;
    rand bit         io_diffCommits_info_25_rfWen;
    rand bit         io_diffCommits_info_25_fpWen;
    rand bit         io_diffCommits_info_25_vecWen;
    rand bit         io_diffCommits_info_25_v0Wen;
    rand bit         io_diffCommits_info_25_vlWen;
    rand bit [5:0]   io_diffCommits_info_26_ldest;
    rand bit [7:0]   io_diffCommits_info_26_pdest;
    rand bit         io_diffCommits_info_26_rfWen;
    rand bit         io_diffCommits_info_26_fpWen;
    rand bit         io_diffCommits_info_26_vecWen;
    rand bit         io_diffCommits_info_26_v0Wen;
    rand bit         io_diffCommits_info_26_vlWen;
    rand bit [5:0]   io_diffCommits_info_27_ldest;
    rand bit [7:0]   io_diffCommits_info_27_pdest;
    rand bit         io_diffCommits_info_27_rfWen;
    rand bit         io_diffCommits_info_27_fpWen;
    rand bit         io_diffCommits_info_27_vecWen;
    rand bit         io_diffCommits_info_27_v0Wen;
    rand bit         io_diffCommits_info_27_vlWen;
    rand bit [5:0]   io_diffCommits_info_28_ldest;
    rand bit [7:0]   io_diffCommits_info_28_pdest;
    rand bit         io_diffCommits_info_28_rfWen;
    rand bit         io_diffCommits_info_28_fpWen;
    rand bit         io_diffCommits_info_28_vecWen;
    rand bit         io_diffCommits_info_28_v0Wen;
    rand bit         io_diffCommits_info_28_vlWen;
    rand bit [5:0]   io_diffCommits_info_29_ldest;
    rand bit [7:0]   io_diffCommits_info_29_pdest;
    rand bit         io_diffCommits_info_29_rfWen;
    rand bit         io_diffCommits_info_29_fpWen;
    rand bit         io_diffCommits_info_29_vecWen;
    rand bit         io_diffCommits_info_29_v0Wen;
    rand bit         io_diffCommits_info_29_vlWen;
    rand bit [5:0]   io_diffCommits_info_30_ldest;
    rand bit [7:0]   io_diffCommits_info_30_pdest;
    rand bit         io_diffCommits_info_30_rfWen;
    rand bit         io_diffCommits_info_30_fpWen;
    rand bit         io_diffCommits_info_30_vecWen;
    rand bit         io_diffCommits_info_30_v0Wen;
    rand bit         io_diffCommits_info_30_vlWen;
    rand bit [5:0]   io_diffCommits_info_31_ldest;
    rand bit [7:0]   io_diffCommits_info_31_pdest;
    rand bit         io_diffCommits_info_31_rfWen;
    rand bit         io_diffCommits_info_31_fpWen;
    rand bit         io_diffCommits_info_31_vecWen;
    rand bit         io_diffCommits_info_31_v0Wen;
    rand bit         io_diffCommits_info_31_vlWen;
    rand bit [5:0]   io_diffCommits_info_32_ldest;
    rand bit [7:0]   io_diffCommits_info_32_pdest;
    rand bit         io_diffCommits_info_32_rfWen;
    rand bit         io_diffCommits_info_32_fpWen;
    rand bit         io_diffCommits_info_32_vecWen;
    rand bit         io_diffCommits_info_32_v0Wen;
    rand bit         io_diffCommits_info_32_vlWen;
    rand bit [5:0]   io_diffCommits_info_33_ldest;
    rand bit [7:0]   io_diffCommits_info_33_pdest;
    rand bit         io_diffCommits_info_33_rfWen;
    rand bit         io_diffCommits_info_33_fpWen;
    rand bit         io_diffCommits_info_33_vecWen;
    rand bit         io_diffCommits_info_33_v0Wen;
    rand bit         io_diffCommits_info_33_vlWen;
    rand bit [5:0]   io_diffCommits_info_34_ldest;
    rand bit [7:0]   io_diffCommits_info_34_pdest;
    rand bit         io_diffCommits_info_34_rfWen;
    rand bit         io_diffCommits_info_34_fpWen;
    rand bit         io_diffCommits_info_34_vecWen;
    rand bit         io_diffCommits_info_34_v0Wen;
    rand bit         io_diffCommits_info_34_vlWen;
    rand bit [5:0]   io_diffCommits_info_35_ldest;
    rand bit [7:0]   io_diffCommits_info_35_pdest;
    rand bit         io_diffCommits_info_35_rfWen;
    rand bit         io_diffCommits_info_35_fpWen;
    rand bit         io_diffCommits_info_35_vecWen;
    rand bit         io_diffCommits_info_35_v0Wen;
    rand bit         io_diffCommits_info_35_vlWen;
    rand bit [5:0]   io_diffCommits_info_36_ldest;
    rand bit [7:0]   io_diffCommits_info_36_pdest;
    rand bit         io_diffCommits_info_36_rfWen;
    rand bit         io_diffCommits_info_36_fpWen;
    rand bit         io_diffCommits_info_36_vecWen;
    rand bit         io_diffCommits_info_36_v0Wen;
    rand bit         io_diffCommits_info_36_vlWen;
    rand bit [5:0]   io_diffCommits_info_37_ldest;
    rand bit [7:0]   io_diffCommits_info_37_pdest;
    rand bit         io_diffCommits_info_37_rfWen;
    rand bit         io_diffCommits_info_37_fpWen;
    rand bit         io_diffCommits_info_37_vecWen;
    rand bit         io_diffCommits_info_37_v0Wen;
    rand bit         io_diffCommits_info_37_vlWen;
    rand bit [5:0]   io_diffCommits_info_38_ldest;
    rand bit [7:0]   io_diffCommits_info_38_pdest;
    rand bit         io_diffCommits_info_38_rfWen;
    rand bit         io_diffCommits_info_38_fpWen;
    rand bit         io_diffCommits_info_38_vecWen;
    rand bit         io_diffCommits_info_38_v0Wen;
    rand bit         io_diffCommits_info_38_vlWen;
    rand bit [5:0]   io_diffCommits_info_39_ldest;
    rand bit [7:0]   io_diffCommits_info_39_pdest;
    rand bit         io_diffCommits_info_39_rfWen;
    rand bit         io_diffCommits_info_39_fpWen;
    rand bit         io_diffCommits_info_39_vecWen;
    rand bit         io_diffCommits_info_39_v0Wen;
    rand bit         io_diffCommits_info_39_vlWen;
    rand bit [5:0]   io_diffCommits_info_40_ldest;
    rand bit [7:0]   io_diffCommits_info_40_pdest;
    rand bit         io_diffCommits_info_40_rfWen;
    rand bit         io_diffCommits_info_40_fpWen;
    rand bit         io_diffCommits_info_40_vecWen;
    rand bit         io_diffCommits_info_40_v0Wen;
    rand bit         io_diffCommits_info_40_vlWen;
    rand bit [5:0]   io_diffCommits_info_41_ldest;
    rand bit [7:0]   io_diffCommits_info_41_pdest;
    rand bit         io_diffCommits_info_41_rfWen;
    rand bit         io_diffCommits_info_41_fpWen;
    rand bit         io_diffCommits_info_41_vecWen;
    rand bit         io_diffCommits_info_41_v0Wen;
    rand bit         io_diffCommits_info_41_vlWen;
    rand bit [5:0]   io_diffCommits_info_42_ldest;
    rand bit [7:0]   io_diffCommits_info_42_pdest;
    rand bit         io_diffCommits_info_42_rfWen;
    rand bit         io_diffCommits_info_42_fpWen;
    rand bit         io_diffCommits_info_42_vecWen;
    rand bit         io_diffCommits_info_42_v0Wen;
    rand bit         io_diffCommits_info_42_vlWen;
    rand bit [5:0]   io_diffCommits_info_43_ldest;
    rand bit [7:0]   io_diffCommits_info_43_pdest;
    rand bit         io_diffCommits_info_43_rfWen;
    rand bit         io_diffCommits_info_43_fpWen;
    rand bit         io_diffCommits_info_43_vecWen;
    rand bit         io_diffCommits_info_43_v0Wen;
    rand bit         io_diffCommits_info_43_vlWen;
    rand bit [5:0]   io_diffCommits_info_44_ldest;
    rand bit [7:0]   io_diffCommits_info_44_pdest;
    rand bit         io_diffCommits_info_44_rfWen;
    rand bit         io_diffCommits_info_44_fpWen;
    rand bit         io_diffCommits_info_44_vecWen;
    rand bit         io_diffCommits_info_44_v0Wen;
    rand bit         io_diffCommits_info_44_vlWen;
    rand bit [5:0]   io_diffCommits_info_45_ldest;
    rand bit [7:0]   io_diffCommits_info_45_pdest;
    rand bit         io_diffCommits_info_45_rfWen;
    rand bit         io_diffCommits_info_45_fpWen;
    rand bit         io_diffCommits_info_45_vecWen;
    rand bit         io_diffCommits_info_45_v0Wen;
    rand bit         io_diffCommits_info_45_vlWen;
    rand bit [5:0]   io_diffCommits_info_46_ldest;
    rand bit [7:0]   io_diffCommits_info_46_pdest;
    rand bit         io_diffCommits_info_46_rfWen;
    rand bit         io_diffCommits_info_46_fpWen;
    rand bit         io_diffCommits_info_46_vecWen;
    rand bit         io_diffCommits_info_46_v0Wen;
    rand bit         io_diffCommits_info_46_vlWen;
    rand bit [5:0]   io_diffCommits_info_47_ldest;
    rand bit [7:0]   io_diffCommits_info_47_pdest;
    rand bit         io_diffCommits_info_47_rfWen;
    rand bit         io_diffCommits_info_47_fpWen;
    rand bit         io_diffCommits_info_47_vecWen;
    rand bit         io_diffCommits_info_47_v0Wen;
    rand bit         io_diffCommits_info_47_vlWen;
    rand bit [5:0]   io_diffCommits_info_48_ldest;
    rand bit [7:0]   io_diffCommits_info_48_pdest;
    rand bit         io_diffCommits_info_48_rfWen;
    rand bit         io_diffCommits_info_48_fpWen;
    rand bit         io_diffCommits_info_48_vecWen;
    rand bit         io_diffCommits_info_48_v0Wen;
    rand bit         io_diffCommits_info_48_vlWen;
    rand bit [5:0]   io_diffCommits_info_49_ldest;
    rand bit [7:0]   io_diffCommits_info_49_pdest;
    rand bit         io_diffCommits_info_49_rfWen;
    rand bit         io_diffCommits_info_49_fpWen;
    rand bit         io_diffCommits_info_49_vecWen;
    rand bit         io_diffCommits_info_49_v0Wen;
    rand bit         io_diffCommits_info_49_vlWen;
    rand bit [5:0]   io_diffCommits_info_50_ldest;
    rand bit [7:0]   io_diffCommits_info_50_pdest;
    rand bit         io_diffCommits_info_50_rfWen;
    rand bit         io_diffCommits_info_50_fpWen;
    rand bit         io_diffCommits_info_50_vecWen;
    rand bit         io_diffCommits_info_50_v0Wen;
    rand bit         io_diffCommits_info_50_vlWen;
    rand bit [5:0]   io_diffCommits_info_51_ldest;
    rand bit [7:0]   io_diffCommits_info_51_pdest;
    rand bit         io_diffCommits_info_51_rfWen;
    rand bit         io_diffCommits_info_51_fpWen;
    rand bit         io_diffCommits_info_51_vecWen;
    rand bit         io_diffCommits_info_51_v0Wen;
    rand bit         io_diffCommits_info_51_vlWen;
    rand bit [5:0]   io_diffCommits_info_52_ldest;
    rand bit [7:0]   io_diffCommits_info_52_pdest;
    rand bit         io_diffCommits_info_52_rfWen;
    rand bit         io_diffCommits_info_52_fpWen;
    rand bit         io_diffCommits_info_52_vecWen;
    rand bit         io_diffCommits_info_52_v0Wen;
    rand bit         io_diffCommits_info_52_vlWen;
    rand bit [5:0]   io_diffCommits_info_53_ldest;
    rand bit [7:0]   io_diffCommits_info_53_pdest;
    rand bit         io_diffCommits_info_53_rfWen;
    rand bit         io_diffCommits_info_53_fpWen;
    rand bit         io_diffCommits_info_53_vecWen;
    rand bit         io_diffCommits_info_53_v0Wen;
    rand bit         io_diffCommits_info_53_vlWen;
    rand bit [5:0]   io_diffCommits_info_54_ldest;
    rand bit [7:0]   io_diffCommits_info_54_pdest;
    rand bit         io_diffCommits_info_54_rfWen;
    rand bit         io_diffCommits_info_54_fpWen;
    rand bit         io_diffCommits_info_54_vecWen;
    rand bit         io_diffCommits_info_54_v0Wen;
    rand bit         io_diffCommits_info_54_vlWen;
    rand bit [5:0]   io_diffCommits_info_55_ldest;
    rand bit [7:0]   io_diffCommits_info_55_pdest;
    rand bit         io_diffCommits_info_55_rfWen;
    rand bit         io_diffCommits_info_55_fpWen;
    rand bit         io_diffCommits_info_55_vecWen;
    rand bit         io_diffCommits_info_55_v0Wen;
    rand bit         io_diffCommits_info_55_vlWen;
    rand bit [5:0]   io_diffCommits_info_56_ldest;
    rand bit [7:0]   io_diffCommits_info_56_pdest;
    rand bit         io_diffCommits_info_56_rfWen;
    rand bit         io_diffCommits_info_56_fpWen;
    rand bit         io_diffCommits_info_56_vecWen;
    rand bit         io_diffCommits_info_56_v0Wen;
    rand bit         io_diffCommits_info_56_vlWen;
    rand bit [5:0]   io_diffCommits_info_57_ldest;
    rand bit [7:0]   io_diffCommits_info_57_pdest;
    rand bit         io_diffCommits_info_57_rfWen;
    rand bit         io_diffCommits_info_57_fpWen;
    rand bit         io_diffCommits_info_57_vecWen;
    rand bit         io_diffCommits_info_57_v0Wen;
    rand bit         io_diffCommits_info_57_vlWen;
    rand bit [5:0]   io_diffCommits_info_58_ldest;
    rand bit [7:0]   io_diffCommits_info_58_pdest;
    rand bit         io_diffCommits_info_58_rfWen;
    rand bit         io_diffCommits_info_58_fpWen;
    rand bit         io_diffCommits_info_58_vecWen;
    rand bit         io_diffCommits_info_58_v0Wen;
    rand bit         io_diffCommits_info_58_vlWen;
    rand bit [5:0]   io_diffCommits_info_59_ldest;
    rand bit [7:0]   io_diffCommits_info_59_pdest;
    rand bit         io_diffCommits_info_59_rfWen;
    rand bit         io_diffCommits_info_59_fpWen;
    rand bit         io_diffCommits_info_59_vecWen;
    rand bit         io_diffCommits_info_59_v0Wen;
    rand bit         io_diffCommits_info_59_vlWen;
    rand bit [5:0]   io_diffCommits_info_60_ldest;
    rand bit [7:0]   io_diffCommits_info_60_pdest;
    rand bit         io_diffCommits_info_60_rfWen;
    rand bit         io_diffCommits_info_60_fpWen;
    rand bit         io_diffCommits_info_60_vecWen;
    rand bit         io_diffCommits_info_60_v0Wen;
    rand bit         io_diffCommits_info_60_vlWen;
    rand bit [5:0]   io_diffCommits_info_61_ldest;
    rand bit [7:0]   io_diffCommits_info_61_pdest;
    rand bit         io_diffCommits_info_61_rfWen;
    rand bit         io_diffCommits_info_61_fpWen;
    rand bit         io_diffCommits_info_61_vecWen;
    rand bit         io_diffCommits_info_61_v0Wen;
    rand bit         io_diffCommits_info_61_vlWen;
    rand bit [5:0]   io_diffCommits_info_62_ldest;
    rand bit [7:0]   io_diffCommits_info_62_pdest;
    rand bit         io_diffCommits_info_62_rfWen;
    rand bit         io_diffCommits_info_62_fpWen;
    rand bit         io_diffCommits_info_62_vecWen;
    rand bit         io_diffCommits_info_62_v0Wen;
    rand bit         io_diffCommits_info_62_vlWen;
    rand bit [5:0]   io_diffCommits_info_63_ldest;
    rand bit [7:0]   io_diffCommits_info_63_pdest;
    rand bit         io_diffCommits_info_63_rfWen;
    rand bit         io_diffCommits_info_63_fpWen;
    rand bit         io_diffCommits_info_63_vecWen;
    rand bit         io_diffCommits_info_63_v0Wen;
    rand bit         io_diffCommits_info_63_vlWen;
    rand bit [5:0]   io_diffCommits_info_64_ldest;
    rand bit [7:0]   io_diffCommits_info_64_pdest;
    rand bit         io_diffCommits_info_64_rfWen;
    rand bit         io_diffCommits_info_64_fpWen;
    rand bit         io_diffCommits_info_64_vecWen;
    rand bit         io_diffCommits_info_64_v0Wen;
    rand bit         io_diffCommits_info_64_vlWen;
    rand bit [5:0]   io_diffCommits_info_65_ldest;
    rand bit [7:0]   io_diffCommits_info_65_pdest;
    rand bit         io_diffCommits_info_65_rfWen;
    rand bit         io_diffCommits_info_65_fpWen;
    rand bit         io_diffCommits_info_65_vecWen;
    rand bit         io_diffCommits_info_65_v0Wen;
    rand bit         io_diffCommits_info_65_vlWen;
    rand bit [5:0]   io_diffCommits_info_66_ldest;
    rand bit [7:0]   io_diffCommits_info_66_pdest;
    rand bit         io_diffCommits_info_66_rfWen;
    rand bit         io_diffCommits_info_66_fpWen;
    rand bit         io_diffCommits_info_66_vecWen;
    rand bit         io_diffCommits_info_66_v0Wen;
    rand bit         io_diffCommits_info_66_vlWen;
    rand bit [5:0]   io_diffCommits_info_67_ldest;
    rand bit [7:0]   io_diffCommits_info_67_pdest;
    rand bit         io_diffCommits_info_67_rfWen;
    rand bit         io_diffCommits_info_67_fpWen;
    rand bit         io_diffCommits_info_67_vecWen;
    rand bit         io_diffCommits_info_67_v0Wen;
    rand bit         io_diffCommits_info_67_vlWen;
    rand bit [5:0]   io_diffCommits_info_68_ldest;
    rand bit [7:0]   io_diffCommits_info_68_pdest;
    rand bit         io_diffCommits_info_68_rfWen;
    rand bit         io_diffCommits_info_68_fpWen;
    rand bit         io_diffCommits_info_68_vecWen;
    rand bit         io_diffCommits_info_68_v0Wen;
    rand bit         io_diffCommits_info_68_vlWen;
    rand bit [5:0]   io_diffCommits_info_69_ldest;
    rand bit [7:0]   io_diffCommits_info_69_pdest;
    rand bit         io_diffCommits_info_69_rfWen;
    rand bit         io_diffCommits_info_69_fpWen;
    rand bit         io_diffCommits_info_69_vecWen;
    rand bit         io_diffCommits_info_69_v0Wen;
    rand bit         io_diffCommits_info_69_vlWen;
    rand bit [5:0]   io_diffCommits_info_70_ldest;
    rand bit [7:0]   io_diffCommits_info_70_pdest;
    rand bit         io_diffCommits_info_70_rfWen;
    rand bit         io_diffCommits_info_70_fpWen;
    rand bit         io_diffCommits_info_70_vecWen;
    rand bit         io_diffCommits_info_70_v0Wen;
    rand bit         io_diffCommits_info_70_vlWen;
    rand bit [5:0]   io_diffCommits_info_71_ldest;
    rand bit [7:0]   io_diffCommits_info_71_pdest;
    rand bit         io_diffCommits_info_71_rfWen;
    rand bit         io_diffCommits_info_71_fpWen;
    rand bit         io_diffCommits_info_71_vecWen;
    rand bit         io_diffCommits_info_71_v0Wen;
    rand bit         io_diffCommits_info_71_vlWen;
    rand bit [5:0]   io_diffCommits_info_72_ldest;
    rand bit [7:0]   io_diffCommits_info_72_pdest;
    rand bit         io_diffCommits_info_72_rfWen;
    rand bit         io_diffCommits_info_72_fpWen;
    rand bit         io_diffCommits_info_72_vecWen;
    rand bit         io_diffCommits_info_72_v0Wen;
    rand bit         io_diffCommits_info_72_vlWen;
    rand bit [5:0]   io_diffCommits_info_73_ldest;
    rand bit [7:0]   io_diffCommits_info_73_pdest;
    rand bit         io_diffCommits_info_73_rfWen;
    rand bit         io_diffCommits_info_73_fpWen;
    rand bit         io_diffCommits_info_73_vecWen;
    rand bit         io_diffCommits_info_73_v0Wen;
    rand bit         io_diffCommits_info_73_vlWen;
    rand bit [5:0]   io_diffCommits_info_74_ldest;
    rand bit [7:0]   io_diffCommits_info_74_pdest;
    rand bit         io_diffCommits_info_74_rfWen;
    rand bit         io_diffCommits_info_74_fpWen;
    rand bit         io_diffCommits_info_74_vecWen;
    rand bit         io_diffCommits_info_74_v0Wen;
    rand bit         io_diffCommits_info_74_vlWen;
    rand bit [5:0]   io_diffCommits_info_75_ldest;
    rand bit [7:0]   io_diffCommits_info_75_pdest;
    rand bit         io_diffCommits_info_75_rfWen;
    rand bit         io_diffCommits_info_75_fpWen;
    rand bit         io_diffCommits_info_75_vecWen;
    rand bit         io_diffCommits_info_75_v0Wen;
    rand bit         io_diffCommits_info_75_vlWen;
    rand bit [5:0]   io_diffCommits_info_76_ldest;
    rand bit [7:0]   io_diffCommits_info_76_pdest;
    rand bit         io_diffCommits_info_76_rfWen;
    rand bit         io_diffCommits_info_76_fpWen;
    rand bit         io_diffCommits_info_76_vecWen;
    rand bit         io_diffCommits_info_76_v0Wen;
    rand bit         io_diffCommits_info_76_vlWen;
    rand bit [5:0]   io_diffCommits_info_77_ldest;
    rand bit [7:0]   io_diffCommits_info_77_pdest;
    rand bit         io_diffCommits_info_77_rfWen;
    rand bit         io_diffCommits_info_77_fpWen;
    rand bit         io_diffCommits_info_77_vecWen;
    rand bit         io_diffCommits_info_77_v0Wen;
    rand bit         io_diffCommits_info_77_vlWen;
    rand bit [5:0]   io_diffCommits_info_78_ldest;
    rand bit [7:0]   io_diffCommits_info_78_pdest;
    rand bit         io_diffCommits_info_78_rfWen;
    rand bit         io_diffCommits_info_78_fpWen;
    rand bit         io_diffCommits_info_78_vecWen;
    rand bit         io_diffCommits_info_78_v0Wen;
    rand bit         io_diffCommits_info_78_vlWen;
    rand bit [5:0]   io_diffCommits_info_79_ldest;
    rand bit [7:0]   io_diffCommits_info_79_pdest;
    rand bit         io_diffCommits_info_79_rfWen;
    rand bit         io_diffCommits_info_79_fpWen;
    rand bit         io_diffCommits_info_79_vecWen;
    rand bit         io_diffCommits_info_79_v0Wen;
    rand bit         io_diffCommits_info_79_vlWen;
    rand bit [5:0]   io_diffCommits_info_80_ldest;
    rand bit [7:0]   io_diffCommits_info_80_pdest;
    rand bit         io_diffCommits_info_80_rfWen;
    rand bit         io_diffCommits_info_80_fpWen;
    rand bit         io_diffCommits_info_80_vecWen;
    rand bit         io_diffCommits_info_80_v0Wen;
    rand bit         io_diffCommits_info_80_vlWen;
    rand bit [5:0]   io_diffCommits_info_81_ldest;
    rand bit [7:0]   io_diffCommits_info_81_pdest;
    rand bit         io_diffCommits_info_81_rfWen;
    rand bit         io_diffCommits_info_81_fpWen;
    rand bit         io_diffCommits_info_81_vecWen;
    rand bit         io_diffCommits_info_81_v0Wen;
    rand bit         io_diffCommits_info_81_vlWen;
    rand bit [5:0]   io_diffCommits_info_82_ldest;
    rand bit [7:0]   io_diffCommits_info_82_pdest;
    rand bit         io_diffCommits_info_82_rfWen;
    rand bit         io_diffCommits_info_82_fpWen;
    rand bit         io_diffCommits_info_82_vecWen;
    rand bit         io_diffCommits_info_82_v0Wen;
    rand bit         io_diffCommits_info_82_vlWen;
    rand bit [5:0]   io_diffCommits_info_83_ldest;
    rand bit [7:0]   io_diffCommits_info_83_pdest;
    rand bit         io_diffCommits_info_83_rfWen;
    rand bit         io_diffCommits_info_83_fpWen;
    rand bit         io_diffCommits_info_83_vecWen;
    rand bit         io_diffCommits_info_83_v0Wen;
    rand bit         io_diffCommits_info_83_vlWen;
    rand bit [5:0]   io_diffCommits_info_84_ldest;
    rand bit [7:0]   io_diffCommits_info_84_pdest;
    rand bit         io_diffCommits_info_84_rfWen;
    rand bit         io_diffCommits_info_84_fpWen;
    rand bit         io_diffCommits_info_84_vecWen;
    rand bit         io_diffCommits_info_84_v0Wen;
    rand bit         io_diffCommits_info_84_vlWen;
    rand bit [5:0]   io_diffCommits_info_85_ldest;
    rand bit [7:0]   io_diffCommits_info_85_pdest;
    rand bit         io_diffCommits_info_85_rfWen;
    rand bit         io_diffCommits_info_85_fpWen;
    rand bit         io_diffCommits_info_85_vecWen;
    rand bit         io_diffCommits_info_85_v0Wen;
    rand bit         io_diffCommits_info_85_vlWen;
    rand bit [5:0]   io_diffCommits_info_86_ldest;
    rand bit [7:0]   io_diffCommits_info_86_pdest;
    rand bit         io_diffCommits_info_86_rfWen;
    rand bit         io_diffCommits_info_86_fpWen;
    rand bit         io_diffCommits_info_86_vecWen;
    rand bit         io_diffCommits_info_86_v0Wen;
    rand bit         io_diffCommits_info_86_vlWen;
    rand bit [5:0]   io_diffCommits_info_87_ldest;
    rand bit [7:0]   io_diffCommits_info_87_pdest;
    rand bit         io_diffCommits_info_87_rfWen;
    rand bit         io_diffCommits_info_87_fpWen;
    rand bit         io_diffCommits_info_87_vecWen;
    rand bit         io_diffCommits_info_87_v0Wen;
    rand bit         io_diffCommits_info_87_vlWen;
    rand bit [5:0]   io_diffCommits_info_88_ldest;
    rand bit [7:0]   io_diffCommits_info_88_pdest;
    rand bit         io_diffCommits_info_88_rfWen;
    rand bit         io_diffCommits_info_88_fpWen;
    rand bit         io_diffCommits_info_88_vecWen;
    rand bit         io_diffCommits_info_88_v0Wen;
    rand bit         io_diffCommits_info_88_vlWen;
    rand bit [5:0]   io_diffCommits_info_89_ldest;
    rand bit [7:0]   io_diffCommits_info_89_pdest;
    rand bit         io_diffCommits_info_89_rfWen;
    rand bit         io_diffCommits_info_89_fpWen;
    rand bit         io_diffCommits_info_89_vecWen;
    rand bit         io_diffCommits_info_89_v0Wen;
    rand bit         io_diffCommits_info_89_vlWen;
    rand bit [5:0]   io_diffCommits_info_90_ldest;
    rand bit [7:0]   io_diffCommits_info_90_pdest;
    rand bit         io_diffCommits_info_90_rfWen;
    rand bit         io_diffCommits_info_90_fpWen;
    rand bit         io_diffCommits_info_90_vecWen;
    rand bit         io_diffCommits_info_90_v0Wen;
    rand bit         io_diffCommits_info_90_vlWen;
    rand bit [5:0]   io_diffCommits_info_91_ldest;
    rand bit [7:0]   io_diffCommits_info_91_pdest;
    rand bit         io_diffCommits_info_91_rfWen;
    rand bit         io_diffCommits_info_91_fpWen;
    rand bit         io_diffCommits_info_91_vecWen;
    rand bit         io_diffCommits_info_91_v0Wen;
    rand bit         io_diffCommits_info_91_vlWen;
    rand bit [5:0]   io_diffCommits_info_92_ldest;
    rand bit [7:0]   io_diffCommits_info_92_pdest;
    rand bit         io_diffCommits_info_92_rfWen;
    rand bit         io_diffCommits_info_92_fpWen;
    rand bit         io_diffCommits_info_92_vecWen;
    rand bit         io_diffCommits_info_92_v0Wen;
    rand bit         io_diffCommits_info_92_vlWen;
    rand bit [5:0]   io_diffCommits_info_93_ldest;
    rand bit [7:0]   io_diffCommits_info_93_pdest;
    rand bit         io_diffCommits_info_93_rfWen;
    rand bit         io_diffCommits_info_93_fpWen;
    rand bit         io_diffCommits_info_93_vecWen;
    rand bit         io_diffCommits_info_93_v0Wen;
    rand bit         io_diffCommits_info_93_vlWen;
    rand bit [5:0]   io_diffCommits_info_94_ldest;
    rand bit [7:0]   io_diffCommits_info_94_pdest;
    rand bit         io_diffCommits_info_94_rfWen;
    rand bit         io_diffCommits_info_94_fpWen;
    rand bit         io_diffCommits_info_94_vecWen;
    rand bit         io_diffCommits_info_94_v0Wen;
    rand bit         io_diffCommits_info_94_vlWen;
    rand bit [5:0]   io_diffCommits_info_95_ldest;
    rand bit [7:0]   io_diffCommits_info_95_pdest;
    rand bit         io_diffCommits_info_95_rfWen;
    rand bit         io_diffCommits_info_95_fpWen;
    rand bit         io_diffCommits_info_95_vecWen;
    rand bit         io_diffCommits_info_95_v0Wen;
    rand bit         io_diffCommits_info_95_vlWen;
    rand bit [5:0]   io_diffCommits_info_96_ldest;
    rand bit [7:0]   io_diffCommits_info_96_pdest;
    rand bit         io_diffCommits_info_96_rfWen;
    rand bit         io_diffCommits_info_96_fpWen;
    rand bit         io_diffCommits_info_96_vecWen;
    rand bit         io_diffCommits_info_96_v0Wen;
    rand bit         io_diffCommits_info_96_vlWen;
    rand bit [5:0]   io_diffCommits_info_97_ldest;
    rand bit [7:0]   io_diffCommits_info_97_pdest;
    rand bit         io_diffCommits_info_97_rfWen;
    rand bit         io_diffCommits_info_97_fpWen;
    rand bit         io_diffCommits_info_97_vecWen;
    rand bit         io_diffCommits_info_97_v0Wen;
    rand bit         io_diffCommits_info_97_vlWen;
    rand bit [5:0]   io_diffCommits_info_98_ldest;
    rand bit [7:0]   io_diffCommits_info_98_pdest;
    rand bit         io_diffCommits_info_98_rfWen;
    rand bit         io_diffCommits_info_98_fpWen;
    rand bit         io_diffCommits_info_98_vecWen;
    rand bit         io_diffCommits_info_98_v0Wen;
    rand bit         io_diffCommits_info_98_vlWen;
    rand bit [5:0]   io_diffCommits_info_99_ldest;
    rand bit [7:0]   io_diffCommits_info_99_pdest;
    rand bit         io_diffCommits_info_99_rfWen;
    rand bit         io_diffCommits_info_99_fpWen;
    rand bit         io_diffCommits_info_99_vecWen;
    rand bit         io_diffCommits_info_99_v0Wen;
    rand bit         io_diffCommits_info_99_vlWen;
    rand bit [5:0]   io_diffCommits_info_100_ldest;
    rand bit [7:0]   io_diffCommits_info_100_pdest;
    rand bit         io_diffCommits_info_100_rfWen;
    rand bit         io_diffCommits_info_100_fpWen;
    rand bit         io_diffCommits_info_100_vecWen;
    rand bit         io_diffCommits_info_100_v0Wen;
    rand bit         io_diffCommits_info_100_vlWen;
    rand bit [5:0]   io_diffCommits_info_101_ldest;
    rand bit [7:0]   io_diffCommits_info_101_pdest;
    rand bit         io_diffCommits_info_101_rfWen;
    rand bit         io_diffCommits_info_101_fpWen;
    rand bit         io_diffCommits_info_101_vecWen;
    rand bit         io_diffCommits_info_101_v0Wen;
    rand bit         io_diffCommits_info_101_vlWen;
    rand bit [5:0]   io_diffCommits_info_102_ldest;
    rand bit [7:0]   io_diffCommits_info_102_pdest;
    rand bit         io_diffCommits_info_102_rfWen;
    rand bit         io_diffCommits_info_102_fpWen;
    rand bit         io_diffCommits_info_102_vecWen;
    rand bit         io_diffCommits_info_102_v0Wen;
    rand bit         io_diffCommits_info_102_vlWen;
    rand bit [5:0]   io_diffCommits_info_103_ldest;
    rand bit [7:0]   io_diffCommits_info_103_pdest;
    rand bit         io_diffCommits_info_103_rfWen;
    rand bit         io_diffCommits_info_103_fpWen;
    rand bit         io_diffCommits_info_103_vecWen;
    rand bit         io_diffCommits_info_103_v0Wen;
    rand bit         io_diffCommits_info_103_vlWen;
    rand bit [5:0]   io_diffCommits_info_104_ldest;
    rand bit [7:0]   io_diffCommits_info_104_pdest;
    rand bit         io_diffCommits_info_104_rfWen;
    rand bit         io_diffCommits_info_104_fpWen;
    rand bit         io_diffCommits_info_104_vecWen;
    rand bit         io_diffCommits_info_104_v0Wen;
    rand bit         io_diffCommits_info_104_vlWen;
    rand bit [5:0]   io_diffCommits_info_105_ldest;
    rand bit [7:0]   io_diffCommits_info_105_pdest;
    rand bit         io_diffCommits_info_105_rfWen;
    rand bit         io_diffCommits_info_105_fpWen;
    rand bit         io_diffCommits_info_105_vecWen;
    rand bit         io_diffCommits_info_105_v0Wen;
    rand bit         io_diffCommits_info_105_vlWen;
    rand bit [5:0]   io_diffCommits_info_106_ldest;
    rand bit [7:0]   io_diffCommits_info_106_pdest;
    rand bit         io_diffCommits_info_106_rfWen;
    rand bit         io_diffCommits_info_106_fpWen;
    rand bit         io_diffCommits_info_106_vecWen;
    rand bit         io_diffCommits_info_106_v0Wen;
    rand bit         io_diffCommits_info_106_vlWen;
    rand bit [5:0]   io_diffCommits_info_107_ldest;
    rand bit [7:0]   io_diffCommits_info_107_pdest;
    rand bit         io_diffCommits_info_107_rfWen;
    rand bit         io_diffCommits_info_107_fpWen;
    rand bit         io_diffCommits_info_107_vecWen;
    rand bit         io_diffCommits_info_107_v0Wen;
    rand bit         io_diffCommits_info_107_vlWen;
    rand bit [5:0]   io_diffCommits_info_108_ldest;
    rand bit [7:0]   io_diffCommits_info_108_pdest;
    rand bit         io_diffCommits_info_108_rfWen;
    rand bit         io_diffCommits_info_108_fpWen;
    rand bit         io_diffCommits_info_108_vecWen;
    rand bit         io_diffCommits_info_108_v0Wen;
    rand bit         io_diffCommits_info_108_vlWen;
    rand bit [5:0]   io_diffCommits_info_109_ldest;
    rand bit [7:0]   io_diffCommits_info_109_pdest;
    rand bit         io_diffCommits_info_109_rfWen;
    rand bit         io_diffCommits_info_109_fpWen;
    rand bit         io_diffCommits_info_109_vecWen;
    rand bit         io_diffCommits_info_109_v0Wen;
    rand bit         io_diffCommits_info_109_vlWen;
    rand bit [5:0]   io_diffCommits_info_110_ldest;
    rand bit [7:0]   io_diffCommits_info_110_pdest;
    rand bit         io_diffCommits_info_110_rfWen;
    rand bit         io_diffCommits_info_110_fpWen;
    rand bit         io_diffCommits_info_110_vecWen;
    rand bit         io_diffCommits_info_110_v0Wen;
    rand bit         io_diffCommits_info_110_vlWen;
    rand bit [5:0]   io_diffCommits_info_111_ldest;
    rand bit [7:0]   io_diffCommits_info_111_pdest;
    rand bit         io_diffCommits_info_111_rfWen;
    rand bit         io_diffCommits_info_111_fpWen;
    rand bit         io_diffCommits_info_111_vecWen;
    rand bit         io_diffCommits_info_111_v0Wen;
    rand bit         io_diffCommits_info_111_vlWen;
    rand bit [5:0]   io_diffCommits_info_112_ldest;
    rand bit [7:0]   io_diffCommits_info_112_pdest;
    rand bit         io_diffCommits_info_112_rfWen;
    rand bit         io_diffCommits_info_112_fpWen;
    rand bit         io_diffCommits_info_112_vecWen;
    rand bit         io_diffCommits_info_112_v0Wen;
    rand bit         io_diffCommits_info_112_vlWen;
    rand bit [5:0]   io_diffCommits_info_113_ldest;
    rand bit [7:0]   io_diffCommits_info_113_pdest;
    rand bit         io_diffCommits_info_113_rfWen;
    rand bit         io_diffCommits_info_113_fpWen;
    rand bit         io_diffCommits_info_113_vecWen;
    rand bit         io_diffCommits_info_113_v0Wen;
    rand bit         io_diffCommits_info_113_vlWen;
    rand bit [5:0]   io_diffCommits_info_114_ldest;
    rand bit [7:0]   io_diffCommits_info_114_pdest;
    rand bit         io_diffCommits_info_114_rfWen;
    rand bit         io_diffCommits_info_114_fpWen;
    rand bit         io_diffCommits_info_114_vecWen;
    rand bit         io_diffCommits_info_114_v0Wen;
    rand bit         io_diffCommits_info_114_vlWen;
    rand bit [5:0]   io_diffCommits_info_115_ldest;
    rand bit [7:0]   io_diffCommits_info_115_pdest;
    rand bit         io_diffCommits_info_115_rfWen;
    rand bit         io_diffCommits_info_115_fpWen;
    rand bit         io_diffCommits_info_115_vecWen;
    rand bit         io_diffCommits_info_115_v0Wen;
    rand bit         io_diffCommits_info_115_vlWen;
    rand bit [5:0]   io_diffCommits_info_116_ldest;
    rand bit [7:0]   io_diffCommits_info_116_pdest;
    rand bit         io_diffCommits_info_116_rfWen;
    rand bit         io_diffCommits_info_116_fpWen;
    rand bit         io_diffCommits_info_116_vecWen;
    rand bit         io_diffCommits_info_116_v0Wen;
    rand bit         io_diffCommits_info_116_vlWen;
    rand bit [5:0]   io_diffCommits_info_117_ldest;
    rand bit [7:0]   io_diffCommits_info_117_pdest;
    rand bit         io_diffCommits_info_117_rfWen;
    rand bit         io_diffCommits_info_117_fpWen;
    rand bit         io_diffCommits_info_117_vecWen;
    rand bit         io_diffCommits_info_117_v0Wen;
    rand bit         io_diffCommits_info_117_vlWen;
    rand bit [5:0]   io_diffCommits_info_118_ldest;
    rand bit [7:0]   io_diffCommits_info_118_pdest;
    rand bit         io_diffCommits_info_118_rfWen;
    rand bit         io_diffCommits_info_118_fpWen;
    rand bit         io_diffCommits_info_118_vecWen;
    rand bit         io_diffCommits_info_118_v0Wen;
    rand bit         io_diffCommits_info_118_vlWen;
    rand bit [5:0]   io_diffCommits_info_119_ldest;
    rand bit [7:0]   io_diffCommits_info_119_pdest;
    rand bit         io_diffCommits_info_119_rfWen;
    rand bit         io_diffCommits_info_119_fpWen;
    rand bit         io_diffCommits_info_119_vecWen;
    rand bit         io_diffCommits_info_119_v0Wen;
    rand bit         io_diffCommits_info_119_vlWen;
    rand bit [5:0]   io_diffCommits_info_120_ldest;
    rand bit [7:0]   io_diffCommits_info_120_pdest;
    rand bit         io_diffCommits_info_120_rfWen;
    rand bit         io_diffCommits_info_120_fpWen;
    rand bit         io_diffCommits_info_120_vecWen;
    rand bit         io_diffCommits_info_120_v0Wen;
    rand bit         io_diffCommits_info_120_vlWen;
    rand bit [5:0]   io_diffCommits_info_121_ldest;
    rand bit [7:0]   io_diffCommits_info_121_pdest;
    rand bit         io_diffCommits_info_121_rfWen;
    rand bit         io_diffCommits_info_121_fpWen;
    rand bit         io_diffCommits_info_121_vecWen;
    rand bit         io_diffCommits_info_121_v0Wen;
    rand bit         io_diffCommits_info_121_vlWen;
    rand bit [5:0]   io_diffCommits_info_122_ldest;
    rand bit [7:0]   io_diffCommits_info_122_pdest;
    rand bit         io_diffCommits_info_122_rfWen;
    rand bit         io_diffCommits_info_122_fpWen;
    rand bit         io_diffCommits_info_122_vecWen;
    rand bit         io_diffCommits_info_122_v0Wen;
    rand bit         io_diffCommits_info_122_vlWen;
    rand bit [5:0]   io_diffCommits_info_123_ldest;
    rand bit [7:0]   io_diffCommits_info_123_pdest;
    rand bit         io_diffCommits_info_123_rfWen;
    rand bit         io_diffCommits_info_123_fpWen;
    rand bit         io_diffCommits_info_123_vecWen;
    rand bit         io_diffCommits_info_123_v0Wen;
    rand bit         io_diffCommits_info_123_vlWen;
    rand bit [5:0]   io_diffCommits_info_124_ldest;
    rand bit [7:0]   io_diffCommits_info_124_pdest;
    rand bit         io_diffCommits_info_124_rfWen;
    rand bit         io_diffCommits_info_124_fpWen;
    rand bit         io_diffCommits_info_124_vecWen;
    rand bit         io_diffCommits_info_124_v0Wen;
    rand bit         io_diffCommits_info_124_vlWen;
    rand bit [5:0]   io_diffCommits_info_125_ldest;
    rand bit [7:0]   io_diffCommits_info_125_pdest;
    rand bit         io_diffCommits_info_125_rfWen;
    rand bit         io_diffCommits_info_125_fpWen;
    rand bit         io_diffCommits_info_125_vecWen;
    rand bit         io_diffCommits_info_125_v0Wen;
    rand bit         io_diffCommits_info_125_vlWen;
    rand bit [5:0]   io_diffCommits_info_126_ldest;
    rand bit [7:0]   io_diffCommits_info_126_pdest;
    rand bit         io_diffCommits_info_126_rfWen;
    rand bit         io_diffCommits_info_126_fpWen;
    rand bit         io_diffCommits_info_126_vecWen;
    rand bit         io_diffCommits_info_126_v0Wen;
    rand bit         io_diffCommits_info_126_vlWen;
    rand bit [5:0]   io_diffCommits_info_127_ldest;
    rand bit [7:0]   io_diffCommits_info_127_pdest;
    rand bit         io_diffCommits_info_127_rfWen;
    rand bit         io_diffCommits_info_127_fpWen;
    rand bit         io_diffCommits_info_127_vecWen;
    rand bit         io_diffCommits_info_127_v0Wen;
    rand bit         io_diffCommits_info_127_vlWen;
    rand bit [5:0]   io_diffCommits_info_128_ldest;
    rand bit [7:0]   io_diffCommits_info_128_pdest;
    rand bit         io_diffCommits_info_128_rfWen;
    rand bit         io_diffCommits_info_128_fpWen;
    rand bit         io_diffCommits_info_128_vecWen;
    rand bit         io_diffCommits_info_128_v0Wen;
    rand bit         io_diffCommits_info_128_vlWen;
    rand bit [5:0]   io_diffCommits_info_129_ldest;
    rand bit [7:0]   io_diffCommits_info_129_pdest;
    rand bit         io_diffCommits_info_129_rfWen;
    rand bit         io_diffCommits_info_129_fpWen;
    rand bit         io_diffCommits_info_129_vecWen;
    rand bit         io_diffCommits_info_129_v0Wen;
    rand bit         io_diffCommits_info_129_vlWen;
    rand bit [5:0]   io_diffCommits_info_130_ldest;
    rand bit [7:0]   io_diffCommits_info_130_pdest;
    rand bit         io_diffCommits_info_130_rfWen;
    rand bit         io_diffCommits_info_130_fpWen;
    rand bit         io_diffCommits_info_130_vecWen;
    rand bit         io_diffCommits_info_130_v0Wen;
    rand bit         io_diffCommits_info_130_vlWen;
    rand bit [5:0]   io_diffCommits_info_131_ldest;
    rand bit [7:0]   io_diffCommits_info_131_pdest;
    rand bit         io_diffCommits_info_131_rfWen;
    rand bit         io_diffCommits_info_131_fpWen;
    rand bit         io_diffCommits_info_131_vecWen;
    rand bit         io_diffCommits_info_131_v0Wen;
    rand bit         io_diffCommits_info_131_vlWen;
    rand bit [5:0]   io_diffCommits_info_132_ldest;
    rand bit [7:0]   io_diffCommits_info_132_pdest;
    rand bit         io_diffCommits_info_132_rfWen;
    rand bit         io_diffCommits_info_132_fpWen;
    rand bit         io_diffCommits_info_132_vecWen;
    rand bit         io_diffCommits_info_132_v0Wen;
    rand bit         io_diffCommits_info_132_vlWen;
    rand bit [5:0]   io_diffCommits_info_133_ldest;
    rand bit [7:0]   io_diffCommits_info_133_pdest;
    rand bit         io_diffCommits_info_133_rfWen;
    rand bit         io_diffCommits_info_133_fpWen;
    rand bit         io_diffCommits_info_133_vecWen;
    rand bit         io_diffCommits_info_133_v0Wen;
    rand bit         io_diffCommits_info_133_vlWen;
    rand bit [5:0]   io_diffCommits_info_134_ldest;
    rand bit [7:0]   io_diffCommits_info_134_pdest;
    rand bit         io_diffCommits_info_134_rfWen;
    rand bit         io_diffCommits_info_134_fpWen;
    rand bit         io_diffCommits_info_134_vecWen;
    rand bit         io_diffCommits_info_134_v0Wen;
    rand bit         io_diffCommits_info_134_vlWen;
    rand bit [5:0]   io_diffCommits_info_135_ldest;
    rand bit [7:0]   io_diffCommits_info_135_pdest;
    rand bit         io_diffCommits_info_135_rfWen;
    rand bit         io_diffCommits_info_135_fpWen;
    rand bit         io_diffCommits_info_135_vecWen;
    rand bit         io_diffCommits_info_135_v0Wen;
    rand bit         io_diffCommits_info_135_vlWen;
    rand bit [5:0]   io_diffCommits_info_136_ldest;
    rand bit [7:0]   io_diffCommits_info_136_pdest;
    rand bit         io_diffCommits_info_136_rfWen;
    rand bit         io_diffCommits_info_136_fpWen;
    rand bit         io_diffCommits_info_136_vecWen;
    rand bit         io_diffCommits_info_136_v0Wen;
    rand bit         io_diffCommits_info_136_vlWen;
    rand bit [5:0]   io_diffCommits_info_137_ldest;
    rand bit [7:0]   io_diffCommits_info_137_pdest;
    rand bit         io_diffCommits_info_137_rfWen;
    rand bit         io_diffCommits_info_137_fpWen;
    rand bit         io_diffCommits_info_137_vecWen;
    rand bit         io_diffCommits_info_137_v0Wen;
    rand bit         io_diffCommits_info_137_vlWen;
    rand bit [5:0]   io_diffCommits_info_138_ldest;
    rand bit [7:0]   io_diffCommits_info_138_pdest;
    rand bit         io_diffCommits_info_138_rfWen;
    rand bit         io_diffCommits_info_138_fpWen;
    rand bit         io_diffCommits_info_138_vecWen;
    rand bit         io_diffCommits_info_138_v0Wen;
    rand bit         io_diffCommits_info_138_vlWen;
    rand bit [5:0]   io_diffCommits_info_139_ldest;
    rand bit [7:0]   io_diffCommits_info_139_pdest;
    rand bit         io_diffCommits_info_139_rfWen;
    rand bit         io_diffCommits_info_139_fpWen;
    rand bit         io_diffCommits_info_139_vecWen;
    rand bit         io_diffCommits_info_139_v0Wen;
    rand bit         io_diffCommits_info_139_vlWen;
    rand bit [5:0]   io_diffCommits_info_140_ldest;
    rand bit [7:0]   io_diffCommits_info_140_pdest;
    rand bit         io_diffCommits_info_140_rfWen;
    rand bit         io_diffCommits_info_140_fpWen;
    rand bit         io_diffCommits_info_140_vecWen;
    rand bit         io_diffCommits_info_140_v0Wen;
    rand bit         io_diffCommits_info_140_vlWen;
    rand bit [5:0]   io_diffCommits_info_141_ldest;
    rand bit [7:0]   io_diffCommits_info_141_pdest;
    rand bit         io_diffCommits_info_141_rfWen;
    rand bit         io_diffCommits_info_141_fpWen;
    rand bit         io_diffCommits_info_141_vecWen;
    rand bit         io_diffCommits_info_141_v0Wen;
    rand bit         io_diffCommits_info_141_vlWen;
    rand bit [5:0]   io_diffCommits_info_142_ldest;
    rand bit [7:0]   io_diffCommits_info_142_pdest;
    rand bit         io_diffCommits_info_142_rfWen;
    rand bit         io_diffCommits_info_142_fpWen;
    rand bit         io_diffCommits_info_142_vecWen;
    rand bit         io_diffCommits_info_142_v0Wen;
    rand bit         io_diffCommits_info_142_vlWen;
    rand bit [5:0]   io_diffCommits_info_143_ldest;
    rand bit [7:0]   io_diffCommits_info_143_pdest;
    rand bit         io_diffCommits_info_143_rfWen;
    rand bit         io_diffCommits_info_143_fpWen;
    rand bit         io_diffCommits_info_143_vecWen;
    rand bit         io_diffCommits_info_143_v0Wen;
    rand bit         io_diffCommits_info_143_vlWen;
    rand bit [5:0]   io_diffCommits_info_144_ldest;
    rand bit [7:0]   io_diffCommits_info_144_pdest;
    rand bit         io_diffCommits_info_144_rfWen;
    rand bit         io_diffCommits_info_144_fpWen;
    rand bit         io_diffCommits_info_144_vecWen;
    rand bit         io_diffCommits_info_144_v0Wen;
    rand bit         io_diffCommits_info_144_vlWen;
    rand bit [5:0]   io_diffCommits_info_145_ldest;
    rand bit [7:0]   io_diffCommits_info_145_pdest;
    rand bit         io_diffCommits_info_145_rfWen;
    rand bit         io_diffCommits_info_145_fpWen;
    rand bit         io_diffCommits_info_145_vecWen;
    rand bit         io_diffCommits_info_145_v0Wen;
    rand bit         io_diffCommits_info_145_vlWen;
    rand bit [5:0]   io_diffCommits_info_146_ldest;
    rand bit [7:0]   io_diffCommits_info_146_pdest;
    rand bit         io_diffCommits_info_146_rfWen;
    rand bit         io_diffCommits_info_146_fpWen;
    rand bit         io_diffCommits_info_146_vecWen;
    rand bit         io_diffCommits_info_146_v0Wen;
    rand bit         io_diffCommits_info_146_vlWen;
    rand bit [5:0]   io_diffCommits_info_147_ldest;
    rand bit [7:0]   io_diffCommits_info_147_pdest;
    rand bit         io_diffCommits_info_147_rfWen;
    rand bit         io_diffCommits_info_147_fpWen;
    rand bit         io_diffCommits_info_147_vecWen;
    rand bit         io_diffCommits_info_147_v0Wen;
    rand bit         io_diffCommits_info_147_vlWen;
    rand bit [5:0]   io_diffCommits_info_148_ldest;
    rand bit [7:0]   io_diffCommits_info_148_pdest;
    rand bit         io_diffCommits_info_148_rfWen;
    rand bit         io_diffCommits_info_148_fpWen;
    rand bit         io_diffCommits_info_148_vecWen;
    rand bit         io_diffCommits_info_148_v0Wen;
    rand bit         io_diffCommits_info_148_vlWen;
    rand bit [5:0]   io_diffCommits_info_149_ldest;
    rand bit [7:0]   io_diffCommits_info_149_pdest;
    rand bit         io_diffCommits_info_149_rfWen;
    rand bit         io_diffCommits_info_149_fpWen;
    rand bit         io_diffCommits_info_149_vecWen;
    rand bit         io_diffCommits_info_149_v0Wen;
    rand bit         io_diffCommits_info_149_vlWen;
    rand bit [5:0]   io_diffCommits_info_150_ldest;
    rand bit [7:0]   io_diffCommits_info_150_pdest;
    rand bit         io_diffCommits_info_150_rfWen;
    rand bit         io_diffCommits_info_150_fpWen;
    rand bit         io_diffCommits_info_150_vecWen;
    rand bit         io_diffCommits_info_150_v0Wen;
    rand bit         io_diffCommits_info_150_vlWen;
    rand bit [5:0]   io_diffCommits_info_151_ldest;
    rand bit [7:0]   io_diffCommits_info_151_pdest;
    rand bit         io_diffCommits_info_151_rfWen;
    rand bit         io_diffCommits_info_151_fpWen;
    rand bit         io_diffCommits_info_151_vecWen;
    rand bit         io_diffCommits_info_151_v0Wen;
    rand bit         io_diffCommits_info_151_vlWen;
    rand bit [5:0]   io_diffCommits_info_152_ldest;
    rand bit [7:0]   io_diffCommits_info_152_pdest;
    rand bit         io_diffCommits_info_152_rfWen;
    rand bit         io_diffCommits_info_152_fpWen;
    rand bit         io_diffCommits_info_152_vecWen;
    rand bit         io_diffCommits_info_152_v0Wen;
    rand bit         io_diffCommits_info_152_vlWen;
    rand bit [5:0]   io_diffCommits_info_153_ldest;
    rand bit [7:0]   io_diffCommits_info_153_pdest;
    rand bit         io_diffCommits_info_153_rfWen;
    rand bit         io_diffCommits_info_153_fpWen;
    rand bit         io_diffCommits_info_153_vecWen;
    rand bit         io_diffCommits_info_153_v0Wen;
    rand bit         io_diffCommits_info_153_vlWen;
    rand bit [5:0]   io_diffCommits_info_154_ldest;
    rand bit [7:0]   io_diffCommits_info_154_pdest;
    rand bit         io_diffCommits_info_154_rfWen;
    rand bit         io_diffCommits_info_154_fpWen;
    rand bit         io_diffCommits_info_154_vecWen;
    rand bit         io_diffCommits_info_154_v0Wen;
    rand bit         io_diffCommits_info_154_vlWen;
    rand bit [5:0]   io_diffCommits_info_155_ldest;
    rand bit [7:0]   io_diffCommits_info_155_pdest;
    rand bit         io_diffCommits_info_155_rfWen;
    rand bit         io_diffCommits_info_155_fpWen;
    rand bit         io_diffCommits_info_155_vecWen;
    rand bit         io_diffCommits_info_155_v0Wen;
    rand bit         io_diffCommits_info_155_vlWen;
    rand bit [5:0]   io_diffCommits_info_156_ldest;
    rand bit [7:0]   io_diffCommits_info_156_pdest;
    rand bit         io_diffCommits_info_156_rfWen;
    rand bit         io_diffCommits_info_156_fpWen;
    rand bit         io_diffCommits_info_156_vecWen;
    rand bit         io_diffCommits_info_156_v0Wen;
    rand bit         io_diffCommits_info_156_vlWen;
    rand bit [5:0]   io_diffCommits_info_157_ldest;
    rand bit [7:0]   io_diffCommits_info_157_pdest;
    rand bit         io_diffCommits_info_157_rfWen;
    rand bit         io_diffCommits_info_157_fpWen;
    rand bit         io_diffCommits_info_157_vecWen;
    rand bit         io_diffCommits_info_157_v0Wen;
    rand bit         io_diffCommits_info_157_vlWen;
    rand bit [5:0]   io_diffCommits_info_158_ldest;
    rand bit [7:0]   io_diffCommits_info_158_pdest;
    rand bit         io_diffCommits_info_158_rfWen;
    rand bit         io_diffCommits_info_158_fpWen;
    rand bit         io_diffCommits_info_158_vecWen;
    rand bit         io_diffCommits_info_158_v0Wen;
    rand bit         io_diffCommits_info_158_vlWen;
    rand bit [5:0]   io_diffCommits_info_159_ldest;
    rand bit [7:0]   io_diffCommits_info_159_pdest;
    rand bit         io_diffCommits_info_159_rfWen;
    rand bit         io_diffCommits_info_159_fpWen;
    rand bit         io_diffCommits_info_159_vecWen;
    rand bit         io_diffCommits_info_159_v0Wen;
    rand bit         io_diffCommits_info_159_vlWen;
    rand bit [5:0]   io_diffCommits_info_160_ldest;
    rand bit [7:0]   io_diffCommits_info_160_pdest;
    rand bit         io_diffCommits_info_160_rfWen;
    rand bit         io_diffCommits_info_160_fpWen;
    rand bit         io_diffCommits_info_160_vecWen;
    rand bit         io_diffCommits_info_160_v0Wen;
    rand bit         io_diffCommits_info_160_vlWen;
    rand bit [5:0]   io_diffCommits_info_161_ldest;
    rand bit [7:0]   io_diffCommits_info_161_pdest;
    rand bit         io_diffCommits_info_161_rfWen;
    rand bit         io_diffCommits_info_161_fpWen;
    rand bit         io_diffCommits_info_161_vecWen;
    rand bit         io_diffCommits_info_161_v0Wen;
    rand bit         io_diffCommits_info_161_vlWen;
    rand bit [5:0]   io_diffCommits_info_162_ldest;
    rand bit [7:0]   io_diffCommits_info_162_pdest;
    rand bit         io_diffCommits_info_162_rfWen;
    rand bit         io_diffCommits_info_162_fpWen;
    rand bit         io_diffCommits_info_162_vecWen;
    rand bit         io_diffCommits_info_162_v0Wen;
    rand bit         io_diffCommits_info_162_vlWen;
    rand bit [5:0]   io_diffCommits_info_163_ldest;
    rand bit [7:0]   io_diffCommits_info_163_pdest;
    rand bit         io_diffCommits_info_163_rfWen;
    rand bit         io_diffCommits_info_163_fpWen;
    rand bit         io_diffCommits_info_163_vecWen;
    rand bit         io_diffCommits_info_163_v0Wen;
    rand bit         io_diffCommits_info_163_vlWen;
    rand bit [5:0]   io_diffCommits_info_164_ldest;
    rand bit [7:0]   io_diffCommits_info_164_pdest;
    rand bit         io_diffCommits_info_164_rfWen;
    rand bit         io_diffCommits_info_164_fpWen;
    rand bit         io_diffCommits_info_164_vecWen;
    rand bit         io_diffCommits_info_164_v0Wen;
    rand bit         io_diffCommits_info_164_vlWen;
    rand bit [5:0]   io_diffCommits_info_165_ldest;
    rand bit [7:0]   io_diffCommits_info_165_pdest;
    rand bit         io_diffCommits_info_165_rfWen;
    rand bit         io_diffCommits_info_165_fpWen;
    rand bit         io_diffCommits_info_165_vecWen;
    rand bit         io_diffCommits_info_165_v0Wen;
    rand bit         io_diffCommits_info_165_vlWen;
    rand bit [5:0]   io_diffCommits_info_166_ldest;
    rand bit [7:0]   io_diffCommits_info_166_pdest;
    rand bit         io_diffCommits_info_166_rfWen;
    rand bit         io_diffCommits_info_166_fpWen;
    rand bit         io_diffCommits_info_166_vecWen;
    rand bit         io_diffCommits_info_166_v0Wen;
    rand bit         io_diffCommits_info_166_vlWen;
    rand bit [5:0]   io_diffCommits_info_167_ldest;
    rand bit [7:0]   io_diffCommits_info_167_pdest;
    rand bit         io_diffCommits_info_167_rfWen;
    rand bit         io_diffCommits_info_167_fpWen;
    rand bit         io_diffCommits_info_167_vecWen;
    rand bit         io_diffCommits_info_167_v0Wen;
    rand bit         io_diffCommits_info_167_vlWen;
    rand bit [5:0]   io_diffCommits_info_168_ldest;
    rand bit [7:0]   io_diffCommits_info_168_pdest;
    rand bit         io_diffCommits_info_168_rfWen;
    rand bit         io_diffCommits_info_168_fpWen;
    rand bit         io_diffCommits_info_168_vecWen;
    rand bit         io_diffCommits_info_168_v0Wen;
    rand bit         io_diffCommits_info_168_vlWen;
    rand bit [5:0]   io_diffCommits_info_169_ldest;
    rand bit [7:0]   io_diffCommits_info_169_pdest;
    rand bit         io_diffCommits_info_169_rfWen;
    rand bit         io_diffCommits_info_169_fpWen;
    rand bit         io_diffCommits_info_169_vecWen;
    rand bit         io_diffCommits_info_169_v0Wen;
    rand bit         io_diffCommits_info_169_vlWen;
    rand bit [5:0]   io_diffCommits_info_170_ldest;
    rand bit [7:0]   io_diffCommits_info_170_pdest;
    rand bit         io_diffCommits_info_170_rfWen;
    rand bit         io_diffCommits_info_170_fpWen;
    rand bit         io_diffCommits_info_170_vecWen;
    rand bit         io_diffCommits_info_170_v0Wen;
    rand bit         io_diffCommits_info_170_vlWen;
    rand bit [5:0]   io_diffCommits_info_171_ldest;
    rand bit [7:0]   io_diffCommits_info_171_pdest;
    rand bit         io_diffCommits_info_171_rfWen;
    rand bit         io_diffCommits_info_171_fpWen;
    rand bit         io_diffCommits_info_171_vecWen;
    rand bit         io_diffCommits_info_171_v0Wen;
    rand bit         io_diffCommits_info_171_vlWen;
    rand bit [5:0]   io_diffCommits_info_172_ldest;
    rand bit [7:0]   io_diffCommits_info_172_pdest;
    rand bit         io_diffCommits_info_172_rfWen;
    rand bit         io_diffCommits_info_172_fpWen;
    rand bit         io_diffCommits_info_172_vecWen;
    rand bit         io_diffCommits_info_172_v0Wen;
    rand bit         io_diffCommits_info_172_vlWen;
    rand bit [5:0]   io_diffCommits_info_173_ldest;
    rand bit [7:0]   io_diffCommits_info_173_pdest;
    rand bit         io_diffCommits_info_173_rfWen;
    rand bit         io_diffCommits_info_173_fpWen;
    rand bit         io_diffCommits_info_173_vecWen;
    rand bit         io_diffCommits_info_173_v0Wen;
    rand bit         io_diffCommits_info_173_vlWen;
    rand bit [5:0]   io_diffCommits_info_174_ldest;
    rand bit [7:0]   io_diffCommits_info_174_pdest;
    rand bit         io_diffCommits_info_174_rfWen;
    rand bit         io_diffCommits_info_174_fpWen;
    rand bit         io_diffCommits_info_174_vecWen;
    rand bit         io_diffCommits_info_174_v0Wen;
    rand bit         io_diffCommits_info_174_vlWen;
    rand bit [5:0]   io_diffCommits_info_175_ldest;
    rand bit [7:0]   io_diffCommits_info_175_pdest;
    rand bit         io_diffCommits_info_175_rfWen;
    rand bit         io_diffCommits_info_175_fpWen;
    rand bit         io_diffCommits_info_175_vecWen;
    rand bit         io_diffCommits_info_175_v0Wen;
    rand bit         io_diffCommits_info_175_vlWen;
    rand bit [5:0]   io_diffCommits_info_176_ldest;
    rand bit [7:0]   io_diffCommits_info_176_pdest;
    rand bit         io_diffCommits_info_176_rfWen;
    rand bit         io_diffCommits_info_176_fpWen;
    rand bit         io_diffCommits_info_176_vecWen;
    rand bit         io_diffCommits_info_176_v0Wen;
    rand bit         io_diffCommits_info_176_vlWen;
    rand bit [5:0]   io_diffCommits_info_177_ldest;
    rand bit [7:0]   io_diffCommits_info_177_pdest;
    rand bit         io_diffCommits_info_177_rfWen;
    rand bit         io_diffCommits_info_177_fpWen;
    rand bit         io_diffCommits_info_177_vecWen;
    rand bit         io_diffCommits_info_177_v0Wen;
    rand bit         io_diffCommits_info_177_vlWen;
    rand bit [5:0]   io_diffCommits_info_178_ldest;
    rand bit [7:0]   io_diffCommits_info_178_pdest;
    rand bit         io_diffCommits_info_178_rfWen;
    rand bit         io_diffCommits_info_178_fpWen;
    rand bit         io_diffCommits_info_178_vecWen;
    rand bit         io_diffCommits_info_178_v0Wen;
    rand bit         io_diffCommits_info_178_vlWen;
    rand bit [5:0]   io_diffCommits_info_179_ldest;
    rand bit [7:0]   io_diffCommits_info_179_pdest;
    rand bit         io_diffCommits_info_179_rfWen;
    rand bit         io_diffCommits_info_179_fpWen;
    rand bit         io_diffCommits_info_179_vecWen;
    rand bit         io_diffCommits_info_179_v0Wen;
    rand bit         io_diffCommits_info_179_vlWen;
    rand bit [5:0]   io_diffCommits_info_180_ldest;
    rand bit [7:0]   io_diffCommits_info_180_pdest;
    rand bit         io_diffCommits_info_180_rfWen;
    rand bit         io_diffCommits_info_180_fpWen;
    rand bit         io_diffCommits_info_180_vecWen;
    rand bit         io_diffCommits_info_180_v0Wen;
    rand bit         io_diffCommits_info_180_vlWen;
    rand bit [5:0]   io_diffCommits_info_181_ldest;
    rand bit [7:0]   io_diffCommits_info_181_pdest;
    rand bit         io_diffCommits_info_181_rfWen;
    rand bit         io_diffCommits_info_181_fpWen;
    rand bit         io_diffCommits_info_181_vecWen;
    rand bit         io_diffCommits_info_181_v0Wen;
    rand bit         io_diffCommits_info_181_vlWen;
    rand bit [5:0]   io_diffCommits_info_182_ldest;
    rand bit [7:0]   io_diffCommits_info_182_pdest;
    rand bit         io_diffCommits_info_182_rfWen;
    rand bit         io_diffCommits_info_182_fpWen;
    rand bit         io_diffCommits_info_182_vecWen;
    rand bit         io_diffCommits_info_182_v0Wen;
    rand bit         io_diffCommits_info_182_vlWen;
    rand bit [5:0]   io_diffCommits_info_183_ldest;
    rand bit [7:0]   io_diffCommits_info_183_pdest;
    rand bit         io_diffCommits_info_183_rfWen;
    rand bit         io_diffCommits_info_183_fpWen;
    rand bit         io_diffCommits_info_183_vecWen;
    rand bit         io_diffCommits_info_183_v0Wen;
    rand bit         io_diffCommits_info_183_vlWen;
    rand bit [5:0]   io_diffCommits_info_184_ldest;
    rand bit [7:0]   io_diffCommits_info_184_pdest;
    rand bit         io_diffCommits_info_184_rfWen;
    rand bit         io_diffCommits_info_184_fpWen;
    rand bit         io_diffCommits_info_184_vecWen;
    rand bit         io_diffCommits_info_184_v0Wen;
    rand bit         io_diffCommits_info_184_vlWen;
    rand bit [5:0]   io_diffCommits_info_185_ldest;
    rand bit [7:0]   io_diffCommits_info_185_pdest;
    rand bit         io_diffCommits_info_185_rfWen;
    rand bit         io_diffCommits_info_185_fpWen;
    rand bit         io_diffCommits_info_185_vecWen;
    rand bit         io_diffCommits_info_185_v0Wen;
    rand bit         io_diffCommits_info_185_vlWen;
    rand bit [5:0]   io_diffCommits_info_186_ldest;
    rand bit [7:0]   io_diffCommits_info_186_pdest;
    rand bit         io_diffCommits_info_186_rfWen;
    rand bit         io_diffCommits_info_186_fpWen;
    rand bit         io_diffCommits_info_186_vecWen;
    rand bit         io_diffCommits_info_186_v0Wen;
    rand bit         io_diffCommits_info_186_vlWen;
    rand bit [5:0]   io_diffCommits_info_187_ldest;
    rand bit [7:0]   io_diffCommits_info_187_pdest;
    rand bit         io_diffCommits_info_187_rfWen;
    rand bit         io_diffCommits_info_187_fpWen;
    rand bit         io_diffCommits_info_187_vecWen;
    rand bit         io_diffCommits_info_187_v0Wen;
    rand bit         io_diffCommits_info_187_vlWen;
    rand bit [5:0]   io_diffCommits_info_188_ldest;
    rand bit [7:0]   io_diffCommits_info_188_pdest;
    rand bit         io_diffCommits_info_188_rfWen;
    rand bit         io_diffCommits_info_188_fpWen;
    rand bit         io_diffCommits_info_188_vecWen;
    rand bit         io_diffCommits_info_188_v0Wen;
    rand bit         io_diffCommits_info_188_vlWen;
    rand bit [5:0]   io_diffCommits_info_189_ldest;
    rand bit [7:0]   io_diffCommits_info_189_pdest;
    rand bit         io_diffCommits_info_189_rfWen;
    rand bit         io_diffCommits_info_189_fpWen;
    rand bit         io_diffCommits_info_189_vecWen;
    rand bit         io_diffCommits_info_189_v0Wen;
    rand bit         io_diffCommits_info_189_vlWen;
    rand bit [5:0]   io_diffCommits_info_190_ldest;
    rand bit [7:0]   io_diffCommits_info_190_pdest;
    rand bit         io_diffCommits_info_190_rfWen;
    rand bit         io_diffCommits_info_190_fpWen;
    rand bit         io_diffCommits_info_190_vecWen;
    rand bit         io_diffCommits_info_190_v0Wen;
    rand bit         io_diffCommits_info_190_vlWen;
    rand bit [5:0]   io_diffCommits_info_191_ldest;
    rand bit [7:0]   io_diffCommits_info_191_pdest;
    rand bit         io_diffCommits_info_191_rfWen;
    rand bit         io_diffCommits_info_191_fpWen;
    rand bit         io_diffCommits_info_191_vecWen;
    rand bit         io_diffCommits_info_191_v0Wen;
    rand bit         io_diffCommits_info_191_vlWen;
    rand bit [5:0]   io_diffCommits_info_192_ldest;
    rand bit [7:0]   io_diffCommits_info_192_pdest;
    rand bit         io_diffCommits_info_192_rfWen;
    rand bit         io_diffCommits_info_192_fpWen;
    rand bit         io_diffCommits_info_192_vecWen;
    rand bit         io_diffCommits_info_192_v0Wen;
    rand bit         io_diffCommits_info_192_vlWen;
    rand bit [5:0]   io_diffCommits_info_193_ldest;
    rand bit [7:0]   io_diffCommits_info_193_pdest;
    rand bit         io_diffCommits_info_193_rfWen;
    rand bit         io_diffCommits_info_193_fpWen;
    rand bit         io_diffCommits_info_193_vecWen;
    rand bit         io_diffCommits_info_193_v0Wen;
    rand bit         io_diffCommits_info_193_vlWen;
    rand bit [5:0]   io_diffCommits_info_194_ldest;
    rand bit [7:0]   io_diffCommits_info_194_pdest;
    rand bit         io_diffCommits_info_194_rfWen;
    rand bit         io_diffCommits_info_194_fpWen;
    rand bit         io_diffCommits_info_194_vecWen;
    rand bit         io_diffCommits_info_194_v0Wen;
    rand bit         io_diffCommits_info_194_vlWen;
    rand bit [5:0]   io_diffCommits_info_195_ldest;
    rand bit [7:0]   io_diffCommits_info_195_pdest;
    rand bit         io_diffCommits_info_195_rfWen;
    rand bit         io_diffCommits_info_195_fpWen;
    rand bit         io_diffCommits_info_195_vecWen;
    rand bit         io_diffCommits_info_195_v0Wen;
    rand bit         io_diffCommits_info_195_vlWen;
    rand bit [5:0]   io_diffCommits_info_196_ldest;
    rand bit [7:0]   io_diffCommits_info_196_pdest;
    rand bit         io_diffCommits_info_196_rfWen;
    rand bit         io_diffCommits_info_196_fpWen;
    rand bit         io_diffCommits_info_196_vecWen;
    rand bit         io_diffCommits_info_196_v0Wen;
    rand bit         io_diffCommits_info_196_vlWen;
    rand bit [5:0]   io_diffCommits_info_197_ldest;
    rand bit [7:0]   io_diffCommits_info_197_pdest;
    rand bit         io_diffCommits_info_197_rfWen;
    rand bit         io_diffCommits_info_197_fpWen;
    rand bit         io_diffCommits_info_197_vecWen;
    rand bit         io_diffCommits_info_197_v0Wen;
    rand bit         io_diffCommits_info_197_vlWen;
    rand bit [5:0]   io_diffCommits_info_198_ldest;
    rand bit [7:0]   io_diffCommits_info_198_pdest;
    rand bit         io_diffCommits_info_198_rfWen;
    rand bit         io_diffCommits_info_198_fpWen;
    rand bit         io_diffCommits_info_198_vecWen;
    rand bit         io_diffCommits_info_198_v0Wen;
    rand bit         io_diffCommits_info_198_vlWen;
    rand bit [5:0]   io_diffCommits_info_199_ldest;
    rand bit [7:0]   io_diffCommits_info_199_pdest;
    rand bit         io_diffCommits_info_199_rfWen;
    rand bit         io_diffCommits_info_199_fpWen;
    rand bit         io_diffCommits_info_199_vecWen;
    rand bit         io_diffCommits_info_199_v0Wen;
    rand bit         io_diffCommits_info_199_vlWen;
    rand bit [5:0]   io_diffCommits_info_200_ldest;
    rand bit [7:0]   io_diffCommits_info_200_pdest;
    rand bit         io_diffCommits_info_200_rfWen;
    rand bit         io_diffCommits_info_200_fpWen;
    rand bit         io_diffCommits_info_200_vecWen;
    rand bit         io_diffCommits_info_200_v0Wen;
    rand bit         io_diffCommits_info_200_vlWen;
    rand bit [5:0]   io_diffCommits_info_201_ldest;
    rand bit [7:0]   io_diffCommits_info_201_pdest;
    rand bit         io_diffCommits_info_201_rfWen;
    rand bit         io_diffCommits_info_201_fpWen;
    rand bit         io_diffCommits_info_201_vecWen;
    rand bit         io_diffCommits_info_201_v0Wen;
    rand bit         io_diffCommits_info_201_vlWen;
    rand bit [5:0]   io_diffCommits_info_202_ldest;
    rand bit [7:0]   io_diffCommits_info_202_pdest;
    rand bit         io_diffCommits_info_202_rfWen;
    rand bit         io_diffCommits_info_202_fpWen;
    rand bit         io_diffCommits_info_202_vecWen;
    rand bit         io_diffCommits_info_202_v0Wen;
    rand bit         io_diffCommits_info_202_vlWen;
    rand bit [5:0]   io_diffCommits_info_203_ldest;
    rand bit [7:0]   io_diffCommits_info_203_pdest;
    rand bit         io_diffCommits_info_203_rfWen;
    rand bit         io_diffCommits_info_203_fpWen;
    rand bit         io_diffCommits_info_203_vecWen;
    rand bit         io_diffCommits_info_203_v0Wen;
    rand bit         io_diffCommits_info_203_vlWen;
    rand bit [5:0]   io_diffCommits_info_204_ldest;
    rand bit [7:0]   io_diffCommits_info_204_pdest;
    rand bit         io_diffCommits_info_204_rfWen;
    rand bit         io_diffCommits_info_204_fpWen;
    rand bit         io_diffCommits_info_204_vecWen;
    rand bit         io_diffCommits_info_204_v0Wen;
    rand bit         io_diffCommits_info_204_vlWen;
    rand bit [5:0]   io_diffCommits_info_205_ldest;
    rand bit [7:0]   io_diffCommits_info_205_pdest;
    rand bit         io_diffCommits_info_205_rfWen;
    rand bit         io_diffCommits_info_205_fpWen;
    rand bit         io_diffCommits_info_205_vecWen;
    rand bit         io_diffCommits_info_205_v0Wen;
    rand bit         io_diffCommits_info_205_vlWen;
    rand bit [5:0]   io_diffCommits_info_206_ldest;
    rand bit [7:0]   io_diffCommits_info_206_pdest;
    rand bit         io_diffCommits_info_206_rfWen;
    rand bit         io_diffCommits_info_206_fpWen;
    rand bit         io_diffCommits_info_206_vecWen;
    rand bit         io_diffCommits_info_206_v0Wen;
    rand bit         io_diffCommits_info_206_vlWen;
    rand bit [5:0]   io_diffCommits_info_207_ldest;
    rand bit [7:0]   io_diffCommits_info_207_pdest;
    rand bit         io_diffCommits_info_207_rfWen;
    rand bit         io_diffCommits_info_207_fpWen;
    rand bit         io_diffCommits_info_207_vecWen;
    rand bit         io_diffCommits_info_207_v0Wen;
    rand bit         io_diffCommits_info_207_vlWen;
    rand bit [5:0]   io_diffCommits_info_208_ldest;
    rand bit [7:0]   io_diffCommits_info_208_pdest;
    rand bit         io_diffCommits_info_208_rfWen;
    rand bit         io_diffCommits_info_208_fpWen;
    rand bit         io_diffCommits_info_208_vecWen;
    rand bit         io_diffCommits_info_208_v0Wen;
    rand bit         io_diffCommits_info_208_vlWen;
    rand bit [5:0]   io_diffCommits_info_209_ldest;
    rand bit [7:0]   io_diffCommits_info_209_pdest;
    rand bit         io_diffCommits_info_209_rfWen;
    rand bit         io_diffCommits_info_209_fpWen;
    rand bit         io_diffCommits_info_209_vecWen;
    rand bit         io_diffCommits_info_209_v0Wen;
    rand bit         io_diffCommits_info_209_vlWen;
    rand bit [5:0]   io_diffCommits_info_210_ldest;
    rand bit [7:0]   io_diffCommits_info_210_pdest;
    rand bit         io_diffCommits_info_210_rfWen;
    rand bit         io_diffCommits_info_210_fpWen;
    rand bit         io_diffCommits_info_210_vecWen;
    rand bit         io_diffCommits_info_210_v0Wen;
    rand bit         io_diffCommits_info_210_vlWen;
    rand bit [5:0]   io_diffCommits_info_211_ldest;
    rand bit [7:0]   io_diffCommits_info_211_pdest;
    rand bit         io_diffCommits_info_211_rfWen;
    rand bit         io_diffCommits_info_211_fpWen;
    rand bit         io_diffCommits_info_211_vecWen;
    rand bit         io_diffCommits_info_211_v0Wen;
    rand bit         io_diffCommits_info_211_vlWen;
    rand bit [5:0]   io_diffCommits_info_212_ldest;
    rand bit [7:0]   io_diffCommits_info_212_pdest;
    rand bit         io_diffCommits_info_212_rfWen;
    rand bit         io_diffCommits_info_212_fpWen;
    rand bit         io_diffCommits_info_212_vecWen;
    rand bit         io_diffCommits_info_212_v0Wen;
    rand bit         io_diffCommits_info_212_vlWen;
    rand bit [5:0]   io_diffCommits_info_213_ldest;
    rand bit [7:0]   io_diffCommits_info_213_pdest;
    rand bit         io_diffCommits_info_213_rfWen;
    rand bit         io_diffCommits_info_213_fpWen;
    rand bit         io_diffCommits_info_213_vecWen;
    rand bit         io_diffCommits_info_213_v0Wen;
    rand bit         io_diffCommits_info_213_vlWen;
    rand bit [5:0]   io_diffCommits_info_214_ldest;
    rand bit [7:0]   io_diffCommits_info_214_pdest;
    rand bit         io_diffCommits_info_214_rfWen;
    rand bit         io_diffCommits_info_214_fpWen;
    rand bit         io_diffCommits_info_214_vecWen;
    rand bit         io_diffCommits_info_214_v0Wen;
    rand bit         io_diffCommits_info_214_vlWen;
    rand bit [5:0]   io_diffCommits_info_215_ldest;
    rand bit [7:0]   io_diffCommits_info_215_pdest;
    rand bit         io_diffCommits_info_215_rfWen;
    rand bit         io_diffCommits_info_215_fpWen;
    rand bit         io_diffCommits_info_215_vecWen;
    rand bit         io_diffCommits_info_215_v0Wen;
    rand bit         io_diffCommits_info_215_vlWen;
    rand bit [5:0]   io_diffCommits_info_216_ldest;
    rand bit [7:0]   io_diffCommits_info_216_pdest;
    rand bit         io_diffCommits_info_216_rfWen;
    rand bit         io_diffCommits_info_216_fpWen;
    rand bit         io_diffCommits_info_216_vecWen;
    rand bit         io_diffCommits_info_216_v0Wen;
    rand bit         io_diffCommits_info_216_vlWen;
    rand bit [5:0]   io_diffCommits_info_217_ldest;
    rand bit [7:0]   io_diffCommits_info_217_pdest;
    rand bit         io_diffCommits_info_217_rfWen;
    rand bit         io_diffCommits_info_217_fpWen;
    rand bit         io_diffCommits_info_217_vecWen;
    rand bit         io_diffCommits_info_217_v0Wen;
    rand bit         io_diffCommits_info_217_vlWen;
    rand bit [5:0]   io_diffCommits_info_218_ldest;
    rand bit [7:0]   io_diffCommits_info_218_pdest;
    rand bit         io_diffCommits_info_218_rfWen;
    rand bit         io_diffCommits_info_218_fpWen;
    rand bit         io_diffCommits_info_218_vecWen;
    rand bit         io_diffCommits_info_218_v0Wen;
    rand bit         io_diffCommits_info_218_vlWen;
    rand bit [5:0]   io_diffCommits_info_219_ldest;
    rand bit [7:0]   io_diffCommits_info_219_pdest;
    rand bit         io_diffCommits_info_219_rfWen;
    rand bit         io_diffCommits_info_219_fpWen;
    rand bit         io_diffCommits_info_219_vecWen;
    rand bit         io_diffCommits_info_219_v0Wen;
    rand bit         io_diffCommits_info_219_vlWen;
    rand bit [5:0]   io_diffCommits_info_220_ldest;
    rand bit [7:0]   io_diffCommits_info_220_pdest;
    rand bit         io_diffCommits_info_220_rfWen;
    rand bit         io_diffCommits_info_220_fpWen;
    rand bit         io_diffCommits_info_220_vecWen;
    rand bit         io_diffCommits_info_220_v0Wen;
    rand bit         io_diffCommits_info_220_vlWen;
    rand bit [5:0]   io_diffCommits_info_221_ldest;
    rand bit [7:0]   io_diffCommits_info_221_pdest;
    rand bit         io_diffCommits_info_221_rfWen;
    rand bit         io_diffCommits_info_221_fpWen;
    rand bit         io_diffCommits_info_221_vecWen;
    rand bit         io_diffCommits_info_221_v0Wen;
    rand bit         io_diffCommits_info_221_vlWen;
    rand bit [5:0]   io_diffCommits_info_222_ldest;
    rand bit [7:0]   io_diffCommits_info_222_pdest;
    rand bit         io_diffCommits_info_222_rfWen;
    rand bit         io_diffCommits_info_222_fpWen;
    rand bit         io_diffCommits_info_222_vecWen;
    rand bit         io_diffCommits_info_222_v0Wen;
    rand bit         io_diffCommits_info_222_vlWen;
    rand bit [5:0]   io_diffCommits_info_223_ldest;
    rand bit [7:0]   io_diffCommits_info_223_pdest;
    rand bit         io_diffCommits_info_223_rfWen;
    rand bit         io_diffCommits_info_223_fpWen;
    rand bit         io_diffCommits_info_223_vecWen;
    rand bit         io_diffCommits_info_223_v0Wen;
    rand bit         io_diffCommits_info_223_vlWen;
    rand bit [5:0]   io_diffCommits_info_224_ldest;
    rand bit [7:0]   io_diffCommits_info_224_pdest;
    rand bit         io_diffCommits_info_224_rfWen;
    rand bit         io_diffCommits_info_224_fpWen;
    rand bit         io_diffCommits_info_224_vecWen;
    rand bit         io_diffCommits_info_224_v0Wen;
    rand bit         io_diffCommits_info_224_vlWen;
    rand bit [5:0]   io_diffCommits_info_225_ldest;
    rand bit [7:0]   io_diffCommits_info_225_pdest;
    rand bit         io_diffCommits_info_225_rfWen;
    rand bit         io_diffCommits_info_225_fpWen;
    rand bit         io_diffCommits_info_225_vecWen;
    rand bit         io_diffCommits_info_225_v0Wen;
    rand bit         io_diffCommits_info_225_vlWen;
    rand bit [5:0]   io_diffCommits_info_226_ldest;
    rand bit [7:0]   io_diffCommits_info_226_pdest;
    rand bit         io_diffCommits_info_226_rfWen;
    rand bit         io_diffCommits_info_226_fpWen;
    rand bit         io_diffCommits_info_226_vecWen;
    rand bit         io_diffCommits_info_226_v0Wen;
    rand bit         io_diffCommits_info_226_vlWen;
    rand bit [5:0]   io_diffCommits_info_227_ldest;
    rand bit [7:0]   io_diffCommits_info_227_pdest;
    rand bit         io_diffCommits_info_227_rfWen;
    rand bit         io_diffCommits_info_227_fpWen;
    rand bit         io_diffCommits_info_227_vecWen;
    rand bit         io_diffCommits_info_227_v0Wen;
    rand bit         io_diffCommits_info_227_vlWen;
    rand bit [5:0]   io_diffCommits_info_228_ldest;
    rand bit [7:0]   io_diffCommits_info_228_pdest;
    rand bit         io_diffCommits_info_228_rfWen;
    rand bit         io_diffCommits_info_228_fpWen;
    rand bit         io_diffCommits_info_228_vecWen;
    rand bit         io_diffCommits_info_228_v0Wen;
    rand bit         io_diffCommits_info_228_vlWen;
    rand bit [5:0]   io_diffCommits_info_229_ldest;
    rand bit [7:0]   io_diffCommits_info_229_pdest;
    rand bit         io_diffCommits_info_229_rfWen;
    rand bit         io_diffCommits_info_229_fpWen;
    rand bit         io_diffCommits_info_229_vecWen;
    rand bit         io_diffCommits_info_229_v0Wen;
    rand bit         io_diffCommits_info_229_vlWen;
    rand bit [5:0]   io_diffCommits_info_230_ldest;
    rand bit [7:0]   io_diffCommits_info_230_pdest;
    rand bit         io_diffCommits_info_230_rfWen;
    rand bit         io_diffCommits_info_230_fpWen;
    rand bit         io_diffCommits_info_230_vecWen;
    rand bit         io_diffCommits_info_230_v0Wen;
    rand bit         io_diffCommits_info_230_vlWen;
    rand bit [5:0]   io_diffCommits_info_231_ldest;
    rand bit [7:0]   io_diffCommits_info_231_pdest;
    rand bit         io_diffCommits_info_231_rfWen;
    rand bit         io_diffCommits_info_231_fpWen;
    rand bit         io_diffCommits_info_231_vecWen;
    rand bit         io_diffCommits_info_231_v0Wen;
    rand bit         io_diffCommits_info_231_vlWen;
    rand bit [5:0]   io_diffCommits_info_232_ldest;
    rand bit [7:0]   io_diffCommits_info_232_pdest;
    rand bit         io_diffCommits_info_232_rfWen;
    rand bit         io_diffCommits_info_232_fpWen;
    rand bit         io_diffCommits_info_232_vecWen;
    rand bit         io_diffCommits_info_232_v0Wen;
    rand bit         io_diffCommits_info_232_vlWen;
    rand bit [5:0]   io_diffCommits_info_233_ldest;
    rand bit [7:0]   io_diffCommits_info_233_pdest;
    rand bit         io_diffCommits_info_233_rfWen;
    rand bit         io_diffCommits_info_233_fpWen;
    rand bit         io_diffCommits_info_233_vecWen;
    rand bit         io_diffCommits_info_233_v0Wen;
    rand bit         io_diffCommits_info_233_vlWen;
    rand bit [5:0]   io_diffCommits_info_234_ldest;
    rand bit [7:0]   io_diffCommits_info_234_pdest;
    rand bit         io_diffCommits_info_234_rfWen;
    rand bit         io_diffCommits_info_234_fpWen;
    rand bit         io_diffCommits_info_234_vecWen;
    rand bit         io_diffCommits_info_234_v0Wen;
    rand bit         io_diffCommits_info_234_vlWen;
    rand bit [5:0]   io_diffCommits_info_235_ldest;
    rand bit [7:0]   io_diffCommits_info_235_pdest;
    rand bit         io_diffCommits_info_235_rfWen;
    rand bit         io_diffCommits_info_235_fpWen;
    rand bit         io_diffCommits_info_235_vecWen;
    rand bit         io_diffCommits_info_235_v0Wen;
    rand bit         io_diffCommits_info_235_vlWen;
    rand bit [5:0]   io_diffCommits_info_236_ldest;
    rand bit [7:0]   io_diffCommits_info_236_pdest;
    rand bit         io_diffCommits_info_236_rfWen;
    rand bit         io_diffCommits_info_236_fpWen;
    rand bit         io_diffCommits_info_236_vecWen;
    rand bit         io_diffCommits_info_236_v0Wen;
    rand bit         io_diffCommits_info_236_vlWen;
    rand bit [5:0]   io_diffCommits_info_237_ldest;
    rand bit [7:0]   io_diffCommits_info_237_pdest;
    rand bit         io_diffCommits_info_237_rfWen;
    rand bit         io_diffCommits_info_237_fpWen;
    rand bit         io_diffCommits_info_237_vecWen;
    rand bit         io_diffCommits_info_237_v0Wen;
    rand bit         io_diffCommits_info_237_vlWen;
    rand bit [5:0]   io_diffCommits_info_238_ldest;
    rand bit [7:0]   io_diffCommits_info_238_pdest;
    rand bit         io_diffCommits_info_238_rfWen;
    rand bit         io_diffCommits_info_238_fpWen;
    rand bit         io_diffCommits_info_238_vecWen;
    rand bit         io_diffCommits_info_238_v0Wen;
    rand bit         io_diffCommits_info_238_vlWen;
    rand bit [5:0]   io_diffCommits_info_239_ldest;
    rand bit [7:0]   io_diffCommits_info_239_pdest;
    rand bit         io_diffCommits_info_239_rfWen;
    rand bit         io_diffCommits_info_239_fpWen;
    rand bit         io_diffCommits_info_239_vecWen;
    rand bit         io_diffCommits_info_239_v0Wen;
    rand bit         io_diffCommits_info_239_vlWen;
    rand bit [5:0]   io_diffCommits_info_240_ldest;
    rand bit [7:0]   io_diffCommits_info_240_pdest;
    rand bit         io_diffCommits_info_240_rfWen;
    rand bit         io_diffCommits_info_240_fpWen;
    rand bit         io_diffCommits_info_240_vecWen;
    rand bit         io_diffCommits_info_240_v0Wen;
    rand bit         io_diffCommits_info_240_vlWen;
    rand bit [5:0]   io_diffCommits_info_241_ldest;
    rand bit [7:0]   io_diffCommits_info_241_pdest;
    rand bit         io_diffCommits_info_241_rfWen;
    rand bit         io_diffCommits_info_241_fpWen;
    rand bit         io_diffCommits_info_241_vecWen;
    rand bit         io_diffCommits_info_241_v0Wen;
    rand bit         io_diffCommits_info_241_vlWen;
    rand bit [5:0]   io_diffCommits_info_242_ldest;
    rand bit [7:0]   io_diffCommits_info_242_pdest;
    rand bit         io_diffCommits_info_242_rfWen;
    rand bit         io_diffCommits_info_242_fpWen;
    rand bit         io_diffCommits_info_242_vecWen;
    rand bit         io_diffCommits_info_242_v0Wen;
    rand bit         io_diffCommits_info_242_vlWen;
    rand bit [5:0]   io_diffCommits_info_243_ldest;
    rand bit [7:0]   io_diffCommits_info_243_pdest;
    rand bit         io_diffCommits_info_243_rfWen;
    rand bit         io_diffCommits_info_243_fpWen;
    rand bit         io_diffCommits_info_243_vecWen;
    rand bit         io_diffCommits_info_243_v0Wen;
    rand bit         io_diffCommits_info_243_vlWen;
    rand bit [5:0]   io_diffCommits_info_244_ldest;
    rand bit [7:0]   io_diffCommits_info_244_pdest;
    rand bit         io_diffCommits_info_244_rfWen;
    rand bit         io_diffCommits_info_244_fpWen;
    rand bit         io_diffCommits_info_244_vecWen;
    rand bit         io_diffCommits_info_244_v0Wen;
    rand bit         io_diffCommits_info_244_vlWen;
    rand bit [5:0]   io_diffCommits_info_245_ldest;
    rand bit [7:0]   io_diffCommits_info_245_pdest;
    rand bit         io_diffCommits_info_245_rfWen;
    rand bit         io_diffCommits_info_245_fpWen;
    rand bit         io_diffCommits_info_245_vecWen;
    rand bit         io_diffCommits_info_245_v0Wen;
    rand bit         io_diffCommits_info_245_vlWen;
    rand bit [5:0]   io_diffCommits_info_246_ldest;
    rand bit [7:0]   io_diffCommits_info_246_pdest;
    rand bit         io_diffCommits_info_246_rfWen;
    rand bit         io_diffCommits_info_246_fpWen;
    rand bit         io_diffCommits_info_246_vecWen;
    rand bit         io_diffCommits_info_246_v0Wen;
    rand bit         io_diffCommits_info_246_vlWen;
    rand bit [5:0]   io_diffCommits_info_247_ldest;
    rand bit [7:0]   io_diffCommits_info_247_pdest;
    rand bit         io_diffCommits_info_247_rfWen;
    rand bit         io_diffCommits_info_247_fpWen;
    rand bit         io_diffCommits_info_247_vecWen;
    rand bit         io_diffCommits_info_247_v0Wen;
    rand bit         io_diffCommits_info_247_vlWen;
    rand bit [5:0]   io_diffCommits_info_248_ldest;
    rand bit [7:0]   io_diffCommits_info_248_pdest;
    rand bit         io_diffCommits_info_248_rfWen;
    rand bit         io_diffCommits_info_248_fpWen;
    rand bit         io_diffCommits_info_248_vecWen;
    rand bit         io_diffCommits_info_248_v0Wen;
    rand bit         io_diffCommits_info_248_vlWen;
    rand bit [5:0]   io_diffCommits_info_249_ldest;
    rand bit [7:0]   io_diffCommits_info_249_pdest;
    rand bit         io_diffCommits_info_249_rfWen;
    rand bit         io_diffCommits_info_249_fpWen;
    rand bit         io_diffCommits_info_249_vecWen;
    rand bit         io_diffCommits_info_249_v0Wen;
    rand bit         io_diffCommits_info_249_vlWen;
    rand bit [5:0]   io_diffCommits_info_250_ldest;
    rand bit [7:0]   io_diffCommits_info_250_pdest;
    rand bit         io_diffCommits_info_250_rfWen;
    rand bit         io_diffCommits_info_250_fpWen;
    rand bit         io_diffCommits_info_250_vecWen;
    rand bit         io_diffCommits_info_250_v0Wen;
    rand bit         io_diffCommits_info_250_vlWen;
    rand bit [5:0]   io_diffCommits_info_251_ldest;
    rand bit [7:0]   io_diffCommits_info_251_pdest;
    rand bit         io_diffCommits_info_251_rfWen;
    rand bit         io_diffCommits_info_251_fpWen;
    rand bit         io_diffCommits_info_251_vecWen;
    rand bit         io_diffCommits_info_251_v0Wen;
    rand bit         io_diffCommits_info_251_vlWen;
    rand bit [5:0]   io_diffCommits_info_252_ldest;
    rand bit [7:0]   io_diffCommits_info_252_pdest;
    rand bit         io_diffCommits_info_252_rfWen;
    rand bit         io_diffCommits_info_252_fpWen;
    rand bit         io_diffCommits_info_252_vecWen;
    rand bit         io_diffCommits_info_252_v0Wen;
    rand bit         io_diffCommits_info_252_vlWen;
    rand bit [5:0]   io_diffCommits_info_253_ldest;
    rand bit [7:0]   io_diffCommits_info_253_pdest;
    rand bit         io_diffCommits_info_253_rfWen;
    rand bit         io_diffCommits_info_253_fpWen;
    rand bit         io_diffCommits_info_253_vecWen;
    rand bit         io_diffCommits_info_253_v0Wen;
    rand bit         io_diffCommits_info_253_vlWen;
    rand bit [5:0]   io_diffCommits_info_254_ldest;
    rand bit [7:0]   io_diffCommits_info_254_pdest;
    rand bit         io_diffCommits_info_254_rfWen;
    rand bit         io_diffCommits_info_254_fpWen;
    rand bit         io_diffCommits_info_254_vecWen;
    rand bit         io_diffCommits_info_254_v0Wen;
    rand bit         io_diffCommits_info_254_vlWen;
    rand bit [5:0]   io_diffCommits_info_255_ldest;
    rand bit [7:0]   io_diffCommits_info_255_pdest;
    rand bit [5:0]   io_diffCommits_info_256_ldest;
    rand bit [7:0]   io_diffCommits_info_256_pdest;
    rand bit [5:0]   io_diffCommits_info_257_ldest;
    rand bit [7:0]   io_diffCommits_info_257_pdest;
    rand bit [5:0]   io_diffCommits_info_258_ldest;
    rand bit [7:0]   io_diffCommits_info_258_pdest;
    rand bit [5:0]   io_diffCommits_info_259_ldest;
    rand bit [7:0]   io_diffCommits_info_259_pdest;
    rand bit [5:0]   io_diffCommits_info_260_ldest;
    rand bit [7:0]   io_diffCommits_info_260_pdest;
    rand bit [5:0]   io_diffCommits_info_261_ldest;
    rand bit [7:0]   io_diffCommits_info_261_pdest;
    rand bit [5:0]   io_diffCommits_info_262_ldest;
    rand bit [7:0]   io_diffCommits_info_262_pdest;
    rand bit [5:0]   io_diffCommits_info_263_ldest;
    rand bit [7:0]   io_diffCommits_info_263_pdest;
    rand bit [5:0]   io_diffCommits_info_264_ldest;
    rand bit [7:0]   io_diffCommits_info_264_pdest;
    rand bit [5:0]   io_diffCommits_info_265_ldest;
    rand bit [7:0]   io_diffCommits_info_265_pdest;
    rand bit [5:0]   io_diffCommits_info_266_ldest;
    rand bit [7:0]   io_diffCommits_info_266_pdest;
    rand bit [5:0]   io_diffCommits_info_267_ldest;
    rand bit [7:0]   io_diffCommits_info_267_pdest;
    rand bit [5:0]   io_diffCommits_info_268_ldest;
    rand bit [7:0]   io_diffCommits_info_268_pdest;
    rand bit [5:0]   io_diffCommits_info_269_ldest;
    rand bit [7:0]   io_diffCommits_info_269_pdest;
    rand bit [5:0]   io_diffCommits_info_270_ldest;
    rand bit [7:0]   io_diffCommits_info_270_pdest;
    rand bit [5:0]   io_diffCommits_info_271_ldest;
    rand bit [7:0]   io_diffCommits_info_271_pdest;
    rand bit [5:0]   io_diffCommits_info_272_ldest;
    rand bit [7:0]   io_diffCommits_info_272_pdest;
    rand bit [5:0]   io_diffCommits_info_273_ldest;
    rand bit [7:0]   io_diffCommits_info_273_pdest;
    rand bit [5:0]   io_diffCommits_info_274_ldest;
    rand bit [7:0]   io_diffCommits_info_274_pdest;
    rand bit [5:0]   io_diffCommits_info_275_ldest;
    rand bit [7:0]   io_diffCommits_info_275_pdest;
    rand bit [5:0]   io_diffCommits_info_276_ldest;
    rand bit [7:0]   io_diffCommits_info_276_pdest;
    rand bit [5:0]   io_diffCommits_info_277_ldest;
    rand bit [7:0]   io_diffCommits_info_277_pdest;
    rand bit [5:0]   io_diffCommits_info_278_ldest;
    rand bit [7:0]   io_diffCommits_info_278_pdest;
    rand bit [5:0]   io_diffCommits_info_279_ldest;
    rand bit [7:0]   io_diffCommits_info_279_pdest;
    rand bit [5:0]   io_diffCommits_info_280_ldest;
    rand bit [7:0]   io_diffCommits_info_280_pdest;
    rand bit [5:0]   io_diffCommits_info_281_ldest;
    rand bit [7:0]   io_diffCommits_info_281_pdest;
    rand bit [5:0]   io_diffCommits_info_282_ldest;
    rand bit [7:0]   io_diffCommits_info_282_pdest;
    rand bit [5:0]   io_diffCommits_info_283_ldest;
    rand bit [7:0]   io_diffCommits_info_283_pdest;
    rand bit [5:0]   io_diffCommits_info_284_ldest;
    rand bit [7:0]   io_diffCommits_info_284_pdest;
    rand bit [5:0]   io_diffCommits_info_285_ldest;
    rand bit [7:0]   io_diffCommits_info_285_pdest;
    rand bit [5:0]   io_diffCommits_info_286_ldest;
    rand bit [7:0]   io_diffCommits_info_286_pdest;
    rand bit [5:0]   io_diffCommits_info_287_ldest;
    rand bit [7:0]   io_diffCommits_info_287_pdest;
    rand bit [5:0]   io_diffCommits_info_288_ldest;
    rand bit [7:0]   io_diffCommits_info_288_pdest;
    rand bit [5:0]   io_diffCommits_info_289_ldest;
    rand bit [7:0]   io_diffCommits_info_289_pdest;
    rand bit [5:0]   io_diffCommits_info_290_ldest;
    rand bit [7:0]   io_diffCommits_info_290_pdest;
    rand bit [5:0]   io_diffCommits_info_291_ldest;
    rand bit [7:0]   io_diffCommits_info_291_pdest;
    rand bit [5:0]   io_diffCommits_info_292_ldest;
    rand bit [7:0]   io_diffCommits_info_292_pdest;
    rand bit [5:0]   io_diffCommits_info_293_ldest;
    rand bit [7:0]   io_diffCommits_info_293_pdest;
    rand bit [5:0]   io_diffCommits_info_294_ldest;
    rand bit [7:0]   io_diffCommits_info_294_pdest;
    rand bit [5:0]   io_diffCommits_info_295_ldest;
    rand bit [7:0]   io_diffCommits_info_295_pdest;
    rand bit [5:0]   io_diffCommits_info_296_ldest;
    rand bit [7:0]   io_diffCommits_info_296_pdest;
    rand bit [5:0]   io_diffCommits_info_297_ldest;
    rand bit [7:0]   io_diffCommits_info_297_pdest;
    rand bit [5:0]   io_diffCommits_info_298_ldest;
    rand bit [7:0]   io_diffCommits_info_298_pdest;
    rand bit [5:0]   io_diffCommits_info_299_ldest;
    rand bit [7:0]   io_diffCommits_info_299_pdest;
    rand bit [5:0]   io_diffCommits_info_300_ldest;
    rand bit [7:0]   io_diffCommits_info_300_pdest;
    rand bit [5:0]   io_diffCommits_info_301_ldest;
    rand bit [7:0]   io_diffCommits_info_301_pdest;
    rand bit [5:0]   io_diffCommits_info_302_ldest;
    rand bit [7:0]   io_diffCommits_info_302_pdest;
    rand bit [5:0]   io_diffCommits_info_303_ldest;
    rand bit [7:0]   io_diffCommits_info_303_pdest;
    rand bit [5:0]   io_diffCommits_info_304_ldest;
    rand bit [7:0]   io_diffCommits_info_304_pdest;
    rand bit [5:0]   io_diffCommits_info_305_ldest;
    rand bit [7:0]   io_diffCommits_info_305_pdest;
    rand bit [5:0]   io_diffCommits_info_306_ldest;
    rand bit [7:0]   io_diffCommits_info_306_pdest;
    rand bit [5:0]   io_diffCommits_info_307_ldest;
    rand bit [7:0]   io_diffCommits_info_307_pdest;
    rand bit [5:0]   io_diffCommits_info_308_ldest;
    rand bit [7:0]   io_diffCommits_info_308_pdest;
    rand bit [5:0]   io_diffCommits_info_309_ldest;
    rand bit [7:0]   io_diffCommits_info_309_pdest;
    rand bit [5:0]   io_diffCommits_info_310_ldest;
    rand bit [7:0]   io_diffCommits_info_310_pdest;
    rand bit [5:0]   io_diffCommits_info_311_ldest;
    rand bit [7:0]   io_diffCommits_info_311_pdest;
    rand bit [5:0]   io_diffCommits_info_312_ldest;
    rand bit [7:0]   io_diffCommits_info_312_pdest;
    rand bit [5:0]   io_diffCommits_info_313_ldest;
    rand bit [7:0]   io_diffCommits_info_313_pdest;
    rand bit [5:0]   io_diffCommits_info_314_ldest;
    rand bit [7:0]   io_diffCommits_info_314_pdest;
    rand bit [5:0]   io_diffCommits_info_315_ldest;
    rand bit [7:0]   io_diffCommits_info_315_pdest;
    rand bit [5:0]   io_diffCommits_info_316_ldest;
    rand bit [7:0]   io_diffCommits_info_316_pdest;
    rand bit [5:0]   io_diffCommits_info_317_ldest;
    rand bit [7:0]   io_diffCommits_info_317_pdest;
    rand bit [5:0]   io_diffCommits_info_318_ldest;
    rand bit [7:0]   io_diffCommits_info_318_pdest;
    rand bit [5:0]   io_diffCommits_info_319_ldest;
    rand bit [7:0]   io_diffCommits_info_319_pdest;
    rand bit [5:0]   io_diffCommits_info_320_ldest;
    rand bit [7:0]   io_diffCommits_info_320_pdest;
    rand bit [5:0]   io_diffCommits_info_321_ldest;
    rand bit [7:0]   io_diffCommits_info_321_pdest;
    rand bit [5:0]   io_diffCommits_info_322_ldest;
    rand bit [7:0]   io_diffCommits_info_322_pdest;
    rand bit [5:0]   io_diffCommits_info_323_ldest;
    rand bit [7:0]   io_diffCommits_info_323_pdest;
    rand bit [5:0]   io_diffCommits_info_324_ldest;
    rand bit [7:0]   io_diffCommits_info_324_pdest;
    rand bit [5:0]   io_diffCommits_info_325_ldest;
    rand bit [7:0]   io_diffCommits_info_325_pdest;
    rand bit [5:0]   io_diffCommits_info_326_ldest;
    rand bit [7:0]   io_diffCommits_info_326_pdest;
    rand bit [5:0]   io_diffCommits_info_327_ldest;
    rand bit [7:0]   io_diffCommits_info_327_pdest;
    rand bit [5:0]   io_diffCommits_info_328_ldest;
    rand bit [7:0]   io_diffCommits_info_328_pdest;
    rand bit [5:0]   io_diffCommits_info_329_ldest;
    rand bit [7:0]   io_diffCommits_info_329_pdest;
    rand bit [5:0]   io_diffCommits_info_330_ldest;
    rand bit [7:0]   io_diffCommits_info_330_pdest;
    rand bit [5:0]   io_diffCommits_info_331_ldest;
    rand bit [7:0]   io_diffCommits_info_331_pdest;
    rand bit [5:0]   io_diffCommits_info_332_ldest;
    rand bit [7:0]   io_diffCommits_info_332_pdest;
    rand bit [5:0]   io_diffCommits_info_333_ldest;
    rand bit [7:0]   io_diffCommits_info_333_pdest;
    rand bit [5:0]   io_diffCommits_info_334_ldest;
    rand bit [7:0]   io_diffCommits_info_334_pdest;
    rand bit [5:0]   io_diffCommits_info_335_ldest;
    rand bit [7:0]   io_diffCommits_info_335_pdest;
    rand bit [5:0]   io_diffCommits_info_336_ldest;
    rand bit [7:0]   io_diffCommits_info_336_pdest;
    rand bit [5:0]   io_diffCommits_info_337_ldest;
    rand bit [7:0]   io_diffCommits_info_337_pdest;
    rand bit [5:0]   io_diffCommits_info_338_ldest;
    rand bit [7:0]   io_diffCommits_info_338_pdest;
    rand bit [5:0]   io_diffCommits_info_339_ldest;
    rand bit [7:0]   io_diffCommits_info_339_pdest;
    rand bit [5:0]   io_diffCommits_info_340_ldest;
    rand bit [7:0]   io_diffCommits_info_340_pdest;
    rand bit [5:0]   io_diffCommits_info_341_ldest;
    rand bit [7:0]   io_diffCommits_info_341_pdest;
    rand bit [5:0]   io_diffCommits_info_342_ldest;
    rand bit [7:0]   io_diffCommits_info_342_pdest;
    rand bit [5:0]   io_diffCommits_info_343_ldest;
    rand bit [7:0]   io_diffCommits_info_343_pdest;
    rand bit [5:0]   io_diffCommits_info_344_ldest;
    rand bit [7:0]   io_diffCommits_info_344_pdest;
    rand bit [5:0]   io_diffCommits_info_345_ldest;
    rand bit [7:0]   io_diffCommits_info_345_pdest;
    rand bit [5:0]   io_diffCommits_info_346_ldest;
    rand bit [7:0]   io_diffCommits_info_346_pdest;
    rand bit [5:0]   io_diffCommits_info_347_ldest;
    rand bit [7:0]   io_diffCommits_info_347_pdest;
    rand bit [5:0]   io_diffCommits_info_348_ldest;
    rand bit [7:0]   io_diffCommits_info_348_pdest;
    rand bit [5:0]   io_diffCommits_info_349_ldest;
    rand bit [7:0]   io_diffCommits_info_349_pdest;
    rand bit [5:0]   io_diffCommits_info_350_ldest;
    rand bit [7:0]   io_diffCommits_info_350_pdest;
    rand bit [5:0]   io_diffCommits_info_351_ldest;
    rand bit [7:0]   io_diffCommits_info_351_pdest;
    rand bit [5:0]   io_diffCommits_info_352_ldest;
    rand bit [7:0]   io_diffCommits_info_352_pdest;
    rand bit [5:0]   io_diffCommits_info_353_ldest;
    rand bit [7:0]   io_diffCommits_info_353_pdest;
    rand bit [5:0]   io_diffCommits_info_354_ldest;
    rand bit [7:0]   io_diffCommits_info_354_pdest;
    rand bit [5:0]   io_diffCommits_info_355_ldest;
    rand bit [7:0]   io_diffCommits_info_355_pdest;
    rand bit [5:0]   io_diffCommits_info_356_ldest;
    rand bit [7:0]   io_diffCommits_info_356_pdest;
    rand bit [5:0]   io_diffCommits_info_357_ldest;
    rand bit [7:0]   io_diffCommits_info_357_pdest;
    rand bit [5:0]   io_diffCommits_info_358_ldest;
    rand bit [7:0]   io_diffCommits_info_358_pdest;
    rand bit [5:0]   io_diffCommits_info_359_ldest;
    rand bit [7:0]   io_diffCommits_info_359_pdest;
    rand bit [5:0]   io_diffCommits_info_360_ldest;
    rand bit [7:0]   io_diffCommits_info_360_pdest;
    rand bit [5:0]   io_diffCommits_info_361_ldest;
    rand bit [7:0]   io_diffCommits_info_361_pdest;
    rand bit [5:0]   io_diffCommits_info_362_ldest;
    rand bit [7:0]   io_diffCommits_info_362_pdest;
    rand bit [5:0]   io_diffCommits_info_363_ldest;
    rand bit [7:0]   io_diffCommits_info_363_pdest;
    rand bit [5:0]   io_diffCommits_info_364_ldest;
    rand bit [7:0]   io_diffCommits_info_364_pdest;
    rand bit [5:0]   io_diffCommits_info_365_ldest;
    rand bit [7:0]   io_diffCommits_info_365_pdest;
    rand bit [5:0]   io_diffCommits_info_366_ldest;
    rand bit [7:0]   io_diffCommits_info_366_pdest;
    rand bit [5:0]   io_diffCommits_info_367_ldest;
    rand bit [7:0]   io_diffCommits_info_367_pdest;
    rand bit [5:0]   io_diffCommits_info_368_ldest;
    rand bit [7:0]   io_diffCommits_info_368_pdest;
    rand bit [5:0]   io_diffCommits_info_369_ldest;
    rand bit [7:0]   io_diffCommits_info_369_pdest;
    rand bit [5:0]   io_diffCommits_info_370_ldest;
    rand bit [7:0]   io_diffCommits_info_370_pdest;
    rand bit [5:0]   io_diffCommits_info_371_ldest;
    rand bit [7:0]   io_diffCommits_info_371_pdest;
    rand bit [5:0]   io_diffCommits_info_372_ldest;
    rand bit [7:0]   io_diffCommits_info_372_pdest;
    rand bit [5:0]   io_diffCommits_info_373_ldest;
    rand bit [7:0]   io_diffCommits_info_373_pdest;
    rand bit [5:0]   io_diffCommits_info_374_ldest;
    rand bit [7:0]   io_diffCommits_info_374_pdest;
    rand bit [5:0]   io_diffCommits_info_375_ldest;
    rand bit [7:0]   io_diffCommits_info_375_pdest;
    rand bit [5:0]   io_diffCommits_info_376_ldest;
    rand bit [7:0]   io_diffCommits_info_376_pdest;
    rand bit [5:0]   io_diffCommits_info_377_ldest;
    rand bit [7:0]   io_diffCommits_info_377_pdest;
    rand bit [5:0]   io_diffCommits_info_378_ldest;
    rand bit [7:0]   io_diffCommits_info_378_pdest;
    rand bit [5:0]   io_diffCommits_info_379_ldest;
    rand bit [7:0]   io_diffCommits_info_379_pdest;
    rand bit [5:0]   io_diffCommits_info_380_ldest;
    rand bit [7:0]   io_diffCommits_info_380_pdest;
    rand bit [5:0]   io_diffCommits_info_381_ldest;
    rand bit [7:0]   io_diffCommits_info_381_pdest;
    rand bit [5:0]   io_diffCommits_info_382_ldest;
    rand bit [7:0]   io_diffCommits_info_382_pdest;
    rand bit [5:0]   io_diffCommits_info_383_ldest;
    rand bit [7:0]   io_diffCommits_info_383_pdest;
    rand bit [5:0]   io_diffCommits_info_384_ldest;
    rand bit [7:0]   io_diffCommits_info_384_pdest;
    rand bit [5:0]   io_diffCommits_info_385_ldest;
    rand bit [7:0]   io_diffCommits_info_385_pdest;
    rand bit [5:0]   io_diffCommits_info_386_ldest;
    rand bit [7:0]   io_diffCommits_info_386_pdest;
    rand bit [5:0]   io_diffCommits_info_387_ldest;
    rand bit [7:0]   io_diffCommits_info_387_pdest;
    rand bit [5:0]   io_diffCommits_info_388_ldest;
    rand bit [7:0]   io_diffCommits_info_388_pdest;
    rand bit [5:0]   io_diffCommits_info_389_ldest;
    rand bit [7:0]   io_diffCommits_info_389_pdest;
    rand bit [3:0]   io_lsq_scommit    ;
    rand bit         io_lsq_pendingMMIOld;
    rand bit         io_lsq_pendingst  ;
    rand bit         io_lsq_pendingPtr_flag;
    rand bit [7:0]   io_lsq_pendingPtr_value;
    rand bit         io_robDeqPtr_flag ;
    rand bit [7:0]   io_robDeqPtr_value;
    rand bit         io_csr_fflags_valid;
    rand bit [4:0]   io_csr_fflags_bits;
    rand bit         io_csr_vxsat_valid;
    rand bit         io_csr_vxsat_bits ;
    rand bit         io_csr_vstart_valid;
    rand bit [63:0]  io_csr_vstart_bits;
    rand bit         io_csr_dirty_fs   ;
    rand bit         io_csr_dirty_vs   ;
    rand bit [6:0]   io_csr_perfinfo_retiredInstr;
    rand bit         io_cpu_halt       ;
    rand bit         io_wfi_wfiReq     ;
    rand bit         io_toDecode_isResumeVType;
    rand bit         io_toDecode_walkToArchVType;
    rand bit         io_toDecode_walkVType_valid;
    rand bit         io_toDecode_walkVType_bits_illegal;
    rand bit         io_toDecode_walkVType_bits_vma;
    rand bit         io_toDecode_walkVType_bits_vta;
    rand bit [1:0]   io_toDecode_walkVType_bits_vsew;
    rand bit [2:0]   io_toDecode_walkVType_bits_vlmul;
    rand bit         io_toDecode_commitVType_vtype_valid;
    rand bit         io_toDecode_commitVType_vtype_bits_illegal;
    rand bit         io_toDecode_commitVType_vtype_bits_vma;
    rand bit         io_toDecode_commitVType_vtype_bits_vta;
    rand bit [1:0]   io_toDecode_commitVType_vtype_bits_vsew;
    rand bit [2:0]   io_toDecode_commitVType_vtype_bits_vlmul;
    rand bit         io_toDecode_commitVType_hasVsetvl;
    rand bit         io_readGPAMemAddr_valid;
    rand bit [5:0]   io_readGPAMemAddr_bits_ftqPtr_value;
    rand bit [3:0]   io_readGPAMemAddr_bits_ftqOffset;
    rand bit         io_toVecExcpMod_logicPhyRegMap_0_valid;
    rand bit [5:0]   io_toVecExcpMod_logicPhyRegMap_0_bits_lreg;
    rand bit [6:0]   io_toVecExcpMod_logicPhyRegMap_0_bits_preg;
    rand bit         io_toVecExcpMod_logicPhyRegMap_1_valid;
    rand bit [5:0]   io_toVecExcpMod_logicPhyRegMap_1_bits_lreg;
    rand bit [6:0]   io_toVecExcpMod_logicPhyRegMap_1_bits_preg;
    rand bit         io_toVecExcpMod_logicPhyRegMap_2_valid;
    rand bit [5:0]   io_toVecExcpMod_logicPhyRegMap_2_bits_lreg;
    rand bit [6:0]   io_toVecExcpMod_logicPhyRegMap_2_bits_preg;
    rand bit         io_toVecExcpMod_logicPhyRegMap_3_valid;
    rand bit [5:0]   io_toVecExcpMod_logicPhyRegMap_3_bits_lreg;
    rand bit [6:0]   io_toVecExcpMod_logicPhyRegMap_3_bits_preg;
    rand bit         io_toVecExcpMod_logicPhyRegMap_4_valid;
    rand bit [5:0]   io_toVecExcpMod_logicPhyRegMap_4_bits_lreg;
    rand bit [6:0]   io_toVecExcpMod_logicPhyRegMap_4_bits_preg;
    rand bit         io_toVecExcpMod_logicPhyRegMap_5_valid;
    rand bit [5:0]   io_toVecExcpMod_logicPhyRegMap_5_bits_lreg;
    rand bit [6:0]   io_toVecExcpMod_logicPhyRegMap_5_bits_preg;
    rand bit         io_toVecExcpMod_excpInfo_valid;
    rand bit [6:0]   io_toVecExcpMod_excpInfo_bits_vstart;
    rand bit [1:0]   io_toVecExcpMod_excpInfo_bits_vsew;
    rand bit [1:0]   io_toVecExcpMod_excpInfo_bits_veew;
    rand bit [2:0]   io_toVecExcpMod_excpInfo_bits_vlmul;
    rand bit [2:0]   io_toVecExcpMod_excpInfo_bits_nf;
    rand bit         io_toVecExcpMod_excpInfo_bits_isStride;
    rand bit         io_toVecExcpMod_excpInfo_bits_isIndexed;
    rand bit         io_toVecExcpMod_excpInfo_bits_isWhole;
    rand bit         io_toVecExcpMod_excpInfo_bits_isVlm;
    rand bit [49:0]  io_storeDebugInfo_1_pc;
    rand bit [5:0]   io_perf_0_value   ;
    rand bit [5:0]   io_perf_1_value   ;
    rand bit [5:0]   io_perf_2_value   ;
    rand bit [5:0]   io_perf_3_value   ;
    rand bit [5:0]   io_perf_4_value   ;
    rand bit [5:0]   io_perf_5_value   ;
    rand bit [5:0]   io_perf_6_value   ;
    rand bit [5:0]   io_perf_7_value   ;
    rand bit [5:0]   io_perf_8_value   ;
    rand bit [5:0]   io_perf_9_value   ;
    rand bit [5:0]   io_perf_10_value  ;
    rand bit [5:0]   io_perf_11_value  ;
    rand bit [5:0]   io_perf_12_value  ;
    rand bit [5:0]   io_perf_13_value  ;
    rand bit [5:0]   io_perf_14_value  ;
    rand bit [5:0]   io_perf_15_value  ;
    rand bit [5:0]   io_perf_16_value  ;
    rand bit [5:0]   io_perf_17_value  ;
    rand bit         io_error_0        ;

    extern constraint default_io_enq_canAccept_cons;
    extern constraint default_io_enq_canAcceptForDispatch_cons;
    extern constraint default_io_enq_isEmpty_cons;
    extern constraint default_io_flushOut_valid_cons;
    extern constraint default_io_flushOut_bits_isRVC_cons;
    extern constraint default_io_flushOut_bits_robIdx_flag_cons;
    extern constraint default_io_flushOut_bits_robIdx_value_cons;
    extern constraint default_io_flushOut_bits_ftqIdx_flag_cons;
    extern constraint default_io_flushOut_bits_ftqIdx_value_cons;
    extern constraint default_io_flushOut_bits_ftqOffset_cons;
    extern constraint default_io_flushOut_bits_level_cons;
    extern constraint default_io_exception_valid_cons;
    extern constraint default_io_exception_bits_instr_cons;
    extern constraint default_io_exception_bits_commitType_cons;
    extern constraint default_io_exception_bits_exceptionVec_0_cons;
    extern constraint default_io_exception_bits_exceptionVec_1_cons;
    extern constraint default_io_exception_bits_exceptionVec_2_cons;
    extern constraint default_io_exception_bits_exceptionVec_3_cons;
    extern constraint default_io_exception_bits_exceptionVec_4_cons;
    extern constraint default_io_exception_bits_exceptionVec_5_cons;
    extern constraint default_io_exception_bits_exceptionVec_6_cons;
    extern constraint default_io_exception_bits_exceptionVec_7_cons;
    extern constraint default_io_exception_bits_exceptionVec_8_cons;
    extern constraint default_io_exception_bits_exceptionVec_9_cons;
    extern constraint default_io_exception_bits_exceptionVec_10_cons;
    extern constraint default_io_exception_bits_exceptionVec_11_cons;
    extern constraint default_io_exception_bits_exceptionVec_12_cons;
    extern constraint default_io_exception_bits_exceptionVec_13_cons;
    extern constraint default_io_exception_bits_exceptionVec_14_cons;
    extern constraint default_io_exception_bits_exceptionVec_15_cons;
    extern constraint default_io_exception_bits_exceptionVec_16_cons;
    extern constraint default_io_exception_bits_exceptionVec_17_cons;
    extern constraint default_io_exception_bits_exceptionVec_18_cons;
    extern constraint default_io_exception_bits_exceptionVec_19_cons;
    extern constraint default_io_exception_bits_exceptionVec_20_cons;
    extern constraint default_io_exception_bits_exceptionVec_21_cons;
    extern constraint default_io_exception_bits_exceptionVec_22_cons;
    extern constraint default_io_exception_bits_exceptionVec_23_cons;
    extern constraint default_io_exception_bits_isPcBkpt_cons;
    extern constraint default_io_exception_bits_isFetchMalAddr_cons;
    extern constraint default_io_exception_bits_gpaddr_cons;
    extern constraint default_io_exception_bits_singleStep_cons;
    extern constraint default_io_exception_bits_crossPageIPFFix_cons;
    extern constraint default_io_exception_bits_isInterrupt_cons;
    extern constraint default_io_exception_bits_isHls_cons;
    extern constraint default_io_exception_bits_trigger_cons;
    extern constraint default_io_exception_bits_isForVSnonLeafPTE_cons;
    extern constraint default_io_commits_isCommit_cons;
    extern constraint default_io_commits_commitValid_0_cons;
    extern constraint default_io_commits_commitValid_1_cons;
    extern constraint default_io_commits_commitValid_2_cons;
    extern constraint default_io_commits_commitValid_3_cons;
    extern constraint default_io_commits_commitValid_4_cons;
    extern constraint default_io_commits_commitValid_5_cons;
    extern constraint default_io_commits_commitValid_6_cons;
    extern constraint default_io_commits_commitValid_7_cons;
    extern constraint default_io_commits_isWalk_cons;
    extern constraint default_io_commits_walkValid_0_cons;
    extern constraint default_io_commits_walkValid_1_cons;
    extern constraint default_io_commits_walkValid_2_cons;
    extern constraint default_io_commits_walkValid_3_cons;
    extern constraint default_io_commits_walkValid_4_cons;
    extern constraint default_io_commits_walkValid_5_cons;
    extern constraint default_io_commits_walkValid_6_cons;
    extern constraint default_io_commits_walkValid_7_cons;
    extern constraint default_io_commits_info_0_walk_v_cons;
    extern constraint default_io_commits_info_0_commit_v_cons;
    extern constraint default_io_commits_info_0_commit_w_cons;
    extern constraint default_io_commits_info_0_realDestSize_cons;
    extern constraint default_io_commits_info_0_interrupt_safe_cons;
    extern constraint default_io_commits_info_0_wflags_cons;
    extern constraint default_io_commits_info_0_fflags_cons;
    extern constraint default_io_commits_info_0_vxsat_cons;
    extern constraint default_io_commits_info_0_isRVC_cons;
    extern constraint default_io_commits_info_0_isVset_cons;
    extern constraint default_io_commits_info_0_isHls_cons;
    extern constraint default_io_commits_info_0_isVls_cons;
    extern constraint default_io_commits_info_0_vls_cons;
    extern constraint default_io_commits_info_0_mmio_cons;
    extern constraint default_io_commits_info_0_commitType_cons;
    extern constraint default_io_commits_info_0_ftqIdx_flag_cons;
    extern constraint default_io_commits_info_0_ftqIdx_value_cons;
    extern constraint default_io_commits_info_0_ftqOffset_cons;
    extern constraint default_io_commits_info_0_instrSize_cons;
    extern constraint default_io_commits_info_0_fpWen_cons;
    extern constraint default_io_commits_info_0_rfWen_cons;
    extern constraint default_io_commits_info_0_needFlush_cons;
    extern constraint default_io_commits_info_0_traceBlockInPipe_itype_cons;
    extern constraint default_io_commits_info_0_traceBlockInPipe_iretire_cons;
    extern constraint default_io_commits_info_0_traceBlockInPipe_ilastsize_cons;
    extern constraint default_io_commits_info_0_debug_pc_cons;
    extern constraint default_io_commits_info_0_debug_instr_cons;
    extern constraint default_io_commits_info_0_debug_ldest_cons;
    extern constraint default_io_commits_info_0_debug_pdest_cons;
    extern constraint default_io_commits_info_0_debug_otherPdest_0_cons;
    extern constraint default_io_commits_info_0_debug_otherPdest_1_cons;
    extern constraint default_io_commits_info_0_debug_otherPdest_2_cons;
    extern constraint default_io_commits_info_0_debug_otherPdest_3_cons;
    extern constraint default_io_commits_info_0_debug_otherPdest_4_cons;
    extern constraint default_io_commits_info_0_debug_otherPdest_5_cons;
    extern constraint default_io_commits_info_0_debug_otherPdest_6_cons;
    extern constraint default_io_commits_info_0_debug_fuType_cons;
    extern constraint default_io_commits_info_0_dirtyFs_cons;
    extern constraint default_io_commits_info_0_dirtyVs_cons;
    extern constraint default_io_commits_info_1_walk_v_cons;
    extern constraint default_io_commits_info_1_commit_v_cons;
    extern constraint default_io_commits_info_1_commit_w_cons;
    extern constraint default_io_commits_info_1_realDestSize_cons;
    extern constraint default_io_commits_info_1_interrupt_safe_cons;
    extern constraint default_io_commits_info_1_wflags_cons;
    extern constraint default_io_commits_info_1_fflags_cons;
    extern constraint default_io_commits_info_1_vxsat_cons;
    extern constraint default_io_commits_info_1_isRVC_cons;
    extern constraint default_io_commits_info_1_isVset_cons;
    extern constraint default_io_commits_info_1_isHls_cons;
    extern constraint default_io_commits_info_1_isVls_cons;
    extern constraint default_io_commits_info_1_vls_cons;
    extern constraint default_io_commits_info_1_mmio_cons;
    extern constraint default_io_commits_info_1_commitType_cons;
    extern constraint default_io_commits_info_1_ftqIdx_flag_cons;
    extern constraint default_io_commits_info_1_ftqIdx_value_cons;
    extern constraint default_io_commits_info_1_ftqOffset_cons;
    extern constraint default_io_commits_info_1_instrSize_cons;
    extern constraint default_io_commits_info_1_fpWen_cons;
    extern constraint default_io_commits_info_1_rfWen_cons;
    extern constraint default_io_commits_info_1_needFlush_cons;
    extern constraint default_io_commits_info_1_traceBlockInPipe_itype_cons;
    extern constraint default_io_commits_info_1_traceBlockInPipe_iretire_cons;
    extern constraint default_io_commits_info_1_traceBlockInPipe_ilastsize_cons;
    extern constraint default_io_commits_info_1_debug_pc_cons;
    extern constraint default_io_commits_info_1_debug_instr_cons;
    extern constraint default_io_commits_info_1_debug_ldest_cons;
    extern constraint default_io_commits_info_1_debug_pdest_cons;
    extern constraint default_io_commits_info_1_debug_otherPdest_0_cons;
    extern constraint default_io_commits_info_1_debug_otherPdest_1_cons;
    extern constraint default_io_commits_info_1_debug_otherPdest_2_cons;
    extern constraint default_io_commits_info_1_debug_otherPdest_3_cons;
    extern constraint default_io_commits_info_1_debug_otherPdest_4_cons;
    extern constraint default_io_commits_info_1_debug_otherPdest_5_cons;
    extern constraint default_io_commits_info_1_debug_otherPdest_6_cons;
    extern constraint default_io_commits_info_1_debug_fuType_cons;
    extern constraint default_io_commits_info_1_dirtyFs_cons;
    extern constraint default_io_commits_info_1_dirtyVs_cons;
    extern constraint default_io_commits_info_2_walk_v_cons;
    extern constraint default_io_commits_info_2_commit_v_cons;
    extern constraint default_io_commits_info_2_commit_w_cons;
    extern constraint default_io_commits_info_2_realDestSize_cons;
    extern constraint default_io_commits_info_2_interrupt_safe_cons;
    extern constraint default_io_commits_info_2_wflags_cons;
    extern constraint default_io_commits_info_2_fflags_cons;
    extern constraint default_io_commits_info_2_vxsat_cons;
    extern constraint default_io_commits_info_2_isRVC_cons;
    extern constraint default_io_commits_info_2_isVset_cons;
    extern constraint default_io_commits_info_2_isHls_cons;
    extern constraint default_io_commits_info_2_isVls_cons;
    extern constraint default_io_commits_info_2_vls_cons;
    extern constraint default_io_commits_info_2_mmio_cons;
    extern constraint default_io_commits_info_2_commitType_cons;
    extern constraint default_io_commits_info_2_ftqIdx_flag_cons;
    extern constraint default_io_commits_info_2_ftqIdx_value_cons;
    extern constraint default_io_commits_info_2_ftqOffset_cons;
    extern constraint default_io_commits_info_2_instrSize_cons;
    extern constraint default_io_commits_info_2_fpWen_cons;
    extern constraint default_io_commits_info_2_rfWen_cons;
    extern constraint default_io_commits_info_2_needFlush_cons;
    extern constraint default_io_commits_info_2_traceBlockInPipe_itype_cons;
    extern constraint default_io_commits_info_2_traceBlockInPipe_iretire_cons;
    extern constraint default_io_commits_info_2_traceBlockInPipe_ilastsize_cons;
    extern constraint default_io_commits_info_2_debug_pc_cons;
    extern constraint default_io_commits_info_2_debug_instr_cons;
    extern constraint default_io_commits_info_2_debug_ldest_cons;
    extern constraint default_io_commits_info_2_debug_pdest_cons;
    extern constraint default_io_commits_info_2_debug_otherPdest_0_cons;
    extern constraint default_io_commits_info_2_debug_otherPdest_1_cons;
    extern constraint default_io_commits_info_2_debug_otherPdest_2_cons;
    extern constraint default_io_commits_info_2_debug_otherPdest_3_cons;
    extern constraint default_io_commits_info_2_debug_otherPdest_4_cons;
    extern constraint default_io_commits_info_2_debug_otherPdest_5_cons;
    extern constraint default_io_commits_info_2_debug_otherPdest_6_cons;
    extern constraint default_io_commits_info_2_debug_fuType_cons;
    extern constraint default_io_commits_info_2_dirtyFs_cons;
    extern constraint default_io_commits_info_2_dirtyVs_cons;
    extern constraint default_io_commits_info_3_walk_v_cons;
    extern constraint default_io_commits_info_3_commit_v_cons;
    extern constraint default_io_commits_info_3_commit_w_cons;
    extern constraint default_io_commits_info_3_realDestSize_cons;
    extern constraint default_io_commits_info_3_interrupt_safe_cons;
    extern constraint default_io_commits_info_3_wflags_cons;
    extern constraint default_io_commits_info_3_fflags_cons;
    extern constraint default_io_commits_info_3_vxsat_cons;
    extern constraint default_io_commits_info_3_isRVC_cons;
    extern constraint default_io_commits_info_3_isVset_cons;
    extern constraint default_io_commits_info_3_isHls_cons;
    extern constraint default_io_commits_info_3_isVls_cons;
    extern constraint default_io_commits_info_3_vls_cons;
    extern constraint default_io_commits_info_3_mmio_cons;
    extern constraint default_io_commits_info_3_commitType_cons;
    extern constraint default_io_commits_info_3_ftqIdx_flag_cons;
    extern constraint default_io_commits_info_3_ftqIdx_value_cons;
    extern constraint default_io_commits_info_3_ftqOffset_cons;
    extern constraint default_io_commits_info_3_instrSize_cons;
    extern constraint default_io_commits_info_3_fpWen_cons;
    extern constraint default_io_commits_info_3_rfWen_cons;
    extern constraint default_io_commits_info_3_needFlush_cons;
    extern constraint default_io_commits_info_3_traceBlockInPipe_itype_cons;
    extern constraint default_io_commits_info_3_traceBlockInPipe_iretire_cons;
    extern constraint default_io_commits_info_3_traceBlockInPipe_ilastsize_cons;
    extern constraint default_io_commits_info_3_debug_pc_cons;
    extern constraint default_io_commits_info_3_debug_instr_cons;
    extern constraint default_io_commits_info_3_debug_ldest_cons;
    extern constraint default_io_commits_info_3_debug_pdest_cons;
    extern constraint default_io_commits_info_3_debug_otherPdest_0_cons;
    extern constraint default_io_commits_info_3_debug_otherPdest_1_cons;
    extern constraint default_io_commits_info_3_debug_otherPdest_2_cons;
    extern constraint default_io_commits_info_3_debug_otherPdest_3_cons;
    extern constraint default_io_commits_info_3_debug_otherPdest_4_cons;
    extern constraint default_io_commits_info_3_debug_otherPdest_5_cons;
    extern constraint default_io_commits_info_3_debug_otherPdest_6_cons;
    extern constraint default_io_commits_info_3_debug_fuType_cons;
    extern constraint default_io_commits_info_3_dirtyFs_cons;
    extern constraint default_io_commits_info_3_dirtyVs_cons;
    extern constraint default_io_commits_info_4_walk_v_cons;
    extern constraint default_io_commits_info_4_commit_v_cons;
    extern constraint default_io_commits_info_4_commit_w_cons;
    extern constraint default_io_commits_info_4_realDestSize_cons;
    extern constraint default_io_commits_info_4_interrupt_safe_cons;
    extern constraint default_io_commits_info_4_wflags_cons;
    extern constraint default_io_commits_info_4_fflags_cons;
    extern constraint default_io_commits_info_4_vxsat_cons;
    extern constraint default_io_commits_info_4_isRVC_cons;
    extern constraint default_io_commits_info_4_isVset_cons;
    extern constraint default_io_commits_info_4_isHls_cons;
    extern constraint default_io_commits_info_4_isVls_cons;
    extern constraint default_io_commits_info_4_vls_cons;
    extern constraint default_io_commits_info_4_mmio_cons;
    extern constraint default_io_commits_info_4_commitType_cons;
    extern constraint default_io_commits_info_4_ftqIdx_flag_cons;
    extern constraint default_io_commits_info_4_ftqIdx_value_cons;
    extern constraint default_io_commits_info_4_ftqOffset_cons;
    extern constraint default_io_commits_info_4_instrSize_cons;
    extern constraint default_io_commits_info_4_fpWen_cons;
    extern constraint default_io_commits_info_4_rfWen_cons;
    extern constraint default_io_commits_info_4_needFlush_cons;
    extern constraint default_io_commits_info_4_traceBlockInPipe_itype_cons;
    extern constraint default_io_commits_info_4_traceBlockInPipe_iretire_cons;
    extern constraint default_io_commits_info_4_traceBlockInPipe_ilastsize_cons;
    extern constraint default_io_commits_info_4_debug_pc_cons;
    extern constraint default_io_commits_info_4_debug_instr_cons;
    extern constraint default_io_commits_info_4_debug_ldest_cons;
    extern constraint default_io_commits_info_4_debug_pdest_cons;
    extern constraint default_io_commits_info_4_debug_otherPdest_0_cons;
    extern constraint default_io_commits_info_4_debug_otherPdest_1_cons;
    extern constraint default_io_commits_info_4_debug_otherPdest_2_cons;
    extern constraint default_io_commits_info_4_debug_otherPdest_3_cons;
    extern constraint default_io_commits_info_4_debug_otherPdest_4_cons;
    extern constraint default_io_commits_info_4_debug_otherPdest_5_cons;
    extern constraint default_io_commits_info_4_debug_otherPdest_6_cons;
    extern constraint default_io_commits_info_4_debug_fuType_cons;
    extern constraint default_io_commits_info_4_dirtyFs_cons;
    extern constraint default_io_commits_info_4_dirtyVs_cons;
    extern constraint default_io_commits_info_5_walk_v_cons;
    extern constraint default_io_commits_info_5_commit_v_cons;
    extern constraint default_io_commits_info_5_commit_w_cons;
    extern constraint default_io_commits_info_5_realDestSize_cons;
    extern constraint default_io_commits_info_5_interrupt_safe_cons;
    extern constraint default_io_commits_info_5_wflags_cons;
    extern constraint default_io_commits_info_5_fflags_cons;
    extern constraint default_io_commits_info_5_vxsat_cons;
    extern constraint default_io_commits_info_5_isRVC_cons;
    extern constraint default_io_commits_info_5_isVset_cons;
    extern constraint default_io_commits_info_5_isHls_cons;
    extern constraint default_io_commits_info_5_isVls_cons;
    extern constraint default_io_commits_info_5_vls_cons;
    extern constraint default_io_commits_info_5_mmio_cons;
    extern constraint default_io_commits_info_5_commitType_cons;
    extern constraint default_io_commits_info_5_ftqIdx_flag_cons;
    extern constraint default_io_commits_info_5_ftqIdx_value_cons;
    extern constraint default_io_commits_info_5_ftqOffset_cons;
    extern constraint default_io_commits_info_5_instrSize_cons;
    extern constraint default_io_commits_info_5_fpWen_cons;
    extern constraint default_io_commits_info_5_rfWen_cons;
    extern constraint default_io_commits_info_5_needFlush_cons;
    extern constraint default_io_commits_info_5_traceBlockInPipe_itype_cons;
    extern constraint default_io_commits_info_5_traceBlockInPipe_iretire_cons;
    extern constraint default_io_commits_info_5_traceBlockInPipe_ilastsize_cons;
    extern constraint default_io_commits_info_5_debug_pc_cons;
    extern constraint default_io_commits_info_5_debug_instr_cons;
    extern constraint default_io_commits_info_5_debug_ldest_cons;
    extern constraint default_io_commits_info_5_debug_pdest_cons;
    extern constraint default_io_commits_info_5_debug_otherPdest_0_cons;
    extern constraint default_io_commits_info_5_debug_otherPdest_1_cons;
    extern constraint default_io_commits_info_5_debug_otherPdest_2_cons;
    extern constraint default_io_commits_info_5_debug_otherPdest_3_cons;
    extern constraint default_io_commits_info_5_debug_otherPdest_4_cons;
    extern constraint default_io_commits_info_5_debug_otherPdest_5_cons;
    extern constraint default_io_commits_info_5_debug_otherPdest_6_cons;
    extern constraint default_io_commits_info_5_debug_fuType_cons;
    extern constraint default_io_commits_info_5_dirtyFs_cons;
    extern constraint default_io_commits_info_5_dirtyVs_cons;
    extern constraint default_io_commits_info_6_walk_v_cons;
    extern constraint default_io_commits_info_6_commit_v_cons;
    extern constraint default_io_commits_info_6_commit_w_cons;
    extern constraint default_io_commits_info_6_realDestSize_cons;
    extern constraint default_io_commits_info_6_interrupt_safe_cons;
    extern constraint default_io_commits_info_6_wflags_cons;
    extern constraint default_io_commits_info_6_fflags_cons;
    extern constraint default_io_commits_info_6_vxsat_cons;
    extern constraint default_io_commits_info_6_isRVC_cons;
    extern constraint default_io_commits_info_6_isVset_cons;
    extern constraint default_io_commits_info_6_isHls_cons;
    extern constraint default_io_commits_info_6_isVls_cons;
    extern constraint default_io_commits_info_6_vls_cons;
    extern constraint default_io_commits_info_6_mmio_cons;
    extern constraint default_io_commits_info_6_commitType_cons;
    extern constraint default_io_commits_info_6_ftqIdx_flag_cons;
    extern constraint default_io_commits_info_6_ftqIdx_value_cons;
    extern constraint default_io_commits_info_6_ftqOffset_cons;
    extern constraint default_io_commits_info_6_instrSize_cons;
    extern constraint default_io_commits_info_6_fpWen_cons;
    extern constraint default_io_commits_info_6_rfWen_cons;
    extern constraint default_io_commits_info_6_needFlush_cons;
    extern constraint default_io_commits_info_6_traceBlockInPipe_itype_cons;
    extern constraint default_io_commits_info_6_traceBlockInPipe_iretire_cons;
    extern constraint default_io_commits_info_6_traceBlockInPipe_ilastsize_cons;
    extern constraint default_io_commits_info_6_debug_pc_cons;
    extern constraint default_io_commits_info_6_debug_instr_cons;
    extern constraint default_io_commits_info_6_debug_ldest_cons;
    extern constraint default_io_commits_info_6_debug_pdest_cons;
    extern constraint default_io_commits_info_6_debug_otherPdest_0_cons;
    extern constraint default_io_commits_info_6_debug_otherPdest_1_cons;
    extern constraint default_io_commits_info_6_debug_otherPdest_2_cons;
    extern constraint default_io_commits_info_6_debug_otherPdest_3_cons;
    extern constraint default_io_commits_info_6_debug_otherPdest_4_cons;
    extern constraint default_io_commits_info_6_debug_otherPdest_5_cons;
    extern constraint default_io_commits_info_6_debug_otherPdest_6_cons;
    extern constraint default_io_commits_info_6_debug_fuType_cons;
    extern constraint default_io_commits_info_6_dirtyFs_cons;
    extern constraint default_io_commits_info_6_dirtyVs_cons;
    extern constraint default_io_commits_info_7_walk_v_cons;
    extern constraint default_io_commits_info_7_commit_v_cons;
    extern constraint default_io_commits_info_7_commit_w_cons;
    extern constraint default_io_commits_info_7_realDestSize_cons;
    extern constraint default_io_commits_info_7_interrupt_safe_cons;
    extern constraint default_io_commits_info_7_wflags_cons;
    extern constraint default_io_commits_info_7_fflags_cons;
    extern constraint default_io_commits_info_7_vxsat_cons;
    extern constraint default_io_commits_info_7_isRVC_cons;
    extern constraint default_io_commits_info_7_isVset_cons;
    extern constraint default_io_commits_info_7_isHls_cons;
    extern constraint default_io_commits_info_7_isVls_cons;
    extern constraint default_io_commits_info_7_vls_cons;
    extern constraint default_io_commits_info_7_mmio_cons;
    extern constraint default_io_commits_info_7_commitType_cons;
    extern constraint default_io_commits_info_7_ftqIdx_flag_cons;
    extern constraint default_io_commits_info_7_ftqIdx_value_cons;
    extern constraint default_io_commits_info_7_ftqOffset_cons;
    extern constraint default_io_commits_info_7_instrSize_cons;
    extern constraint default_io_commits_info_7_fpWen_cons;
    extern constraint default_io_commits_info_7_rfWen_cons;
    extern constraint default_io_commits_info_7_needFlush_cons;
    extern constraint default_io_commits_info_7_traceBlockInPipe_itype_cons;
    extern constraint default_io_commits_info_7_traceBlockInPipe_iretire_cons;
    extern constraint default_io_commits_info_7_traceBlockInPipe_ilastsize_cons;
    extern constraint default_io_commits_info_7_debug_pc_cons;
    extern constraint default_io_commits_info_7_debug_instr_cons;
    extern constraint default_io_commits_info_7_debug_ldest_cons;
    extern constraint default_io_commits_info_7_debug_pdest_cons;
    extern constraint default_io_commits_info_7_debug_otherPdest_0_cons;
    extern constraint default_io_commits_info_7_debug_otherPdest_1_cons;
    extern constraint default_io_commits_info_7_debug_otherPdest_2_cons;
    extern constraint default_io_commits_info_7_debug_otherPdest_3_cons;
    extern constraint default_io_commits_info_7_debug_otherPdest_4_cons;
    extern constraint default_io_commits_info_7_debug_otherPdest_5_cons;
    extern constraint default_io_commits_info_7_debug_otherPdest_6_cons;
    extern constraint default_io_commits_info_7_debug_fuType_cons;
    extern constraint default_io_commits_info_7_dirtyFs_cons;
    extern constraint default_io_commits_info_7_dirtyVs_cons;
    extern constraint default_io_commits_robIdx_0_flag_cons;
    extern constraint default_io_commits_robIdx_0_value_cons;
    extern constraint default_io_commits_robIdx_1_flag_cons;
    extern constraint default_io_commits_robIdx_1_value_cons;
    extern constraint default_io_commits_robIdx_2_flag_cons;
    extern constraint default_io_commits_robIdx_2_value_cons;
    extern constraint default_io_commits_robIdx_3_flag_cons;
    extern constraint default_io_commits_robIdx_3_value_cons;
    extern constraint default_io_commits_robIdx_4_flag_cons;
    extern constraint default_io_commits_robIdx_4_value_cons;
    extern constraint default_io_commits_robIdx_5_flag_cons;
    extern constraint default_io_commits_robIdx_5_value_cons;
    extern constraint default_io_commits_robIdx_6_flag_cons;
    extern constraint default_io_commits_robIdx_6_value_cons;
    extern constraint default_io_commits_robIdx_7_flag_cons;
    extern constraint default_io_commits_robIdx_7_value_cons;
    extern constraint default_io_trace_blockCommit_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_0_valid_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_0_bits_ftqOffset_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_1_valid_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_1_bits_ftqOffset_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_2_valid_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_2_bits_ftqOffset_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_3_valid_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_3_bits_ftqOffset_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_4_valid_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_4_bits_ftqOffset_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_5_valid_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_5_bits_ftqOffset_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_6_valid_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_6_bits_ftqOffset_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_7_valid_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_7_bits_ftqOffset_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire_cons;
    extern constraint default_io_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize_cons;
    extern constraint default_io_rabCommits_isCommit_cons;
    extern constraint default_io_rabCommits_commitValid_0_cons;
    extern constraint default_io_rabCommits_commitValid_1_cons;
    extern constraint default_io_rabCommits_commitValid_2_cons;
    extern constraint default_io_rabCommits_commitValid_3_cons;
    extern constraint default_io_rabCommits_commitValid_4_cons;
    extern constraint default_io_rabCommits_commitValid_5_cons;
    extern constraint default_io_rabCommits_isWalk_cons;
    extern constraint default_io_rabCommits_walkValid_0_cons;
    extern constraint default_io_rabCommits_walkValid_1_cons;
    extern constraint default_io_rabCommits_walkValid_2_cons;
    extern constraint default_io_rabCommits_walkValid_3_cons;
    extern constraint default_io_rabCommits_walkValid_4_cons;
    extern constraint default_io_rabCommits_walkValid_5_cons;
    extern constraint default_io_rabCommits_info_0_ldest_cons;
    extern constraint default_io_rabCommits_info_0_pdest_cons;
    extern constraint default_io_rabCommits_info_0_rfWen_cons;
    extern constraint default_io_rabCommits_info_0_fpWen_cons;
    extern constraint default_io_rabCommits_info_0_vecWen_cons;
    extern constraint default_io_rabCommits_info_0_v0Wen_cons;
    extern constraint default_io_rabCommits_info_0_vlWen_cons;
    extern constraint default_io_rabCommits_info_0_isMove_cons;
    extern constraint default_io_rabCommits_info_1_ldest_cons;
    extern constraint default_io_rabCommits_info_1_pdest_cons;
    extern constraint default_io_rabCommits_info_1_rfWen_cons;
    extern constraint default_io_rabCommits_info_1_fpWen_cons;
    extern constraint default_io_rabCommits_info_1_vecWen_cons;
    extern constraint default_io_rabCommits_info_1_v0Wen_cons;
    extern constraint default_io_rabCommits_info_1_vlWen_cons;
    extern constraint default_io_rabCommits_info_1_isMove_cons;
    extern constraint default_io_rabCommits_info_2_ldest_cons;
    extern constraint default_io_rabCommits_info_2_pdest_cons;
    extern constraint default_io_rabCommits_info_2_rfWen_cons;
    extern constraint default_io_rabCommits_info_2_fpWen_cons;
    extern constraint default_io_rabCommits_info_2_vecWen_cons;
    extern constraint default_io_rabCommits_info_2_v0Wen_cons;
    extern constraint default_io_rabCommits_info_2_vlWen_cons;
    extern constraint default_io_rabCommits_info_2_isMove_cons;
    extern constraint default_io_rabCommits_info_3_ldest_cons;
    extern constraint default_io_rabCommits_info_3_pdest_cons;
    extern constraint default_io_rabCommits_info_3_rfWen_cons;
    extern constraint default_io_rabCommits_info_3_fpWen_cons;
    extern constraint default_io_rabCommits_info_3_vecWen_cons;
    extern constraint default_io_rabCommits_info_3_v0Wen_cons;
    extern constraint default_io_rabCommits_info_3_vlWen_cons;
    extern constraint default_io_rabCommits_info_3_isMove_cons;
    extern constraint default_io_rabCommits_info_4_ldest_cons;
    extern constraint default_io_rabCommits_info_4_pdest_cons;
    extern constraint default_io_rabCommits_info_4_rfWen_cons;
    extern constraint default_io_rabCommits_info_4_fpWen_cons;
    extern constraint default_io_rabCommits_info_4_vecWen_cons;
    extern constraint default_io_rabCommits_info_4_v0Wen_cons;
    extern constraint default_io_rabCommits_info_4_vlWen_cons;
    extern constraint default_io_rabCommits_info_4_isMove_cons;
    extern constraint default_io_rabCommits_info_5_ldest_cons;
    extern constraint default_io_rabCommits_info_5_pdest_cons;
    extern constraint default_io_rabCommits_info_5_rfWen_cons;
    extern constraint default_io_rabCommits_info_5_fpWen_cons;
    extern constraint default_io_rabCommits_info_5_vecWen_cons;
    extern constraint default_io_rabCommits_info_5_v0Wen_cons;
    extern constraint default_io_rabCommits_info_5_vlWen_cons;
    extern constraint default_io_rabCommits_info_5_isMove_cons;
    extern constraint default_io_diffCommits_commitValid_0_cons;
    extern constraint default_io_diffCommits_commitValid_1_cons;
    extern constraint default_io_diffCommits_commitValid_2_cons;
    extern constraint default_io_diffCommits_commitValid_3_cons;
    extern constraint default_io_diffCommits_commitValid_4_cons;
    extern constraint default_io_diffCommits_commitValid_5_cons;
    extern constraint default_io_diffCommits_commitValid_6_cons;
    extern constraint default_io_diffCommits_commitValid_7_cons;
    extern constraint default_io_diffCommits_commitValid_8_cons;
    extern constraint default_io_diffCommits_commitValid_9_cons;
    extern constraint default_io_diffCommits_commitValid_10_cons;
    extern constraint default_io_diffCommits_commitValid_11_cons;
    extern constraint default_io_diffCommits_commitValid_12_cons;
    extern constraint default_io_diffCommits_commitValid_13_cons;
    extern constraint default_io_diffCommits_commitValid_14_cons;
    extern constraint default_io_diffCommits_commitValid_15_cons;
    extern constraint default_io_diffCommits_commitValid_16_cons;
    extern constraint default_io_diffCommits_commitValid_17_cons;
    extern constraint default_io_diffCommits_commitValid_18_cons;
    extern constraint default_io_diffCommits_commitValid_19_cons;
    extern constraint default_io_diffCommits_commitValid_20_cons;
    extern constraint default_io_diffCommits_commitValid_21_cons;
    extern constraint default_io_diffCommits_commitValid_22_cons;
    extern constraint default_io_diffCommits_commitValid_23_cons;
    extern constraint default_io_diffCommits_commitValid_24_cons;
    extern constraint default_io_diffCommits_commitValid_25_cons;
    extern constraint default_io_diffCommits_commitValid_26_cons;
    extern constraint default_io_diffCommits_commitValid_27_cons;
    extern constraint default_io_diffCommits_commitValid_28_cons;
    extern constraint default_io_diffCommits_commitValid_29_cons;
    extern constraint default_io_diffCommits_commitValid_30_cons;
    extern constraint default_io_diffCommits_commitValid_31_cons;
    extern constraint default_io_diffCommits_commitValid_32_cons;
    extern constraint default_io_diffCommits_commitValid_33_cons;
    extern constraint default_io_diffCommits_commitValid_34_cons;
    extern constraint default_io_diffCommits_commitValid_35_cons;
    extern constraint default_io_diffCommits_commitValid_36_cons;
    extern constraint default_io_diffCommits_commitValid_37_cons;
    extern constraint default_io_diffCommits_commitValid_38_cons;
    extern constraint default_io_diffCommits_commitValid_39_cons;
    extern constraint default_io_diffCommits_commitValid_40_cons;
    extern constraint default_io_diffCommits_commitValid_41_cons;
    extern constraint default_io_diffCommits_commitValid_42_cons;
    extern constraint default_io_diffCommits_commitValid_43_cons;
    extern constraint default_io_diffCommits_commitValid_44_cons;
    extern constraint default_io_diffCommits_commitValid_45_cons;
    extern constraint default_io_diffCommits_commitValid_46_cons;
    extern constraint default_io_diffCommits_commitValid_47_cons;
    extern constraint default_io_diffCommits_commitValid_48_cons;
    extern constraint default_io_diffCommits_commitValid_49_cons;
    extern constraint default_io_diffCommits_commitValid_50_cons;
    extern constraint default_io_diffCommits_commitValid_51_cons;
    extern constraint default_io_diffCommits_commitValid_52_cons;
    extern constraint default_io_diffCommits_commitValid_53_cons;
    extern constraint default_io_diffCommits_commitValid_54_cons;
    extern constraint default_io_diffCommits_commitValid_55_cons;
    extern constraint default_io_diffCommits_commitValid_56_cons;
    extern constraint default_io_diffCommits_commitValid_57_cons;
    extern constraint default_io_diffCommits_commitValid_58_cons;
    extern constraint default_io_diffCommits_commitValid_59_cons;
    extern constraint default_io_diffCommits_commitValid_60_cons;
    extern constraint default_io_diffCommits_commitValid_61_cons;
    extern constraint default_io_diffCommits_commitValid_62_cons;
    extern constraint default_io_diffCommits_commitValid_63_cons;
    extern constraint default_io_diffCommits_commitValid_64_cons;
    extern constraint default_io_diffCommits_commitValid_65_cons;
    extern constraint default_io_diffCommits_commitValid_66_cons;
    extern constraint default_io_diffCommits_commitValid_67_cons;
    extern constraint default_io_diffCommits_commitValid_68_cons;
    extern constraint default_io_diffCommits_commitValid_69_cons;
    extern constraint default_io_diffCommits_commitValid_70_cons;
    extern constraint default_io_diffCommits_commitValid_71_cons;
    extern constraint default_io_diffCommits_commitValid_72_cons;
    extern constraint default_io_diffCommits_commitValid_73_cons;
    extern constraint default_io_diffCommits_commitValid_74_cons;
    extern constraint default_io_diffCommits_commitValid_75_cons;
    extern constraint default_io_diffCommits_commitValid_76_cons;
    extern constraint default_io_diffCommits_commitValid_77_cons;
    extern constraint default_io_diffCommits_commitValid_78_cons;
    extern constraint default_io_diffCommits_commitValid_79_cons;
    extern constraint default_io_diffCommits_commitValid_80_cons;
    extern constraint default_io_diffCommits_commitValid_81_cons;
    extern constraint default_io_diffCommits_commitValid_82_cons;
    extern constraint default_io_diffCommits_commitValid_83_cons;
    extern constraint default_io_diffCommits_commitValid_84_cons;
    extern constraint default_io_diffCommits_commitValid_85_cons;
    extern constraint default_io_diffCommits_commitValid_86_cons;
    extern constraint default_io_diffCommits_commitValid_87_cons;
    extern constraint default_io_diffCommits_commitValid_88_cons;
    extern constraint default_io_diffCommits_commitValid_89_cons;
    extern constraint default_io_diffCommits_commitValid_90_cons;
    extern constraint default_io_diffCommits_commitValid_91_cons;
    extern constraint default_io_diffCommits_commitValid_92_cons;
    extern constraint default_io_diffCommits_commitValid_93_cons;
    extern constraint default_io_diffCommits_commitValid_94_cons;
    extern constraint default_io_diffCommits_commitValid_95_cons;
    extern constraint default_io_diffCommits_commitValid_96_cons;
    extern constraint default_io_diffCommits_commitValid_97_cons;
    extern constraint default_io_diffCommits_commitValid_98_cons;
    extern constraint default_io_diffCommits_commitValid_99_cons;
    extern constraint default_io_diffCommits_commitValid_100_cons;
    extern constraint default_io_diffCommits_commitValid_101_cons;
    extern constraint default_io_diffCommits_commitValid_102_cons;
    extern constraint default_io_diffCommits_commitValid_103_cons;
    extern constraint default_io_diffCommits_commitValid_104_cons;
    extern constraint default_io_diffCommits_commitValid_105_cons;
    extern constraint default_io_diffCommits_commitValid_106_cons;
    extern constraint default_io_diffCommits_commitValid_107_cons;
    extern constraint default_io_diffCommits_commitValid_108_cons;
    extern constraint default_io_diffCommits_commitValid_109_cons;
    extern constraint default_io_diffCommits_commitValid_110_cons;
    extern constraint default_io_diffCommits_commitValid_111_cons;
    extern constraint default_io_diffCommits_commitValid_112_cons;
    extern constraint default_io_diffCommits_commitValid_113_cons;
    extern constraint default_io_diffCommits_commitValid_114_cons;
    extern constraint default_io_diffCommits_commitValid_115_cons;
    extern constraint default_io_diffCommits_commitValid_116_cons;
    extern constraint default_io_diffCommits_commitValid_117_cons;
    extern constraint default_io_diffCommits_commitValid_118_cons;
    extern constraint default_io_diffCommits_commitValid_119_cons;
    extern constraint default_io_diffCommits_commitValid_120_cons;
    extern constraint default_io_diffCommits_commitValid_121_cons;
    extern constraint default_io_diffCommits_commitValid_122_cons;
    extern constraint default_io_diffCommits_commitValid_123_cons;
    extern constraint default_io_diffCommits_commitValid_124_cons;
    extern constraint default_io_diffCommits_commitValid_125_cons;
    extern constraint default_io_diffCommits_commitValid_126_cons;
    extern constraint default_io_diffCommits_commitValid_127_cons;
    extern constraint default_io_diffCommits_commitValid_128_cons;
    extern constraint default_io_diffCommits_commitValid_129_cons;
    extern constraint default_io_diffCommits_commitValid_130_cons;
    extern constraint default_io_diffCommits_commitValid_131_cons;
    extern constraint default_io_diffCommits_commitValid_132_cons;
    extern constraint default_io_diffCommits_commitValid_133_cons;
    extern constraint default_io_diffCommits_commitValid_134_cons;
    extern constraint default_io_diffCommits_commitValid_135_cons;
    extern constraint default_io_diffCommits_commitValid_136_cons;
    extern constraint default_io_diffCommits_commitValid_137_cons;
    extern constraint default_io_diffCommits_commitValid_138_cons;
    extern constraint default_io_diffCommits_commitValid_139_cons;
    extern constraint default_io_diffCommits_commitValid_140_cons;
    extern constraint default_io_diffCommits_commitValid_141_cons;
    extern constraint default_io_diffCommits_commitValid_142_cons;
    extern constraint default_io_diffCommits_commitValid_143_cons;
    extern constraint default_io_diffCommits_commitValid_144_cons;
    extern constraint default_io_diffCommits_commitValid_145_cons;
    extern constraint default_io_diffCommits_commitValid_146_cons;
    extern constraint default_io_diffCommits_commitValid_147_cons;
    extern constraint default_io_diffCommits_commitValid_148_cons;
    extern constraint default_io_diffCommits_commitValid_149_cons;
    extern constraint default_io_diffCommits_commitValid_150_cons;
    extern constraint default_io_diffCommits_commitValid_151_cons;
    extern constraint default_io_diffCommits_commitValid_152_cons;
    extern constraint default_io_diffCommits_commitValid_153_cons;
    extern constraint default_io_diffCommits_commitValid_154_cons;
    extern constraint default_io_diffCommits_commitValid_155_cons;
    extern constraint default_io_diffCommits_commitValid_156_cons;
    extern constraint default_io_diffCommits_commitValid_157_cons;
    extern constraint default_io_diffCommits_commitValid_158_cons;
    extern constraint default_io_diffCommits_commitValid_159_cons;
    extern constraint default_io_diffCommits_commitValid_160_cons;
    extern constraint default_io_diffCommits_commitValid_161_cons;
    extern constraint default_io_diffCommits_commitValid_162_cons;
    extern constraint default_io_diffCommits_commitValid_163_cons;
    extern constraint default_io_diffCommits_commitValid_164_cons;
    extern constraint default_io_diffCommits_commitValid_165_cons;
    extern constraint default_io_diffCommits_commitValid_166_cons;
    extern constraint default_io_diffCommits_commitValid_167_cons;
    extern constraint default_io_diffCommits_commitValid_168_cons;
    extern constraint default_io_diffCommits_commitValid_169_cons;
    extern constraint default_io_diffCommits_commitValid_170_cons;
    extern constraint default_io_diffCommits_commitValid_171_cons;
    extern constraint default_io_diffCommits_commitValid_172_cons;
    extern constraint default_io_diffCommits_commitValid_173_cons;
    extern constraint default_io_diffCommits_commitValid_174_cons;
    extern constraint default_io_diffCommits_commitValid_175_cons;
    extern constraint default_io_diffCommits_commitValid_176_cons;
    extern constraint default_io_diffCommits_commitValid_177_cons;
    extern constraint default_io_diffCommits_commitValid_178_cons;
    extern constraint default_io_diffCommits_commitValid_179_cons;
    extern constraint default_io_diffCommits_commitValid_180_cons;
    extern constraint default_io_diffCommits_commitValid_181_cons;
    extern constraint default_io_diffCommits_commitValid_182_cons;
    extern constraint default_io_diffCommits_commitValid_183_cons;
    extern constraint default_io_diffCommits_commitValid_184_cons;
    extern constraint default_io_diffCommits_commitValid_185_cons;
    extern constraint default_io_diffCommits_commitValid_186_cons;
    extern constraint default_io_diffCommits_commitValid_187_cons;
    extern constraint default_io_diffCommits_commitValid_188_cons;
    extern constraint default_io_diffCommits_commitValid_189_cons;
    extern constraint default_io_diffCommits_commitValid_190_cons;
    extern constraint default_io_diffCommits_commitValid_191_cons;
    extern constraint default_io_diffCommits_commitValid_192_cons;
    extern constraint default_io_diffCommits_commitValid_193_cons;
    extern constraint default_io_diffCommits_commitValid_194_cons;
    extern constraint default_io_diffCommits_commitValid_195_cons;
    extern constraint default_io_diffCommits_commitValid_196_cons;
    extern constraint default_io_diffCommits_commitValid_197_cons;
    extern constraint default_io_diffCommits_commitValid_198_cons;
    extern constraint default_io_diffCommits_commitValid_199_cons;
    extern constraint default_io_diffCommits_commitValid_200_cons;
    extern constraint default_io_diffCommits_commitValid_201_cons;
    extern constraint default_io_diffCommits_commitValid_202_cons;
    extern constraint default_io_diffCommits_commitValid_203_cons;
    extern constraint default_io_diffCommits_commitValid_204_cons;
    extern constraint default_io_diffCommits_commitValid_205_cons;
    extern constraint default_io_diffCommits_commitValid_206_cons;
    extern constraint default_io_diffCommits_commitValid_207_cons;
    extern constraint default_io_diffCommits_commitValid_208_cons;
    extern constraint default_io_diffCommits_commitValid_209_cons;
    extern constraint default_io_diffCommits_commitValid_210_cons;
    extern constraint default_io_diffCommits_commitValid_211_cons;
    extern constraint default_io_diffCommits_commitValid_212_cons;
    extern constraint default_io_diffCommits_commitValid_213_cons;
    extern constraint default_io_diffCommits_commitValid_214_cons;
    extern constraint default_io_diffCommits_commitValid_215_cons;
    extern constraint default_io_diffCommits_commitValid_216_cons;
    extern constraint default_io_diffCommits_commitValid_217_cons;
    extern constraint default_io_diffCommits_commitValid_218_cons;
    extern constraint default_io_diffCommits_commitValid_219_cons;
    extern constraint default_io_diffCommits_commitValid_220_cons;
    extern constraint default_io_diffCommits_commitValid_221_cons;
    extern constraint default_io_diffCommits_commitValid_222_cons;
    extern constraint default_io_diffCommits_commitValid_223_cons;
    extern constraint default_io_diffCommits_commitValid_224_cons;
    extern constraint default_io_diffCommits_commitValid_225_cons;
    extern constraint default_io_diffCommits_commitValid_226_cons;
    extern constraint default_io_diffCommits_commitValid_227_cons;
    extern constraint default_io_diffCommits_commitValid_228_cons;
    extern constraint default_io_diffCommits_commitValid_229_cons;
    extern constraint default_io_diffCommits_commitValid_230_cons;
    extern constraint default_io_diffCommits_commitValid_231_cons;
    extern constraint default_io_diffCommits_commitValid_232_cons;
    extern constraint default_io_diffCommits_commitValid_233_cons;
    extern constraint default_io_diffCommits_commitValid_234_cons;
    extern constraint default_io_diffCommits_commitValid_235_cons;
    extern constraint default_io_diffCommits_commitValid_236_cons;
    extern constraint default_io_diffCommits_commitValid_237_cons;
    extern constraint default_io_diffCommits_commitValid_238_cons;
    extern constraint default_io_diffCommits_commitValid_239_cons;
    extern constraint default_io_diffCommits_commitValid_240_cons;
    extern constraint default_io_diffCommits_commitValid_241_cons;
    extern constraint default_io_diffCommits_commitValid_242_cons;
    extern constraint default_io_diffCommits_commitValid_243_cons;
    extern constraint default_io_diffCommits_commitValid_244_cons;
    extern constraint default_io_diffCommits_commitValid_245_cons;
    extern constraint default_io_diffCommits_commitValid_246_cons;
    extern constraint default_io_diffCommits_commitValid_247_cons;
    extern constraint default_io_diffCommits_commitValid_248_cons;
    extern constraint default_io_diffCommits_commitValid_249_cons;
    extern constraint default_io_diffCommits_commitValid_250_cons;
    extern constraint default_io_diffCommits_commitValid_251_cons;
    extern constraint default_io_diffCommits_commitValid_252_cons;
    extern constraint default_io_diffCommits_commitValid_253_cons;
    extern constraint default_io_diffCommits_commitValid_254_cons;
    extern constraint default_io_diffCommits_info_0_ldest_cons;
    extern constraint default_io_diffCommits_info_0_pdest_cons;
    extern constraint default_io_diffCommits_info_0_rfWen_cons;
    extern constraint default_io_diffCommits_info_0_fpWen_cons;
    extern constraint default_io_diffCommits_info_0_vecWen_cons;
    extern constraint default_io_diffCommits_info_0_v0Wen_cons;
    extern constraint default_io_diffCommits_info_0_vlWen_cons;
    extern constraint default_io_diffCommits_info_1_ldest_cons;
    extern constraint default_io_diffCommits_info_1_pdest_cons;
    extern constraint default_io_diffCommits_info_1_rfWen_cons;
    extern constraint default_io_diffCommits_info_1_fpWen_cons;
    extern constraint default_io_diffCommits_info_1_vecWen_cons;
    extern constraint default_io_diffCommits_info_1_v0Wen_cons;
    extern constraint default_io_diffCommits_info_1_vlWen_cons;
    extern constraint default_io_diffCommits_info_2_ldest_cons;
    extern constraint default_io_diffCommits_info_2_pdest_cons;
    extern constraint default_io_diffCommits_info_2_rfWen_cons;
    extern constraint default_io_diffCommits_info_2_fpWen_cons;
    extern constraint default_io_diffCommits_info_2_vecWen_cons;
    extern constraint default_io_diffCommits_info_2_v0Wen_cons;
    extern constraint default_io_diffCommits_info_2_vlWen_cons;
    extern constraint default_io_diffCommits_info_3_ldest_cons;
    extern constraint default_io_diffCommits_info_3_pdest_cons;
    extern constraint default_io_diffCommits_info_3_rfWen_cons;
    extern constraint default_io_diffCommits_info_3_fpWen_cons;
    extern constraint default_io_diffCommits_info_3_vecWen_cons;
    extern constraint default_io_diffCommits_info_3_v0Wen_cons;
    extern constraint default_io_diffCommits_info_3_vlWen_cons;
    extern constraint default_io_diffCommits_info_4_ldest_cons;
    extern constraint default_io_diffCommits_info_4_pdest_cons;
    extern constraint default_io_diffCommits_info_4_rfWen_cons;
    extern constraint default_io_diffCommits_info_4_fpWen_cons;
    extern constraint default_io_diffCommits_info_4_vecWen_cons;
    extern constraint default_io_diffCommits_info_4_v0Wen_cons;
    extern constraint default_io_diffCommits_info_4_vlWen_cons;
    extern constraint default_io_diffCommits_info_5_ldest_cons;
    extern constraint default_io_diffCommits_info_5_pdest_cons;
    extern constraint default_io_diffCommits_info_5_rfWen_cons;
    extern constraint default_io_diffCommits_info_5_fpWen_cons;
    extern constraint default_io_diffCommits_info_5_vecWen_cons;
    extern constraint default_io_diffCommits_info_5_v0Wen_cons;
    extern constraint default_io_diffCommits_info_5_vlWen_cons;
    extern constraint default_io_diffCommits_info_6_ldest_cons;
    extern constraint default_io_diffCommits_info_6_pdest_cons;
    extern constraint default_io_diffCommits_info_6_rfWen_cons;
    extern constraint default_io_diffCommits_info_6_fpWen_cons;
    extern constraint default_io_diffCommits_info_6_vecWen_cons;
    extern constraint default_io_diffCommits_info_6_v0Wen_cons;
    extern constraint default_io_diffCommits_info_6_vlWen_cons;
    extern constraint default_io_diffCommits_info_7_ldest_cons;
    extern constraint default_io_diffCommits_info_7_pdest_cons;
    extern constraint default_io_diffCommits_info_7_rfWen_cons;
    extern constraint default_io_diffCommits_info_7_fpWen_cons;
    extern constraint default_io_diffCommits_info_7_vecWen_cons;
    extern constraint default_io_diffCommits_info_7_v0Wen_cons;
    extern constraint default_io_diffCommits_info_7_vlWen_cons;
    extern constraint default_io_diffCommits_info_8_ldest_cons;
    extern constraint default_io_diffCommits_info_8_pdest_cons;
    extern constraint default_io_diffCommits_info_8_rfWen_cons;
    extern constraint default_io_diffCommits_info_8_fpWen_cons;
    extern constraint default_io_diffCommits_info_8_vecWen_cons;
    extern constraint default_io_diffCommits_info_8_v0Wen_cons;
    extern constraint default_io_diffCommits_info_8_vlWen_cons;
    extern constraint default_io_diffCommits_info_9_ldest_cons;
    extern constraint default_io_diffCommits_info_9_pdest_cons;
    extern constraint default_io_diffCommits_info_9_rfWen_cons;
    extern constraint default_io_diffCommits_info_9_fpWen_cons;
    extern constraint default_io_diffCommits_info_9_vecWen_cons;
    extern constraint default_io_diffCommits_info_9_v0Wen_cons;
    extern constraint default_io_diffCommits_info_9_vlWen_cons;
    extern constraint default_io_diffCommits_info_10_ldest_cons;
    extern constraint default_io_diffCommits_info_10_pdest_cons;
    extern constraint default_io_diffCommits_info_10_rfWen_cons;
    extern constraint default_io_diffCommits_info_10_fpWen_cons;
    extern constraint default_io_diffCommits_info_10_vecWen_cons;
    extern constraint default_io_diffCommits_info_10_v0Wen_cons;
    extern constraint default_io_diffCommits_info_10_vlWen_cons;
    extern constraint default_io_diffCommits_info_11_ldest_cons;
    extern constraint default_io_diffCommits_info_11_pdest_cons;
    extern constraint default_io_diffCommits_info_11_rfWen_cons;
    extern constraint default_io_diffCommits_info_11_fpWen_cons;
    extern constraint default_io_diffCommits_info_11_vecWen_cons;
    extern constraint default_io_diffCommits_info_11_v0Wen_cons;
    extern constraint default_io_diffCommits_info_11_vlWen_cons;
    extern constraint default_io_diffCommits_info_12_ldest_cons;
    extern constraint default_io_diffCommits_info_12_pdest_cons;
    extern constraint default_io_diffCommits_info_12_rfWen_cons;
    extern constraint default_io_diffCommits_info_12_fpWen_cons;
    extern constraint default_io_diffCommits_info_12_vecWen_cons;
    extern constraint default_io_diffCommits_info_12_v0Wen_cons;
    extern constraint default_io_diffCommits_info_12_vlWen_cons;
    extern constraint default_io_diffCommits_info_13_ldest_cons;
    extern constraint default_io_diffCommits_info_13_pdest_cons;
    extern constraint default_io_diffCommits_info_13_rfWen_cons;
    extern constraint default_io_diffCommits_info_13_fpWen_cons;
    extern constraint default_io_diffCommits_info_13_vecWen_cons;
    extern constraint default_io_diffCommits_info_13_v0Wen_cons;
    extern constraint default_io_diffCommits_info_13_vlWen_cons;
    extern constraint default_io_diffCommits_info_14_ldest_cons;
    extern constraint default_io_diffCommits_info_14_pdest_cons;
    extern constraint default_io_diffCommits_info_14_rfWen_cons;
    extern constraint default_io_diffCommits_info_14_fpWen_cons;
    extern constraint default_io_diffCommits_info_14_vecWen_cons;
    extern constraint default_io_diffCommits_info_14_v0Wen_cons;
    extern constraint default_io_diffCommits_info_14_vlWen_cons;
    extern constraint default_io_diffCommits_info_15_ldest_cons;
    extern constraint default_io_diffCommits_info_15_pdest_cons;
    extern constraint default_io_diffCommits_info_15_rfWen_cons;
    extern constraint default_io_diffCommits_info_15_fpWen_cons;
    extern constraint default_io_diffCommits_info_15_vecWen_cons;
    extern constraint default_io_diffCommits_info_15_v0Wen_cons;
    extern constraint default_io_diffCommits_info_15_vlWen_cons;
    extern constraint default_io_diffCommits_info_16_ldest_cons;
    extern constraint default_io_diffCommits_info_16_pdest_cons;
    extern constraint default_io_diffCommits_info_16_rfWen_cons;
    extern constraint default_io_diffCommits_info_16_fpWen_cons;
    extern constraint default_io_diffCommits_info_16_vecWen_cons;
    extern constraint default_io_diffCommits_info_16_v0Wen_cons;
    extern constraint default_io_diffCommits_info_16_vlWen_cons;
    extern constraint default_io_diffCommits_info_17_ldest_cons;
    extern constraint default_io_diffCommits_info_17_pdest_cons;
    extern constraint default_io_diffCommits_info_17_rfWen_cons;
    extern constraint default_io_diffCommits_info_17_fpWen_cons;
    extern constraint default_io_diffCommits_info_17_vecWen_cons;
    extern constraint default_io_diffCommits_info_17_v0Wen_cons;
    extern constraint default_io_diffCommits_info_17_vlWen_cons;
    extern constraint default_io_diffCommits_info_18_ldest_cons;
    extern constraint default_io_diffCommits_info_18_pdest_cons;
    extern constraint default_io_diffCommits_info_18_rfWen_cons;
    extern constraint default_io_diffCommits_info_18_fpWen_cons;
    extern constraint default_io_diffCommits_info_18_vecWen_cons;
    extern constraint default_io_diffCommits_info_18_v0Wen_cons;
    extern constraint default_io_diffCommits_info_18_vlWen_cons;
    extern constraint default_io_diffCommits_info_19_ldest_cons;
    extern constraint default_io_diffCommits_info_19_pdest_cons;
    extern constraint default_io_diffCommits_info_19_rfWen_cons;
    extern constraint default_io_diffCommits_info_19_fpWen_cons;
    extern constraint default_io_diffCommits_info_19_vecWen_cons;
    extern constraint default_io_diffCommits_info_19_v0Wen_cons;
    extern constraint default_io_diffCommits_info_19_vlWen_cons;
    extern constraint default_io_diffCommits_info_20_ldest_cons;
    extern constraint default_io_diffCommits_info_20_pdest_cons;
    extern constraint default_io_diffCommits_info_20_rfWen_cons;
    extern constraint default_io_diffCommits_info_20_fpWen_cons;
    extern constraint default_io_diffCommits_info_20_vecWen_cons;
    extern constraint default_io_diffCommits_info_20_v0Wen_cons;
    extern constraint default_io_diffCommits_info_20_vlWen_cons;
    extern constraint default_io_diffCommits_info_21_ldest_cons;
    extern constraint default_io_diffCommits_info_21_pdest_cons;
    extern constraint default_io_diffCommits_info_21_rfWen_cons;
    extern constraint default_io_diffCommits_info_21_fpWen_cons;
    extern constraint default_io_diffCommits_info_21_vecWen_cons;
    extern constraint default_io_diffCommits_info_21_v0Wen_cons;
    extern constraint default_io_diffCommits_info_21_vlWen_cons;
    extern constraint default_io_diffCommits_info_22_ldest_cons;
    extern constraint default_io_diffCommits_info_22_pdest_cons;
    extern constraint default_io_diffCommits_info_22_rfWen_cons;
    extern constraint default_io_diffCommits_info_22_fpWen_cons;
    extern constraint default_io_diffCommits_info_22_vecWen_cons;
    extern constraint default_io_diffCommits_info_22_v0Wen_cons;
    extern constraint default_io_diffCommits_info_22_vlWen_cons;
    extern constraint default_io_diffCommits_info_23_ldest_cons;
    extern constraint default_io_diffCommits_info_23_pdest_cons;
    extern constraint default_io_diffCommits_info_23_rfWen_cons;
    extern constraint default_io_diffCommits_info_23_fpWen_cons;
    extern constraint default_io_diffCommits_info_23_vecWen_cons;
    extern constraint default_io_diffCommits_info_23_v0Wen_cons;
    extern constraint default_io_diffCommits_info_23_vlWen_cons;
    extern constraint default_io_diffCommits_info_24_ldest_cons;
    extern constraint default_io_diffCommits_info_24_pdest_cons;
    extern constraint default_io_diffCommits_info_24_rfWen_cons;
    extern constraint default_io_diffCommits_info_24_fpWen_cons;
    extern constraint default_io_diffCommits_info_24_vecWen_cons;
    extern constraint default_io_diffCommits_info_24_v0Wen_cons;
    extern constraint default_io_diffCommits_info_24_vlWen_cons;
    extern constraint default_io_diffCommits_info_25_ldest_cons;
    extern constraint default_io_diffCommits_info_25_pdest_cons;
    extern constraint default_io_diffCommits_info_25_rfWen_cons;
    extern constraint default_io_diffCommits_info_25_fpWen_cons;
    extern constraint default_io_diffCommits_info_25_vecWen_cons;
    extern constraint default_io_diffCommits_info_25_v0Wen_cons;
    extern constraint default_io_diffCommits_info_25_vlWen_cons;
    extern constraint default_io_diffCommits_info_26_ldest_cons;
    extern constraint default_io_diffCommits_info_26_pdest_cons;
    extern constraint default_io_diffCommits_info_26_rfWen_cons;
    extern constraint default_io_diffCommits_info_26_fpWen_cons;
    extern constraint default_io_diffCommits_info_26_vecWen_cons;
    extern constraint default_io_diffCommits_info_26_v0Wen_cons;
    extern constraint default_io_diffCommits_info_26_vlWen_cons;
    extern constraint default_io_diffCommits_info_27_ldest_cons;
    extern constraint default_io_diffCommits_info_27_pdest_cons;
    extern constraint default_io_diffCommits_info_27_rfWen_cons;
    extern constraint default_io_diffCommits_info_27_fpWen_cons;
    extern constraint default_io_diffCommits_info_27_vecWen_cons;
    extern constraint default_io_diffCommits_info_27_v0Wen_cons;
    extern constraint default_io_diffCommits_info_27_vlWen_cons;
    extern constraint default_io_diffCommits_info_28_ldest_cons;
    extern constraint default_io_diffCommits_info_28_pdest_cons;
    extern constraint default_io_diffCommits_info_28_rfWen_cons;
    extern constraint default_io_diffCommits_info_28_fpWen_cons;
    extern constraint default_io_diffCommits_info_28_vecWen_cons;
    extern constraint default_io_diffCommits_info_28_v0Wen_cons;
    extern constraint default_io_diffCommits_info_28_vlWen_cons;
    extern constraint default_io_diffCommits_info_29_ldest_cons;
    extern constraint default_io_diffCommits_info_29_pdest_cons;
    extern constraint default_io_diffCommits_info_29_rfWen_cons;
    extern constraint default_io_diffCommits_info_29_fpWen_cons;
    extern constraint default_io_diffCommits_info_29_vecWen_cons;
    extern constraint default_io_diffCommits_info_29_v0Wen_cons;
    extern constraint default_io_diffCommits_info_29_vlWen_cons;
    extern constraint default_io_diffCommits_info_30_ldest_cons;
    extern constraint default_io_diffCommits_info_30_pdest_cons;
    extern constraint default_io_diffCommits_info_30_rfWen_cons;
    extern constraint default_io_diffCommits_info_30_fpWen_cons;
    extern constraint default_io_diffCommits_info_30_vecWen_cons;
    extern constraint default_io_diffCommits_info_30_v0Wen_cons;
    extern constraint default_io_diffCommits_info_30_vlWen_cons;
    extern constraint default_io_diffCommits_info_31_ldest_cons;
    extern constraint default_io_diffCommits_info_31_pdest_cons;
    extern constraint default_io_diffCommits_info_31_rfWen_cons;
    extern constraint default_io_diffCommits_info_31_fpWen_cons;
    extern constraint default_io_diffCommits_info_31_vecWen_cons;
    extern constraint default_io_diffCommits_info_31_v0Wen_cons;
    extern constraint default_io_diffCommits_info_31_vlWen_cons;
    extern constraint default_io_diffCommits_info_32_ldest_cons;
    extern constraint default_io_diffCommits_info_32_pdest_cons;
    extern constraint default_io_diffCommits_info_32_rfWen_cons;
    extern constraint default_io_diffCommits_info_32_fpWen_cons;
    extern constraint default_io_diffCommits_info_32_vecWen_cons;
    extern constraint default_io_diffCommits_info_32_v0Wen_cons;
    extern constraint default_io_diffCommits_info_32_vlWen_cons;
    extern constraint default_io_diffCommits_info_33_ldest_cons;
    extern constraint default_io_diffCommits_info_33_pdest_cons;
    extern constraint default_io_diffCommits_info_33_rfWen_cons;
    extern constraint default_io_diffCommits_info_33_fpWen_cons;
    extern constraint default_io_diffCommits_info_33_vecWen_cons;
    extern constraint default_io_diffCommits_info_33_v0Wen_cons;
    extern constraint default_io_diffCommits_info_33_vlWen_cons;
    extern constraint default_io_diffCommits_info_34_ldest_cons;
    extern constraint default_io_diffCommits_info_34_pdest_cons;
    extern constraint default_io_diffCommits_info_34_rfWen_cons;
    extern constraint default_io_diffCommits_info_34_fpWen_cons;
    extern constraint default_io_diffCommits_info_34_vecWen_cons;
    extern constraint default_io_diffCommits_info_34_v0Wen_cons;
    extern constraint default_io_diffCommits_info_34_vlWen_cons;
    extern constraint default_io_diffCommits_info_35_ldest_cons;
    extern constraint default_io_diffCommits_info_35_pdest_cons;
    extern constraint default_io_diffCommits_info_35_rfWen_cons;
    extern constraint default_io_diffCommits_info_35_fpWen_cons;
    extern constraint default_io_diffCommits_info_35_vecWen_cons;
    extern constraint default_io_diffCommits_info_35_v0Wen_cons;
    extern constraint default_io_diffCommits_info_35_vlWen_cons;
    extern constraint default_io_diffCommits_info_36_ldest_cons;
    extern constraint default_io_diffCommits_info_36_pdest_cons;
    extern constraint default_io_diffCommits_info_36_rfWen_cons;
    extern constraint default_io_diffCommits_info_36_fpWen_cons;
    extern constraint default_io_diffCommits_info_36_vecWen_cons;
    extern constraint default_io_diffCommits_info_36_v0Wen_cons;
    extern constraint default_io_diffCommits_info_36_vlWen_cons;
    extern constraint default_io_diffCommits_info_37_ldest_cons;
    extern constraint default_io_diffCommits_info_37_pdest_cons;
    extern constraint default_io_diffCommits_info_37_rfWen_cons;
    extern constraint default_io_diffCommits_info_37_fpWen_cons;
    extern constraint default_io_diffCommits_info_37_vecWen_cons;
    extern constraint default_io_diffCommits_info_37_v0Wen_cons;
    extern constraint default_io_diffCommits_info_37_vlWen_cons;
    extern constraint default_io_diffCommits_info_38_ldest_cons;
    extern constraint default_io_diffCommits_info_38_pdest_cons;
    extern constraint default_io_diffCommits_info_38_rfWen_cons;
    extern constraint default_io_diffCommits_info_38_fpWen_cons;
    extern constraint default_io_diffCommits_info_38_vecWen_cons;
    extern constraint default_io_diffCommits_info_38_v0Wen_cons;
    extern constraint default_io_diffCommits_info_38_vlWen_cons;
    extern constraint default_io_diffCommits_info_39_ldest_cons;
    extern constraint default_io_diffCommits_info_39_pdest_cons;
    extern constraint default_io_diffCommits_info_39_rfWen_cons;
    extern constraint default_io_diffCommits_info_39_fpWen_cons;
    extern constraint default_io_diffCommits_info_39_vecWen_cons;
    extern constraint default_io_diffCommits_info_39_v0Wen_cons;
    extern constraint default_io_diffCommits_info_39_vlWen_cons;
    extern constraint default_io_diffCommits_info_40_ldest_cons;
    extern constraint default_io_diffCommits_info_40_pdest_cons;
    extern constraint default_io_diffCommits_info_40_rfWen_cons;
    extern constraint default_io_diffCommits_info_40_fpWen_cons;
    extern constraint default_io_diffCommits_info_40_vecWen_cons;
    extern constraint default_io_diffCommits_info_40_v0Wen_cons;
    extern constraint default_io_diffCommits_info_40_vlWen_cons;
    extern constraint default_io_diffCommits_info_41_ldest_cons;
    extern constraint default_io_diffCommits_info_41_pdest_cons;
    extern constraint default_io_diffCommits_info_41_rfWen_cons;
    extern constraint default_io_diffCommits_info_41_fpWen_cons;
    extern constraint default_io_diffCommits_info_41_vecWen_cons;
    extern constraint default_io_diffCommits_info_41_v0Wen_cons;
    extern constraint default_io_diffCommits_info_41_vlWen_cons;
    extern constraint default_io_diffCommits_info_42_ldest_cons;
    extern constraint default_io_diffCommits_info_42_pdest_cons;
    extern constraint default_io_diffCommits_info_42_rfWen_cons;
    extern constraint default_io_diffCommits_info_42_fpWen_cons;
    extern constraint default_io_diffCommits_info_42_vecWen_cons;
    extern constraint default_io_diffCommits_info_42_v0Wen_cons;
    extern constraint default_io_diffCommits_info_42_vlWen_cons;
    extern constraint default_io_diffCommits_info_43_ldest_cons;
    extern constraint default_io_diffCommits_info_43_pdest_cons;
    extern constraint default_io_diffCommits_info_43_rfWen_cons;
    extern constraint default_io_diffCommits_info_43_fpWen_cons;
    extern constraint default_io_diffCommits_info_43_vecWen_cons;
    extern constraint default_io_diffCommits_info_43_v0Wen_cons;
    extern constraint default_io_diffCommits_info_43_vlWen_cons;
    extern constraint default_io_diffCommits_info_44_ldest_cons;
    extern constraint default_io_diffCommits_info_44_pdest_cons;
    extern constraint default_io_diffCommits_info_44_rfWen_cons;
    extern constraint default_io_diffCommits_info_44_fpWen_cons;
    extern constraint default_io_diffCommits_info_44_vecWen_cons;
    extern constraint default_io_diffCommits_info_44_v0Wen_cons;
    extern constraint default_io_diffCommits_info_44_vlWen_cons;
    extern constraint default_io_diffCommits_info_45_ldest_cons;
    extern constraint default_io_diffCommits_info_45_pdest_cons;
    extern constraint default_io_diffCommits_info_45_rfWen_cons;
    extern constraint default_io_diffCommits_info_45_fpWen_cons;
    extern constraint default_io_diffCommits_info_45_vecWen_cons;
    extern constraint default_io_diffCommits_info_45_v0Wen_cons;
    extern constraint default_io_diffCommits_info_45_vlWen_cons;
    extern constraint default_io_diffCommits_info_46_ldest_cons;
    extern constraint default_io_diffCommits_info_46_pdest_cons;
    extern constraint default_io_diffCommits_info_46_rfWen_cons;
    extern constraint default_io_diffCommits_info_46_fpWen_cons;
    extern constraint default_io_diffCommits_info_46_vecWen_cons;
    extern constraint default_io_diffCommits_info_46_v0Wen_cons;
    extern constraint default_io_diffCommits_info_46_vlWen_cons;
    extern constraint default_io_diffCommits_info_47_ldest_cons;
    extern constraint default_io_diffCommits_info_47_pdest_cons;
    extern constraint default_io_diffCommits_info_47_rfWen_cons;
    extern constraint default_io_diffCommits_info_47_fpWen_cons;
    extern constraint default_io_diffCommits_info_47_vecWen_cons;
    extern constraint default_io_diffCommits_info_47_v0Wen_cons;
    extern constraint default_io_diffCommits_info_47_vlWen_cons;
    extern constraint default_io_diffCommits_info_48_ldest_cons;
    extern constraint default_io_diffCommits_info_48_pdest_cons;
    extern constraint default_io_diffCommits_info_48_rfWen_cons;
    extern constraint default_io_diffCommits_info_48_fpWen_cons;
    extern constraint default_io_diffCommits_info_48_vecWen_cons;
    extern constraint default_io_diffCommits_info_48_v0Wen_cons;
    extern constraint default_io_diffCommits_info_48_vlWen_cons;
    extern constraint default_io_diffCommits_info_49_ldest_cons;
    extern constraint default_io_diffCommits_info_49_pdest_cons;
    extern constraint default_io_diffCommits_info_49_rfWen_cons;
    extern constraint default_io_diffCommits_info_49_fpWen_cons;
    extern constraint default_io_diffCommits_info_49_vecWen_cons;
    extern constraint default_io_diffCommits_info_49_v0Wen_cons;
    extern constraint default_io_diffCommits_info_49_vlWen_cons;
    extern constraint default_io_diffCommits_info_50_ldest_cons;
    extern constraint default_io_diffCommits_info_50_pdest_cons;
    extern constraint default_io_diffCommits_info_50_rfWen_cons;
    extern constraint default_io_diffCommits_info_50_fpWen_cons;
    extern constraint default_io_diffCommits_info_50_vecWen_cons;
    extern constraint default_io_diffCommits_info_50_v0Wen_cons;
    extern constraint default_io_diffCommits_info_50_vlWen_cons;
    extern constraint default_io_diffCommits_info_51_ldest_cons;
    extern constraint default_io_diffCommits_info_51_pdest_cons;
    extern constraint default_io_diffCommits_info_51_rfWen_cons;
    extern constraint default_io_diffCommits_info_51_fpWen_cons;
    extern constraint default_io_diffCommits_info_51_vecWen_cons;
    extern constraint default_io_diffCommits_info_51_v0Wen_cons;
    extern constraint default_io_diffCommits_info_51_vlWen_cons;
    extern constraint default_io_diffCommits_info_52_ldest_cons;
    extern constraint default_io_diffCommits_info_52_pdest_cons;
    extern constraint default_io_diffCommits_info_52_rfWen_cons;
    extern constraint default_io_diffCommits_info_52_fpWen_cons;
    extern constraint default_io_diffCommits_info_52_vecWen_cons;
    extern constraint default_io_diffCommits_info_52_v0Wen_cons;
    extern constraint default_io_diffCommits_info_52_vlWen_cons;
    extern constraint default_io_diffCommits_info_53_ldest_cons;
    extern constraint default_io_diffCommits_info_53_pdest_cons;
    extern constraint default_io_diffCommits_info_53_rfWen_cons;
    extern constraint default_io_diffCommits_info_53_fpWen_cons;
    extern constraint default_io_diffCommits_info_53_vecWen_cons;
    extern constraint default_io_diffCommits_info_53_v0Wen_cons;
    extern constraint default_io_diffCommits_info_53_vlWen_cons;
    extern constraint default_io_diffCommits_info_54_ldest_cons;
    extern constraint default_io_diffCommits_info_54_pdest_cons;
    extern constraint default_io_diffCommits_info_54_rfWen_cons;
    extern constraint default_io_diffCommits_info_54_fpWen_cons;
    extern constraint default_io_diffCommits_info_54_vecWen_cons;
    extern constraint default_io_diffCommits_info_54_v0Wen_cons;
    extern constraint default_io_diffCommits_info_54_vlWen_cons;
    extern constraint default_io_diffCommits_info_55_ldest_cons;
    extern constraint default_io_diffCommits_info_55_pdest_cons;
    extern constraint default_io_diffCommits_info_55_rfWen_cons;
    extern constraint default_io_diffCommits_info_55_fpWen_cons;
    extern constraint default_io_diffCommits_info_55_vecWen_cons;
    extern constraint default_io_diffCommits_info_55_v0Wen_cons;
    extern constraint default_io_diffCommits_info_55_vlWen_cons;
    extern constraint default_io_diffCommits_info_56_ldest_cons;
    extern constraint default_io_diffCommits_info_56_pdest_cons;
    extern constraint default_io_diffCommits_info_56_rfWen_cons;
    extern constraint default_io_diffCommits_info_56_fpWen_cons;
    extern constraint default_io_diffCommits_info_56_vecWen_cons;
    extern constraint default_io_diffCommits_info_56_v0Wen_cons;
    extern constraint default_io_diffCommits_info_56_vlWen_cons;
    extern constraint default_io_diffCommits_info_57_ldest_cons;
    extern constraint default_io_diffCommits_info_57_pdest_cons;
    extern constraint default_io_diffCommits_info_57_rfWen_cons;
    extern constraint default_io_diffCommits_info_57_fpWen_cons;
    extern constraint default_io_diffCommits_info_57_vecWen_cons;
    extern constraint default_io_diffCommits_info_57_v0Wen_cons;
    extern constraint default_io_diffCommits_info_57_vlWen_cons;
    extern constraint default_io_diffCommits_info_58_ldest_cons;
    extern constraint default_io_diffCommits_info_58_pdest_cons;
    extern constraint default_io_diffCommits_info_58_rfWen_cons;
    extern constraint default_io_diffCommits_info_58_fpWen_cons;
    extern constraint default_io_diffCommits_info_58_vecWen_cons;
    extern constraint default_io_diffCommits_info_58_v0Wen_cons;
    extern constraint default_io_diffCommits_info_58_vlWen_cons;
    extern constraint default_io_diffCommits_info_59_ldest_cons;
    extern constraint default_io_diffCommits_info_59_pdest_cons;
    extern constraint default_io_diffCommits_info_59_rfWen_cons;
    extern constraint default_io_diffCommits_info_59_fpWen_cons;
    extern constraint default_io_diffCommits_info_59_vecWen_cons;
    extern constraint default_io_diffCommits_info_59_v0Wen_cons;
    extern constraint default_io_diffCommits_info_59_vlWen_cons;
    extern constraint default_io_diffCommits_info_60_ldest_cons;
    extern constraint default_io_diffCommits_info_60_pdest_cons;
    extern constraint default_io_diffCommits_info_60_rfWen_cons;
    extern constraint default_io_diffCommits_info_60_fpWen_cons;
    extern constraint default_io_diffCommits_info_60_vecWen_cons;
    extern constraint default_io_diffCommits_info_60_v0Wen_cons;
    extern constraint default_io_diffCommits_info_60_vlWen_cons;
    extern constraint default_io_diffCommits_info_61_ldest_cons;
    extern constraint default_io_diffCommits_info_61_pdest_cons;
    extern constraint default_io_diffCommits_info_61_rfWen_cons;
    extern constraint default_io_diffCommits_info_61_fpWen_cons;
    extern constraint default_io_diffCommits_info_61_vecWen_cons;
    extern constraint default_io_diffCommits_info_61_v0Wen_cons;
    extern constraint default_io_diffCommits_info_61_vlWen_cons;
    extern constraint default_io_diffCommits_info_62_ldest_cons;
    extern constraint default_io_diffCommits_info_62_pdest_cons;
    extern constraint default_io_diffCommits_info_62_rfWen_cons;
    extern constraint default_io_diffCommits_info_62_fpWen_cons;
    extern constraint default_io_diffCommits_info_62_vecWen_cons;
    extern constraint default_io_diffCommits_info_62_v0Wen_cons;
    extern constraint default_io_diffCommits_info_62_vlWen_cons;
    extern constraint default_io_diffCommits_info_63_ldest_cons;
    extern constraint default_io_diffCommits_info_63_pdest_cons;
    extern constraint default_io_diffCommits_info_63_rfWen_cons;
    extern constraint default_io_diffCommits_info_63_fpWen_cons;
    extern constraint default_io_diffCommits_info_63_vecWen_cons;
    extern constraint default_io_diffCommits_info_63_v0Wen_cons;
    extern constraint default_io_diffCommits_info_63_vlWen_cons;
    extern constraint default_io_diffCommits_info_64_ldest_cons;
    extern constraint default_io_diffCommits_info_64_pdest_cons;
    extern constraint default_io_diffCommits_info_64_rfWen_cons;
    extern constraint default_io_diffCommits_info_64_fpWen_cons;
    extern constraint default_io_diffCommits_info_64_vecWen_cons;
    extern constraint default_io_diffCommits_info_64_v0Wen_cons;
    extern constraint default_io_diffCommits_info_64_vlWen_cons;
    extern constraint default_io_diffCommits_info_65_ldest_cons;
    extern constraint default_io_diffCommits_info_65_pdest_cons;
    extern constraint default_io_diffCommits_info_65_rfWen_cons;
    extern constraint default_io_diffCommits_info_65_fpWen_cons;
    extern constraint default_io_diffCommits_info_65_vecWen_cons;
    extern constraint default_io_diffCommits_info_65_v0Wen_cons;
    extern constraint default_io_diffCommits_info_65_vlWen_cons;
    extern constraint default_io_diffCommits_info_66_ldest_cons;
    extern constraint default_io_diffCommits_info_66_pdest_cons;
    extern constraint default_io_diffCommits_info_66_rfWen_cons;
    extern constraint default_io_diffCommits_info_66_fpWen_cons;
    extern constraint default_io_diffCommits_info_66_vecWen_cons;
    extern constraint default_io_diffCommits_info_66_v0Wen_cons;
    extern constraint default_io_diffCommits_info_66_vlWen_cons;
    extern constraint default_io_diffCommits_info_67_ldest_cons;
    extern constraint default_io_diffCommits_info_67_pdest_cons;
    extern constraint default_io_diffCommits_info_67_rfWen_cons;
    extern constraint default_io_diffCommits_info_67_fpWen_cons;
    extern constraint default_io_diffCommits_info_67_vecWen_cons;
    extern constraint default_io_diffCommits_info_67_v0Wen_cons;
    extern constraint default_io_diffCommits_info_67_vlWen_cons;
    extern constraint default_io_diffCommits_info_68_ldest_cons;
    extern constraint default_io_diffCommits_info_68_pdest_cons;
    extern constraint default_io_diffCommits_info_68_rfWen_cons;
    extern constraint default_io_diffCommits_info_68_fpWen_cons;
    extern constraint default_io_diffCommits_info_68_vecWen_cons;
    extern constraint default_io_diffCommits_info_68_v0Wen_cons;
    extern constraint default_io_diffCommits_info_68_vlWen_cons;
    extern constraint default_io_diffCommits_info_69_ldest_cons;
    extern constraint default_io_diffCommits_info_69_pdest_cons;
    extern constraint default_io_diffCommits_info_69_rfWen_cons;
    extern constraint default_io_diffCommits_info_69_fpWen_cons;
    extern constraint default_io_diffCommits_info_69_vecWen_cons;
    extern constraint default_io_diffCommits_info_69_v0Wen_cons;
    extern constraint default_io_diffCommits_info_69_vlWen_cons;
    extern constraint default_io_diffCommits_info_70_ldest_cons;
    extern constraint default_io_diffCommits_info_70_pdest_cons;
    extern constraint default_io_diffCommits_info_70_rfWen_cons;
    extern constraint default_io_diffCommits_info_70_fpWen_cons;
    extern constraint default_io_diffCommits_info_70_vecWen_cons;
    extern constraint default_io_diffCommits_info_70_v0Wen_cons;
    extern constraint default_io_diffCommits_info_70_vlWen_cons;
    extern constraint default_io_diffCommits_info_71_ldest_cons;
    extern constraint default_io_diffCommits_info_71_pdest_cons;
    extern constraint default_io_diffCommits_info_71_rfWen_cons;
    extern constraint default_io_diffCommits_info_71_fpWen_cons;
    extern constraint default_io_diffCommits_info_71_vecWen_cons;
    extern constraint default_io_diffCommits_info_71_v0Wen_cons;
    extern constraint default_io_diffCommits_info_71_vlWen_cons;
    extern constraint default_io_diffCommits_info_72_ldest_cons;
    extern constraint default_io_diffCommits_info_72_pdest_cons;
    extern constraint default_io_diffCommits_info_72_rfWen_cons;
    extern constraint default_io_diffCommits_info_72_fpWen_cons;
    extern constraint default_io_diffCommits_info_72_vecWen_cons;
    extern constraint default_io_diffCommits_info_72_v0Wen_cons;
    extern constraint default_io_diffCommits_info_72_vlWen_cons;
    extern constraint default_io_diffCommits_info_73_ldest_cons;
    extern constraint default_io_diffCommits_info_73_pdest_cons;
    extern constraint default_io_diffCommits_info_73_rfWen_cons;
    extern constraint default_io_diffCommits_info_73_fpWen_cons;
    extern constraint default_io_diffCommits_info_73_vecWen_cons;
    extern constraint default_io_diffCommits_info_73_v0Wen_cons;
    extern constraint default_io_diffCommits_info_73_vlWen_cons;
    extern constraint default_io_diffCommits_info_74_ldest_cons;
    extern constraint default_io_diffCommits_info_74_pdest_cons;
    extern constraint default_io_diffCommits_info_74_rfWen_cons;
    extern constraint default_io_diffCommits_info_74_fpWen_cons;
    extern constraint default_io_diffCommits_info_74_vecWen_cons;
    extern constraint default_io_diffCommits_info_74_v0Wen_cons;
    extern constraint default_io_diffCommits_info_74_vlWen_cons;
    extern constraint default_io_diffCommits_info_75_ldest_cons;
    extern constraint default_io_diffCommits_info_75_pdest_cons;
    extern constraint default_io_diffCommits_info_75_rfWen_cons;
    extern constraint default_io_diffCommits_info_75_fpWen_cons;
    extern constraint default_io_diffCommits_info_75_vecWen_cons;
    extern constraint default_io_diffCommits_info_75_v0Wen_cons;
    extern constraint default_io_diffCommits_info_75_vlWen_cons;
    extern constraint default_io_diffCommits_info_76_ldest_cons;
    extern constraint default_io_diffCommits_info_76_pdest_cons;
    extern constraint default_io_diffCommits_info_76_rfWen_cons;
    extern constraint default_io_diffCommits_info_76_fpWen_cons;
    extern constraint default_io_diffCommits_info_76_vecWen_cons;
    extern constraint default_io_diffCommits_info_76_v0Wen_cons;
    extern constraint default_io_diffCommits_info_76_vlWen_cons;
    extern constraint default_io_diffCommits_info_77_ldest_cons;
    extern constraint default_io_diffCommits_info_77_pdest_cons;
    extern constraint default_io_diffCommits_info_77_rfWen_cons;
    extern constraint default_io_diffCommits_info_77_fpWen_cons;
    extern constraint default_io_diffCommits_info_77_vecWen_cons;
    extern constraint default_io_diffCommits_info_77_v0Wen_cons;
    extern constraint default_io_diffCommits_info_77_vlWen_cons;
    extern constraint default_io_diffCommits_info_78_ldest_cons;
    extern constraint default_io_diffCommits_info_78_pdest_cons;
    extern constraint default_io_diffCommits_info_78_rfWen_cons;
    extern constraint default_io_diffCommits_info_78_fpWen_cons;
    extern constraint default_io_diffCommits_info_78_vecWen_cons;
    extern constraint default_io_diffCommits_info_78_v0Wen_cons;
    extern constraint default_io_diffCommits_info_78_vlWen_cons;
    extern constraint default_io_diffCommits_info_79_ldest_cons;
    extern constraint default_io_diffCommits_info_79_pdest_cons;
    extern constraint default_io_diffCommits_info_79_rfWen_cons;
    extern constraint default_io_diffCommits_info_79_fpWen_cons;
    extern constraint default_io_diffCommits_info_79_vecWen_cons;
    extern constraint default_io_diffCommits_info_79_v0Wen_cons;
    extern constraint default_io_diffCommits_info_79_vlWen_cons;
    extern constraint default_io_diffCommits_info_80_ldest_cons;
    extern constraint default_io_diffCommits_info_80_pdest_cons;
    extern constraint default_io_diffCommits_info_80_rfWen_cons;
    extern constraint default_io_diffCommits_info_80_fpWen_cons;
    extern constraint default_io_diffCommits_info_80_vecWen_cons;
    extern constraint default_io_diffCommits_info_80_v0Wen_cons;
    extern constraint default_io_diffCommits_info_80_vlWen_cons;
    extern constraint default_io_diffCommits_info_81_ldest_cons;
    extern constraint default_io_diffCommits_info_81_pdest_cons;
    extern constraint default_io_diffCommits_info_81_rfWen_cons;
    extern constraint default_io_diffCommits_info_81_fpWen_cons;
    extern constraint default_io_diffCommits_info_81_vecWen_cons;
    extern constraint default_io_diffCommits_info_81_v0Wen_cons;
    extern constraint default_io_diffCommits_info_81_vlWen_cons;
    extern constraint default_io_diffCommits_info_82_ldest_cons;
    extern constraint default_io_diffCommits_info_82_pdest_cons;
    extern constraint default_io_diffCommits_info_82_rfWen_cons;
    extern constraint default_io_diffCommits_info_82_fpWen_cons;
    extern constraint default_io_diffCommits_info_82_vecWen_cons;
    extern constraint default_io_diffCommits_info_82_v0Wen_cons;
    extern constraint default_io_diffCommits_info_82_vlWen_cons;
    extern constraint default_io_diffCommits_info_83_ldest_cons;
    extern constraint default_io_diffCommits_info_83_pdest_cons;
    extern constraint default_io_diffCommits_info_83_rfWen_cons;
    extern constraint default_io_diffCommits_info_83_fpWen_cons;
    extern constraint default_io_diffCommits_info_83_vecWen_cons;
    extern constraint default_io_diffCommits_info_83_v0Wen_cons;
    extern constraint default_io_diffCommits_info_83_vlWen_cons;
    extern constraint default_io_diffCommits_info_84_ldest_cons;
    extern constraint default_io_diffCommits_info_84_pdest_cons;
    extern constraint default_io_diffCommits_info_84_rfWen_cons;
    extern constraint default_io_diffCommits_info_84_fpWen_cons;
    extern constraint default_io_diffCommits_info_84_vecWen_cons;
    extern constraint default_io_diffCommits_info_84_v0Wen_cons;
    extern constraint default_io_diffCommits_info_84_vlWen_cons;
    extern constraint default_io_diffCommits_info_85_ldest_cons;
    extern constraint default_io_diffCommits_info_85_pdest_cons;
    extern constraint default_io_diffCommits_info_85_rfWen_cons;
    extern constraint default_io_diffCommits_info_85_fpWen_cons;
    extern constraint default_io_diffCommits_info_85_vecWen_cons;
    extern constraint default_io_diffCommits_info_85_v0Wen_cons;
    extern constraint default_io_diffCommits_info_85_vlWen_cons;
    extern constraint default_io_diffCommits_info_86_ldest_cons;
    extern constraint default_io_diffCommits_info_86_pdest_cons;
    extern constraint default_io_diffCommits_info_86_rfWen_cons;
    extern constraint default_io_diffCommits_info_86_fpWen_cons;
    extern constraint default_io_diffCommits_info_86_vecWen_cons;
    extern constraint default_io_diffCommits_info_86_v0Wen_cons;
    extern constraint default_io_diffCommits_info_86_vlWen_cons;
    extern constraint default_io_diffCommits_info_87_ldest_cons;
    extern constraint default_io_diffCommits_info_87_pdest_cons;
    extern constraint default_io_diffCommits_info_87_rfWen_cons;
    extern constraint default_io_diffCommits_info_87_fpWen_cons;
    extern constraint default_io_diffCommits_info_87_vecWen_cons;
    extern constraint default_io_diffCommits_info_87_v0Wen_cons;
    extern constraint default_io_diffCommits_info_87_vlWen_cons;
    extern constraint default_io_diffCommits_info_88_ldest_cons;
    extern constraint default_io_diffCommits_info_88_pdest_cons;
    extern constraint default_io_diffCommits_info_88_rfWen_cons;
    extern constraint default_io_diffCommits_info_88_fpWen_cons;
    extern constraint default_io_diffCommits_info_88_vecWen_cons;
    extern constraint default_io_diffCommits_info_88_v0Wen_cons;
    extern constraint default_io_diffCommits_info_88_vlWen_cons;
    extern constraint default_io_diffCommits_info_89_ldest_cons;
    extern constraint default_io_diffCommits_info_89_pdest_cons;
    extern constraint default_io_diffCommits_info_89_rfWen_cons;
    extern constraint default_io_diffCommits_info_89_fpWen_cons;
    extern constraint default_io_diffCommits_info_89_vecWen_cons;
    extern constraint default_io_diffCommits_info_89_v0Wen_cons;
    extern constraint default_io_diffCommits_info_89_vlWen_cons;
    extern constraint default_io_diffCommits_info_90_ldest_cons;
    extern constraint default_io_diffCommits_info_90_pdest_cons;
    extern constraint default_io_diffCommits_info_90_rfWen_cons;
    extern constraint default_io_diffCommits_info_90_fpWen_cons;
    extern constraint default_io_diffCommits_info_90_vecWen_cons;
    extern constraint default_io_diffCommits_info_90_v0Wen_cons;
    extern constraint default_io_diffCommits_info_90_vlWen_cons;
    extern constraint default_io_diffCommits_info_91_ldest_cons;
    extern constraint default_io_diffCommits_info_91_pdest_cons;
    extern constraint default_io_diffCommits_info_91_rfWen_cons;
    extern constraint default_io_diffCommits_info_91_fpWen_cons;
    extern constraint default_io_diffCommits_info_91_vecWen_cons;
    extern constraint default_io_diffCommits_info_91_v0Wen_cons;
    extern constraint default_io_diffCommits_info_91_vlWen_cons;
    extern constraint default_io_diffCommits_info_92_ldest_cons;
    extern constraint default_io_diffCommits_info_92_pdest_cons;
    extern constraint default_io_diffCommits_info_92_rfWen_cons;
    extern constraint default_io_diffCommits_info_92_fpWen_cons;
    extern constraint default_io_diffCommits_info_92_vecWen_cons;
    extern constraint default_io_diffCommits_info_92_v0Wen_cons;
    extern constraint default_io_diffCommits_info_92_vlWen_cons;
    extern constraint default_io_diffCommits_info_93_ldest_cons;
    extern constraint default_io_diffCommits_info_93_pdest_cons;
    extern constraint default_io_diffCommits_info_93_rfWen_cons;
    extern constraint default_io_diffCommits_info_93_fpWen_cons;
    extern constraint default_io_diffCommits_info_93_vecWen_cons;
    extern constraint default_io_diffCommits_info_93_v0Wen_cons;
    extern constraint default_io_diffCommits_info_93_vlWen_cons;
    extern constraint default_io_diffCommits_info_94_ldest_cons;
    extern constraint default_io_diffCommits_info_94_pdest_cons;
    extern constraint default_io_diffCommits_info_94_rfWen_cons;
    extern constraint default_io_diffCommits_info_94_fpWen_cons;
    extern constraint default_io_diffCommits_info_94_vecWen_cons;
    extern constraint default_io_diffCommits_info_94_v0Wen_cons;
    extern constraint default_io_diffCommits_info_94_vlWen_cons;
    extern constraint default_io_diffCommits_info_95_ldest_cons;
    extern constraint default_io_diffCommits_info_95_pdest_cons;
    extern constraint default_io_diffCommits_info_95_rfWen_cons;
    extern constraint default_io_diffCommits_info_95_fpWen_cons;
    extern constraint default_io_diffCommits_info_95_vecWen_cons;
    extern constraint default_io_diffCommits_info_95_v0Wen_cons;
    extern constraint default_io_diffCommits_info_95_vlWen_cons;
    extern constraint default_io_diffCommits_info_96_ldest_cons;
    extern constraint default_io_diffCommits_info_96_pdest_cons;
    extern constraint default_io_diffCommits_info_96_rfWen_cons;
    extern constraint default_io_diffCommits_info_96_fpWen_cons;
    extern constraint default_io_diffCommits_info_96_vecWen_cons;
    extern constraint default_io_diffCommits_info_96_v0Wen_cons;
    extern constraint default_io_diffCommits_info_96_vlWen_cons;
    extern constraint default_io_diffCommits_info_97_ldest_cons;
    extern constraint default_io_diffCommits_info_97_pdest_cons;
    extern constraint default_io_diffCommits_info_97_rfWen_cons;
    extern constraint default_io_diffCommits_info_97_fpWen_cons;
    extern constraint default_io_diffCommits_info_97_vecWen_cons;
    extern constraint default_io_diffCommits_info_97_v0Wen_cons;
    extern constraint default_io_diffCommits_info_97_vlWen_cons;
    extern constraint default_io_diffCommits_info_98_ldest_cons;
    extern constraint default_io_diffCommits_info_98_pdest_cons;
    extern constraint default_io_diffCommits_info_98_rfWen_cons;
    extern constraint default_io_diffCommits_info_98_fpWen_cons;
    extern constraint default_io_diffCommits_info_98_vecWen_cons;
    extern constraint default_io_diffCommits_info_98_v0Wen_cons;
    extern constraint default_io_diffCommits_info_98_vlWen_cons;
    extern constraint default_io_diffCommits_info_99_ldest_cons;
    extern constraint default_io_diffCommits_info_99_pdest_cons;
    extern constraint default_io_diffCommits_info_99_rfWen_cons;
    extern constraint default_io_diffCommits_info_99_fpWen_cons;
    extern constraint default_io_diffCommits_info_99_vecWen_cons;
    extern constraint default_io_diffCommits_info_99_v0Wen_cons;
    extern constraint default_io_diffCommits_info_99_vlWen_cons;
    extern constraint default_io_diffCommits_info_100_ldest_cons;
    extern constraint default_io_diffCommits_info_100_pdest_cons;
    extern constraint default_io_diffCommits_info_100_rfWen_cons;
    extern constraint default_io_diffCommits_info_100_fpWen_cons;
    extern constraint default_io_diffCommits_info_100_vecWen_cons;
    extern constraint default_io_diffCommits_info_100_v0Wen_cons;
    extern constraint default_io_diffCommits_info_100_vlWen_cons;
    extern constraint default_io_diffCommits_info_101_ldest_cons;
    extern constraint default_io_diffCommits_info_101_pdest_cons;
    extern constraint default_io_diffCommits_info_101_rfWen_cons;
    extern constraint default_io_diffCommits_info_101_fpWen_cons;
    extern constraint default_io_diffCommits_info_101_vecWen_cons;
    extern constraint default_io_diffCommits_info_101_v0Wen_cons;
    extern constraint default_io_diffCommits_info_101_vlWen_cons;
    extern constraint default_io_diffCommits_info_102_ldest_cons;
    extern constraint default_io_diffCommits_info_102_pdest_cons;
    extern constraint default_io_diffCommits_info_102_rfWen_cons;
    extern constraint default_io_diffCommits_info_102_fpWen_cons;
    extern constraint default_io_diffCommits_info_102_vecWen_cons;
    extern constraint default_io_diffCommits_info_102_v0Wen_cons;
    extern constraint default_io_diffCommits_info_102_vlWen_cons;
    extern constraint default_io_diffCommits_info_103_ldest_cons;
    extern constraint default_io_diffCommits_info_103_pdest_cons;
    extern constraint default_io_diffCommits_info_103_rfWen_cons;
    extern constraint default_io_diffCommits_info_103_fpWen_cons;
    extern constraint default_io_diffCommits_info_103_vecWen_cons;
    extern constraint default_io_diffCommits_info_103_v0Wen_cons;
    extern constraint default_io_diffCommits_info_103_vlWen_cons;
    extern constraint default_io_diffCommits_info_104_ldest_cons;
    extern constraint default_io_diffCommits_info_104_pdest_cons;
    extern constraint default_io_diffCommits_info_104_rfWen_cons;
    extern constraint default_io_diffCommits_info_104_fpWen_cons;
    extern constraint default_io_diffCommits_info_104_vecWen_cons;
    extern constraint default_io_diffCommits_info_104_v0Wen_cons;
    extern constraint default_io_diffCommits_info_104_vlWen_cons;
    extern constraint default_io_diffCommits_info_105_ldest_cons;
    extern constraint default_io_diffCommits_info_105_pdest_cons;
    extern constraint default_io_diffCommits_info_105_rfWen_cons;
    extern constraint default_io_diffCommits_info_105_fpWen_cons;
    extern constraint default_io_diffCommits_info_105_vecWen_cons;
    extern constraint default_io_diffCommits_info_105_v0Wen_cons;
    extern constraint default_io_diffCommits_info_105_vlWen_cons;
    extern constraint default_io_diffCommits_info_106_ldest_cons;
    extern constraint default_io_diffCommits_info_106_pdest_cons;
    extern constraint default_io_diffCommits_info_106_rfWen_cons;
    extern constraint default_io_diffCommits_info_106_fpWen_cons;
    extern constraint default_io_diffCommits_info_106_vecWen_cons;
    extern constraint default_io_diffCommits_info_106_v0Wen_cons;
    extern constraint default_io_diffCommits_info_106_vlWen_cons;
    extern constraint default_io_diffCommits_info_107_ldest_cons;
    extern constraint default_io_diffCommits_info_107_pdest_cons;
    extern constraint default_io_diffCommits_info_107_rfWen_cons;
    extern constraint default_io_diffCommits_info_107_fpWen_cons;
    extern constraint default_io_diffCommits_info_107_vecWen_cons;
    extern constraint default_io_diffCommits_info_107_v0Wen_cons;
    extern constraint default_io_diffCommits_info_107_vlWen_cons;
    extern constraint default_io_diffCommits_info_108_ldest_cons;
    extern constraint default_io_diffCommits_info_108_pdest_cons;
    extern constraint default_io_diffCommits_info_108_rfWen_cons;
    extern constraint default_io_diffCommits_info_108_fpWen_cons;
    extern constraint default_io_diffCommits_info_108_vecWen_cons;
    extern constraint default_io_diffCommits_info_108_v0Wen_cons;
    extern constraint default_io_diffCommits_info_108_vlWen_cons;
    extern constraint default_io_diffCommits_info_109_ldest_cons;
    extern constraint default_io_diffCommits_info_109_pdest_cons;
    extern constraint default_io_diffCommits_info_109_rfWen_cons;
    extern constraint default_io_diffCommits_info_109_fpWen_cons;
    extern constraint default_io_diffCommits_info_109_vecWen_cons;
    extern constraint default_io_diffCommits_info_109_v0Wen_cons;
    extern constraint default_io_diffCommits_info_109_vlWen_cons;
    extern constraint default_io_diffCommits_info_110_ldest_cons;
    extern constraint default_io_diffCommits_info_110_pdest_cons;
    extern constraint default_io_diffCommits_info_110_rfWen_cons;
    extern constraint default_io_diffCommits_info_110_fpWen_cons;
    extern constraint default_io_diffCommits_info_110_vecWen_cons;
    extern constraint default_io_diffCommits_info_110_v0Wen_cons;
    extern constraint default_io_diffCommits_info_110_vlWen_cons;
    extern constraint default_io_diffCommits_info_111_ldest_cons;
    extern constraint default_io_diffCommits_info_111_pdest_cons;
    extern constraint default_io_diffCommits_info_111_rfWen_cons;
    extern constraint default_io_diffCommits_info_111_fpWen_cons;
    extern constraint default_io_diffCommits_info_111_vecWen_cons;
    extern constraint default_io_diffCommits_info_111_v0Wen_cons;
    extern constraint default_io_diffCommits_info_111_vlWen_cons;
    extern constraint default_io_diffCommits_info_112_ldest_cons;
    extern constraint default_io_diffCommits_info_112_pdest_cons;
    extern constraint default_io_diffCommits_info_112_rfWen_cons;
    extern constraint default_io_diffCommits_info_112_fpWen_cons;
    extern constraint default_io_diffCommits_info_112_vecWen_cons;
    extern constraint default_io_diffCommits_info_112_v0Wen_cons;
    extern constraint default_io_diffCommits_info_112_vlWen_cons;
    extern constraint default_io_diffCommits_info_113_ldest_cons;
    extern constraint default_io_diffCommits_info_113_pdest_cons;
    extern constraint default_io_diffCommits_info_113_rfWen_cons;
    extern constraint default_io_diffCommits_info_113_fpWen_cons;
    extern constraint default_io_diffCommits_info_113_vecWen_cons;
    extern constraint default_io_diffCommits_info_113_v0Wen_cons;
    extern constraint default_io_diffCommits_info_113_vlWen_cons;
    extern constraint default_io_diffCommits_info_114_ldest_cons;
    extern constraint default_io_diffCommits_info_114_pdest_cons;
    extern constraint default_io_diffCommits_info_114_rfWen_cons;
    extern constraint default_io_diffCommits_info_114_fpWen_cons;
    extern constraint default_io_diffCommits_info_114_vecWen_cons;
    extern constraint default_io_diffCommits_info_114_v0Wen_cons;
    extern constraint default_io_diffCommits_info_114_vlWen_cons;
    extern constraint default_io_diffCommits_info_115_ldest_cons;
    extern constraint default_io_diffCommits_info_115_pdest_cons;
    extern constraint default_io_diffCommits_info_115_rfWen_cons;
    extern constraint default_io_diffCommits_info_115_fpWen_cons;
    extern constraint default_io_diffCommits_info_115_vecWen_cons;
    extern constraint default_io_diffCommits_info_115_v0Wen_cons;
    extern constraint default_io_diffCommits_info_115_vlWen_cons;
    extern constraint default_io_diffCommits_info_116_ldest_cons;
    extern constraint default_io_diffCommits_info_116_pdest_cons;
    extern constraint default_io_diffCommits_info_116_rfWen_cons;
    extern constraint default_io_diffCommits_info_116_fpWen_cons;
    extern constraint default_io_diffCommits_info_116_vecWen_cons;
    extern constraint default_io_diffCommits_info_116_v0Wen_cons;
    extern constraint default_io_diffCommits_info_116_vlWen_cons;
    extern constraint default_io_diffCommits_info_117_ldest_cons;
    extern constraint default_io_diffCommits_info_117_pdest_cons;
    extern constraint default_io_diffCommits_info_117_rfWen_cons;
    extern constraint default_io_diffCommits_info_117_fpWen_cons;
    extern constraint default_io_diffCommits_info_117_vecWen_cons;
    extern constraint default_io_diffCommits_info_117_v0Wen_cons;
    extern constraint default_io_diffCommits_info_117_vlWen_cons;
    extern constraint default_io_diffCommits_info_118_ldest_cons;
    extern constraint default_io_diffCommits_info_118_pdest_cons;
    extern constraint default_io_diffCommits_info_118_rfWen_cons;
    extern constraint default_io_diffCommits_info_118_fpWen_cons;
    extern constraint default_io_diffCommits_info_118_vecWen_cons;
    extern constraint default_io_diffCommits_info_118_v0Wen_cons;
    extern constraint default_io_diffCommits_info_118_vlWen_cons;
    extern constraint default_io_diffCommits_info_119_ldest_cons;
    extern constraint default_io_diffCommits_info_119_pdest_cons;
    extern constraint default_io_diffCommits_info_119_rfWen_cons;
    extern constraint default_io_diffCommits_info_119_fpWen_cons;
    extern constraint default_io_diffCommits_info_119_vecWen_cons;
    extern constraint default_io_diffCommits_info_119_v0Wen_cons;
    extern constraint default_io_diffCommits_info_119_vlWen_cons;
    extern constraint default_io_diffCommits_info_120_ldest_cons;
    extern constraint default_io_diffCommits_info_120_pdest_cons;
    extern constraint default_io_diffCommits_info_120_rfWen_cons;
    extern constraint default_io_diffCommits_info_120_fpWen_cons;
    extern constraint default_io_diffCommits_info_120_vecWen_cons;
    extern constraint default_io_diffCommits_info_120_v0Wen_cons;
    extern constraint default_io_diffCommits_info_120_vlWen_cons;
    extern constraint default_io_diffCommits_info_121_ldest_cons;
    extern constraint default_io_diffCommits_info_121_pdest_cons;
    extern constraint default_io_diffCommits_info_121_rfWen_cons;
    extern constraint default_io_diffCommits_info_121_fpWen_cons;
    extern constraint default_io_diffCommits_info_121_vecWen_cons;
    extern constraint default_io_diffCommits_info_121_v0Wen_cons;
    extern constraint default_io_diffCommits_info_121_vlWen_cons;
    extern constraint default_io_diffCommits_info_122_ldest_cons;
    extern constraint default_io_diffCommits_info_122_pdest_cons;
    extern constraint default_io_diffCommits_info_122_rfWen_cons;
    extern constraint default_io_diffCommits_info_122_fpWen_cons;
    extern constraint default_io_diffCommits_info_122_vecWen_cons;
    extern constraint default_io_diffCommits_info_122_v0Wen_cons;
    extern constraint default_io_diffCommits_info_122_vlWen_cons;
    extern constraint default_io_diffCommits_info_123_ldest_cons;
    extern constraint default_io_diffCommits_info_123_pdest_cons;
    extern constraint default_io_diffCommits_info_123_rfWen_cons;
    extern constraint default_io_diffCommits_info_123_fpWen_cons;
    extern constraint default_io_diffCommits_info_123_vecWen_cons;
    extern constraint default_io_diffCommits_info_123_v0Wen_cons;
    extern constraint default_io_diffCommits_info_123_vlWen_cons;
    extern constraint default_io_diffCommits_info_124_ldest_cons;
    extern constraint default_io_diffCommits_info_124_pdest_cons;
    extern constraint default_io_diffCommits_info_124_rfWen_cons;
    extern constraint default_io_diffCommits_info_124_fpWen_cons;
    extern constraint default_io_diffCommits_info_124_vecWen_cons;
    extern constraint default_io_diffCommits_info_124_v0Wen_cons;
    extern constraint default_io_diffCommits_info_124_vlWen_cons;
    extern constraint default_io_diffCommits_info_125_ldest_cons;
    extern constraint default_io_diffCommits_info_125_pdest_cons;
    extern constraint default_io_diffCommits_info_125_rfWen_cons;
    extern constraint default_io_diffCommits_info_125_fpWen_cons;
    extern constraint default_io_diffCommits_info_125_vecWen_cons;
    extern constraint default_io_diffCommits_info_125_v0Wen_cons;
    extern constraint default_io_diffCommits_info_125_vlWen_cons;
    extern constraint default_io_diffCommits_info_126_ldest_cons;
    extern constraint default_io_diffCommits_info_126_pdest_cons;
    extern constraint default_io_diffCommits_info_126_rfWen_cons;
    extern constraint default_io_diffCommits_info_126_fpWen_cons;
    extern constraint default_io_diffCommits_info_126_vecWen_cons;
    extern constraint default_io_diffCommits_info_126_v0Wen_cons;
    extern constraint default_io_diffCommits_info_126_vlWen_cons;
    extern constraint default_io_diffCommits_info_127_ldest_cons;
    extern constraint default_io_diffCommits_info_127_pdest_cons;
    extern constraint default_io_diffCommits_info_127_rfWen_cons;
    extern constraint default_io_diffCommits_info_127_fpWen_cons;
    extern constraint default_io_diffCommits_info_127_vecWen_cons;
    extern constraint default_io_diffCommits_info_127_v0Wen_cons;
    extern constraint default_io_diffCommits_info_127_vlWen_cons;
    extern constraint default_io_diffCommits_info_128_ldest_cons;
    extern constraint default_io_diffCommits_info_128_pdest_cons;
    extern constraint default_io_diffCommits_info_128_rfWen_cons;
    extern constraint default_io_diffCommits_info_128_fpWen_cons;
    extern constraint default_io_diffCommits_info_128_vecWen_cons;
    extern constraint default_io_diffCommits_info_128_v0Wen_cons;
    extern constraint default_io_diffCommits_info_128_vlWen_cons;
    extern constraint default_io_diffCommits_info_129_ldest_cons;
    extern constraint default_io_diffCommits_info_129_pdest_cons;
    extern constraint default_io_diffCommits_info_129_rfWen_cons;
    extern constraint default_io_diffCommits_info_129_fpWen_cons;
    extern constraint default_io_diffCommits_info_129_vecWen_cons;
    extern constraint default_io_diffCommits_info_129_v0Wen_cons;
    extern constraint default_io_diffCommits_info_129_vlWen_cons;
    extern constraint default_io_diffCommits_info_130_ldest_cons;
    extern constraint default_io_diffCommits_info_130_pdest_cons;
    extern constraint default_io_diffCommits_info_130_rfWen_cons;
    extern constraint default_io_diffCommits_info_130_fpWen_cons;
    extern constraint default_io_diffCommits_info_130_vecWen_cons;
    extern constraint default_io_diffCommits_info_130_v0Wen_cons;
    extern constraint default_io_diffCommits_info_130_vlWen_cons;
    extern constraint default_io_diffCommits_info_131_ldest_cons;
    extern constraint default_io_diffCommits_info_131_pdest_cons;
    extern constraint default_io_diffCommits_info_131_rfWen_cons;
    extern constraint default_io_diffCommits_info_131_fpWen_cons;
    extern constraint default_io_diffCommits_info_131_vecWen_cons;
    extern constraint default_io_diffCommits_info_131_v0Wen_cons;
    extern constraint default_io_diffCommits_info_131_vlWen_cons;
    extern constraint default_io_diffCommits_info_132_ldest_cons;
    extern constraint default_io_diffCommits_info_132_pdest_cons;
    extern constraint default_io_diffCommits_info_132_rfWen_cons;
    extern constraint default_io_diffCommits_info_132_fpWen_cons;
    extern constraint default_io_diffCommits_info_132_vecWen_cons;
    extern constraint default_io_diffCommits_info_132_v0Wen_cons;
    extern constraint default_io_diffCommits_info_132_vlWen_cons;
    extern constraint default_io_diffCommits_info_133_ldest_cons;
    extern constraint default_io_diffCommits_info_133_pdest_cons;
    extern constraint default_io_diffCommits_info_133_rfWen_cons;
    extern constraint default_io_diffCommits_info_133_fpWen_cons;
    extern constraint default_io_diffCommits_info_133_vecWen_cons;
    extern constraint default_io_diffCommits_info_133_v0Wen_cons;
    extern constraint default_io_diffCommits_info_133_vlWen_cons;
    extern constraint default_io_diffCommits_info_134_ldest_cons;
    extern constraint default_io_diffCommits_info_134_pdest_cons;
    extern constraint default_io_diffCommits_info_134_rfWen_cons;
    extern constraint default_io_diffCommits_info_134_fpWen_cons;
    extern constraint default_io_diffCommits_info_134_vecWen_cons;
    extern constraint default_io_diffCommits_info_134_v0Wen_cons;
    extern constraint default_io_diffCommits_info_134_vlWen_cons;
    extern constraint default_io_diffCommits_info_135_ldest_cons;
    extern constraint default_io_diffCommits_info_135_pdest_cons;
    extern constraint default_io_diffCommits_info_135_rfWen_cons;
    extern constraint default_io_diffCommits_info_135_fpWen_cons;
    extern constraint default_io_diffCommits_info_135_vecWen_cons;
    extern constraint default_io_diffCommits_info_135_v0Wen_cons;
    extern constraint default_io_diffCommits_info_135_vlWen_cons;
    extern constraint default_io_diffCommits_info_136_ldest_cons;
    extern constraint default_io_diffCommits_info_136_pdest_cons;
    extern constraint default_io_diffCommits_info_136_rfWen_cons;
    extern constraint default_io_diffCommits_info_136_fpWen_cons;
    extern constraint default_io_diffCommits_info_136_vecWen_cons;
    extern constraint default_io_diffCommits_info_136_v0Wen_cons;
    extern constraint default_io_diffCommits_info_136_vlWen_cons;
    extern constraint default_io_diffCommits_info_137_ldest_cons;
    extern constraint default_io_diffCommits_info_137_pdest_cons;
    extern constraint default_io_diffCommits_info_137_rfWen_cons;
    extern constraint default_io_diffCommits_info_137_fpWen_cons;
    extern constraint default_io_diffCommits_info_137_vecWen_cons;
    extern constraint default_io_diffCommits_info_137_v0Wen_cons;
    extern constraint default_io_diffCommits_info_137_vlWen_cons;
    extern constraint default_io_diffCommits_info_138_ldest_cons;
    extern constraint default_io_diffCommits_info_138_pdest_cons;
    extern constraint default_io_diffCommits_info_138_rfWen_cons;
    extern constraint default_io_diffCommits_info_138_fpWen_cons;
    extern constraint default_io_diffCommits_info_138_vecWen_cons;
    extern constraint default_io_diffCommits_info_138_v0Wen_cons;
    extern constraint default_io_diffCommits_info_138_vlWen_cons;
    extern constraint default_io_diffCommits_info_139_ldest_cons;
    extern constraint default_io_diffCommits_info_139_pdest_cons;
    extern constraint default_io_diffCommits_info_139_rfWen_cons;
    extern constraint default_io_diffCommits_info_139_fpWen_cons;
    extern constraint default_io_diffCommits_info_139_vecWen_cons;
    extern constraint default_io_diffCommits_info_139_v0Wen_cons;
    extern constraint default_io_diffCommits_info_139_vlWen_cons;
    extern constraint default_io_diffCommits_info_140_ldest_cons;
    extern constraint default_io_diffCommits_info_140_pdest_cons;
    extern constraint default_io_diffCommits_info_140_rfWen_cons;
    extern constraint default_io_diffCommits_info_140_fpWen_cons;
    extern constraint default_io_diffCommits_info_140_vecWen_cons;
    extern constraint default_io_diffCommits_info_140_v0Wen_cons;
    extern constraint default_io_diffCommits_info_140_vlWen_cons;
    extern constraint default_io_diffCommits_info_141_ldest_cons;
    extern constraint default_io_diffCommits_info_141_pdest_cons;
    extern constraint default_io_diffCommits_info_141_rfWen_cons;
    extern constraint default_io_diffCommits_info_141_fpWen_cons;
    extern constraint default_io_diffCommits_info_141_vecWen_cons;
    extern constraint default_io_diffCommits_info_141_v0Wen_cons;
    extern constraint default_io_diffCommits_info_141_vlWen_cons;
    extern constraint default_io_diffCommits_info_142_ldest_cons;
    extern constraint default_io_diffCommits_info_142_pdest_cons;
    extern constraint default_io_diffCommits_info_142_rfWen_cons;
    extern constraint default_io_diffCommits_info_142_fpWen_cons;
    extern constraint default_io_diffCommits_info_142_vecWen_cons;
    extern constraint default_io_diffCommits_info_142_v0Wen_cons;
    extern constraint default_io_diffCommits_info_142_vlWen_cons;
    extern constraint default_io_diffCommits_info_143_ldest_cons;
    extern constraint default_io_diffCommits_info_143_pdest_cons;
    extern constraint default_io_diffCommits_info_143_rfWen_cons;
    extern constraint default_io_diffCommits_info_143_fpWen_cons;
    extern constraint default_io_diffCommits_info_143_vecWen_cons;
    extern constraint default_io_diffCommits_info_143_v0Wen_cons;
    extern constraint default_io_diffCommits_info_143_vlWen_cons;
    extern constraint default_io_diffCommits_info_144_ldest_cons;
    extern constraint default_io_diffCommits_info_144_pdest_cons;
    extern constraint default_io_diffCommits_info_144_rfWen_cons;
    extern constraint default_io_diffCommits_info_144_fpWen_cons;
    extern constraint default_io_diffCommits_info_144_vecWen_cons;
    extern constraint default_io_diffCommits_info_144_v0Wen_cons;
    extern constraint default_io_diffCommits_info_144_vlWen_cons;
    extern constraint default_io_diffCommits_info_145_ldest_cons;
    extern constraint default_io_diffCommits_info_145_pdest_cons;
    extern constraint default_io_diffCommits_info_145_rfWen_cons;
    extern constraint default_io_diffCommits_info_145_fpWen_cons;
    extern constraint default_io_diffCommits_info_145_vecWen_cons;
    extern constraint default_io_diffCommits_info_145_v0Wen_cons;
    extern constraint default_io_diffCommits_info_145_vlWen_cons;
    extern constraint default_io_diffCommits_info_146_ldest_cons;
    extern constraint default_io_diffCommits_info_146_pdest_cons;
    extern constraint default_io_diffCommits_info_146_rfWen_cons;
    extern constraint default_io_diffCommits_info_146_fpWen_cons;
    extern constraint default_io_diffCommits_info_146_vecWen_cons;
    extern constraint default_io_diffCommits_info_146_v0Wen_cons;
    extern constraint default_io_diffCommits_info_146_vlWen_cons;
    extern constraint default_io_diffCommits_info_147_ldest_cons;
    extern constraint default_io_diffCommits_info_147_pdest_cons;
    extern constraint default_io_diffCommits_info_147_rfWen_cons;
    extern constraint default_io_diffCommits_info_147_fpWen_cons;
    extern constraint default_io_diffCommits_info_147_vecWen_cons;
    extern constraint default_io_diffCommits_info_147_v0Wen_cons;
    extern constraint default_io_diffCommits_info_147_vlWen_cons;
    extern constraint default_io_diffCommits_info_148_ldest_cons;
    extern constraint default_io_diffCommits_info_148_pdest_cons;
    extern constraint default_io_diffCommits_info_148_rfWen_cons;
    extern constraint default_io_diffCommits_info_148_fpWen_cons;
    extern constraint default_io_diffCommits_info_148_vecWen_cons;
    extern constraint default_io_diffCommits_info_148_v0Wen_cons;
    extern constraint default_io_diffCommits_info_148_vlWen_cons;
    extern constraint default_io_diffCommits_info_149_ldest_cons;
    extern constraint default_io_diffCommits_info_149_pdest_cons;
    extern constraint default_io_diffCommits_info_149_rfWen_cons;
    extern constraint default_io_diffCommits_info_149_fpWen_cons;
    extern constraint default_io_diffCommits_info_149_vecWen_cons;
    extern constraint default_io_diffCommits_info_149_v0Wen_cons;
    extern constraint default_io_diffCommits_info_149_vlWen_cons;
    extern constraint default_io_diffCommits_info_150_ldest_cons;
    extern constraint default_io_diffCommits_info_150_pdest_cons;
    extern constraint default_io_diffCommits_info_150_rfWen_cons;
    extern constraint default_io_diffCommits_info_150_fpWen_cons;
    extern constraint default_io_diffCommits_info_150_vecWen_cons;
    extern constraint default_io_diffCommits_info_150_v0Wen_cons;
    extern constraint default_io_diffCommits_info_150_vlWen_cons;
    extern constraint default_io_diffCommits_info_151_ldest_cons;
    extern constraint default_io_diffCommits_info_151_pdest_cons;
    extern constraint default_io_diffCommits_info_151_rfWen_cons;
    extern constraint default_io_diffCommits_info_151_fpWen_cons;
    extern constraint default_io_diffCommits_info_151_vecWen_cons;
    extern constraint default_io_diffCommits_info_151_v0Wen_cons;
    extern constraint default_io_diffCommits_info_151_vlWen_cons;
    extern constraint default_io_diffCommits_info_152_ldest_cons;
    extern constraint default_io_diffCommits_info_152_pdest_cons;
    extern constraint default_io_diffCommits_info_152_rfWen_cons;
    extern constraint default_io_diffCommits_info_152_fpWen_cons;
    extern constraint default_io_diffCommits_info_152_vecWen_cons;
    extern constraint default_io_diffCommits_info_152_v0Wen_cons;
    extern constraint default_io_diffCommits_info_152_vlWen_cons;
    extern constraint default_io_diffCommits_info_153_ldest_cons;
    extern constraint default_io_diffCommits_info_153_pdest_cons;
    extern constraint default_io_diffCommits_info_153_rfWen_cons;
    extern constraint default_io_diffCommits_info_153_fpWen_cons;
    extern constraint default_io_diffCommits_info_153_vecWen_cons;
    extern constraint default_io_diffCommits_info_153_v0Wen_cons;
    extern constraint default_io_diffCommits_info_153_vlWen_cons;
    extern constraint default_io_diffCommits_info_154_ldest_cons;
    extern constraint default_io_diffCommits_info_154_pdest_cons;
    extern constraint default_io_diffCommits_info_154_rfWen_cons;
    extern constraint default_io_diffCommits_info_154_fpWen_cons;
    extern constraint default_io_diffCommits_info_154_vecWen_cons;
    extern constraint default_io_diffCommits_info_154_v0Wen_cons;
    extern constraint default_io_diffCommits_info_154_vlWen_cons;
    extern constraint default_io_diffCommits_info_155_ldest_cons;
    extern constraint default_io_diffCommits_info_155_pdest_cons;
    extern constraint default_io_diffCommits_info_155_rfWen_cons;
    extern constraint default_io_diffCommits_info_155_fpWen_cons;
    extern constraint default_io_diffCommits_info_155_vecWen_cons;
    extern constraint default_io_diffCommits_info_155_v0Wen_cons;
    extern constraint default_io_diffCommits_info_155_vlWen_cons;
    extern constraint default_io_diffCommits_info_156_ldest_cons;
    extern constraint default_io_diffCommits_info_156_pdest_cons;
    extern constraint default_io_diffCommits_info_156_rfWen_cons;
    extern constraint default_io_diffCommits_info_156_fpWen_cons;
    extern constraint default_io_diffCommits_info_156_vecWen_cons;
    extern constraint default_io_diffCommits_info_156_v0Wen_cons;
    extern constraint default_io_diffCommits_info_156_vlWen_cons;
    extern constraint default_io_diffCommits_info_157_ldest_cons;
    extern constraint default_io_diffCommits_info_157_pdest_cons;
    extern constraint default_io_diffCommits_info_157_rfWen_cons;
    extern constraint default_io_diffCommits_info_157_fpWen_cons;
    extern constraint default_io_diffCommits_info_157_vecWen_cons;
    extern constraint default_io_diffCommits_info_157_v0Wen_cons;
    extern constraint default_io_diffCommits_info_157_vlWen_cons;
    extern constraint default_io_diffCommits_info_158_ldest_cons;
    extern constraint default_io_diffCommits_info_158_pdest_cons;
    extern constraint default_io_diffCommits_info_158_rfWen_cons;
    extern constraint default_io_diffCommits_info_158_fpWen_cons;
    extern constraint default_io_diffCommits_info_158_vecWen_cons;
    extern constraint default_io_diffCommits_info_158_v0Wen_cons;
    extern constraint default_io_diffCommits_info_158_vlWen_cons;
    extern constraint default_io_diffCommits_info_159_ldest_cons;
    extern constraint default_io_diffCommits_info_159_pdest_cons;
    extern constraint default_io_diffCommits_info_159_rfWen_cons;
    extern constraint default_io_diffCommits_info_159_fpWen_cons;
    extern constraint default_io_diffCommits_info_159_vecWen_cons;
    extern constraint default_io_diffCommits_info_159_v0Wen_cons;
    extern constraint default_io_diffCommits_info_159_vlWen_cons;
    extern constraint default_io_diffCommits_info_160_ldest_cons;
    extern constraint default_io_diffCommits_info_160_pdest_cons;
    extern constraint default_io_diffCommits_info_160_rfWen_cons;
    extern constraint default_io_diffCommits_info_160_fpWen_cons;
    extern constraint default_io_diffCommits_info_160_vecWen_cons;
    extern constraint default_io_diffCommits_info_160_v0Wen_cons;
    extern constraint default_io_diffCommits_info_160_vlWen_cons;
    extern constraint default_io_diffCommits_info_161_ldest_cons;
    extern constraint default_io_diffCommits_info_161_pdest_cons;
    extern constraint default_io_diffCommits_info_161_rfWen_cons;
    extern constraint default_io_diffCommits_info_161_fpWen_cons;
    extern constraint default_io_diffCommits_info_161_vecWen_cons;
    extern constraint default_io_diffCommits_info_161_v0Wen_cons;
    extern constraint default_io_diffCommits_info_161_vlWen_cons;
    extern constraint default_io_diffCommits_info_162_ldest_cons;
    extern constraint default_io_diffCommits_info_162_pdest_cons;
    extern constraint default_io_diffCommits_info_162_rfWen_cons;
    extern constraint default_io_diffCommits_info_162_fpWen_cons;
    extern constraint default_io_diffCommits_info_162_vecWen_cons;
    extern constraint default_io_diffCommits_info_162_v0Wen_cons;
    extern constraint default_io_diffCommits_info_162_vlWen_cons;
    extern constraint default_io_diffCommits_info_163_ldest_cons;
    extern constraint default_io_diffCommits_info_163_pdest_cons;
    extern constraint default_io_diffCommits_info_163_rfWen_cons;
    extern constraint default_io_diffCommits_info_163_fpWen_cons;
    extern constraint default_io_diffCommits_info_163_vecWen_cons;
    extern constraint default_io_diffCommits_info_163_v0Wen_cons;
    extern constraint default_io_diffCommits_info_163_vlWen_cons;
    extern constraint default_io_diffCommits_info_164_ldest_cons;
    extern constraint default_io_diffCommits_info_164_pdest_cons;
    extern constraint default_io_diffCommits_info_164_rfWen_cons;
    extern constraint default_io_diffCommits_info_164_fpWen_cons;
    extern constraint default_io_diffCommits_info_164_vecWen_cons;
    extern constraint default_io_diffCommits_info_164_v0Wen_cons;
    extern constraint default_io_diffCommits_info_164_vlWen_cons;
    extern constraint default_io_diffCommits_info_165_ldest_cons;
    extern constraint default_io_diffCommits_info_165_pdest_cons;
    extern constraint default_io_diffCommits_info_165_rfWen_cons;
    extern constraint default_io_diffCommits_info_165_fpWen_cons;
    extern constraint default_io_diffCommits_info_165_vecWen_cons;
    extern constraint default_io_diffCommits_info_165_v0Wen_cons;
    extern constraint default_io_diffCommits_info_165_vlWen_cons;
    extern constraint default_io_diffCommits_info_166_ldest_cons;
    extern constraint default_io_diffCommits_info_166_pdest_cons;
    extern constraint default_io_diffCommits_info_166_rfWen_cons;
    extern constraint default_io_diffCommits_info_166_fpWen_cons;
    extern constraint default_io_diffCommits_info_166_vecWen_cons;
    extern constraint default_io_diffCommits_info_166_v0Wen_cons;
    extern constraint default_io_diffCommits_info_166_vlWen_cons;
    extern constraint default_io_diffCommits_info_167_ldest_cons;
    extern constraint default_io_diffCommits_info_167_pdest_cons;
    extern constraint default_io_diffCommits_info_167_rfWen_cons;
    extern constraint default_io_diffCommits_info_167_fpWen_cons;
    extern constraint default_io_diffCommits_info_167_vecWen_cons;
    extern constraint default_io_diffCommits_info_167_v0Wen_cons;
    extern constraint default_io_diffCommits_info_167_vlWen_cons;
    extern constraint default_io_diffCommits_info_168_ldest_cons;
    extern constraint default_io_diffCommits_info_168_pdest_cons;
    extern constraint default_io_diffCommits_info_168_rfWen_cons;
    extern constraint default_io_diffCommits_info_168_fpWen_cons;
    extern constraint default_io_diffCommits_info_168_vecWen_cons;
    extern constraint default_io_diffCommits_info_168_v0Wen_cons;
    extern constraint default_io_diffCommits_info_168_vlWen_cons;
    extern constraint default_io_diffCommits_info_169_ldest_cons;
    extern constraint default_io_diffCommits_info_169_pdest_cons;
    extern constraint default_io_diffCommits_info_169_rfWen_cons;
    extern constraint default_io_diffCommits_info_169_fpWen_cons;
    extern constraint default_io_diffCommits_info_169_vecWen_cons;
    extern constraint default_io_diffCommits_info_169_v0Wen_cons;
    extern constraint default_io_diffCommits_info_169_vlWen_cons;
    extern constraint default_io_diffCommits_info_170_ldest_cons;
    extern constraint default_io_diffCommits_info_170_pdest_cons;
    extern constraint default_io_diffCommits_info_170_rfWen_cons;
    extern constraint default_io_diffCommits_info_170_fpWen_cons;
    extern constraint default_io_diffCommits_info_170_vecWen_cons;
    extern constraint default_io_diffCommits_info_170_v0Wen_cons;
    extern constraint default_io_diffCommits_info_170_vlWen_cons;
    extern constraint default_io_diffCommits_info_171_ldest_cons;
    extern constraint default_io_diffCommits_info_171_pdest_cons;
    extern constraint default_io_diffCommits_info_171_rfWen_cons;
    extern constraint default_io_diffCommits_info_171_fpWen_cons;
    extern constraint default_io_diffCommits_info_171_vecWen_cons;
    extern constraint default_io_diffCommits_info_171_v0Wen_cons;
    extern constraint default_io_diffCommits_info_171_vlWen_cons;
    extern constraint default_io_diffCommits_info_172_ldest_cons;
    extern constraint default_io_diffCommits_info_172_pdest_cons;
    extern constraint default_io_diffCommits_info_172_rfWen_cons;
    extern constraint default_io_diffCommits_info_172_fpWen_cons;
    extern constraint default_io_diffCommits_info_172_vecWen_cons;
    extern constraint default_io_diffCommits_info_172_v0Wen_cons;
    extern constraint default_io_diffCommits_info_172_vlWen_cons;
    extern constraint default_io_diffCommits_info_173_ldest_cons;
    extern constraint default_io_diffCommits_info_173_pdest_cons;
    extern constraint default_io_diffCommits_info_173_rfWen_cons;
    extern constraint default_io_diffCommits_info_173_fpWen_cons;
    extern constraint default_io_diffCommits_info_173_vecWen_cons;
    extern constraint default_io_diffCommits_info_173_v0Wen_cons;
    extern constraint default_io_diffCommits_info_173_vlWen_cons;
    extern constraint default_io_diffCommits_info_174_ldest_cons;
    extern constraint default_io_diffCommits_info_174_pdest_cons;
    extern constraint default_io_diffCommits_info_174_rfWen_cons;
    extern constraint default_io_diffCommits_info_174_fpWen_cons;
    extern constraint default_io_diffCommits_info_174_vecWen_cons;
    extern constraint default_io_diffCommits_info_174_v0Wen_cons;
    extern constraint default_io_diffCommits_info_174_vlWen_cons;
    extern constraint default_io_diffCommits_info_175_ldest_cons;
    extern constraint default_io_diffCommits_info_175_pdest_cons;
    extern constraint default_io_diffCommits_info_175_rfWen_cons;
    extern constraint default_io_diffCommits_info_175_fpWen_cons;
    extern constraint default_io_diffCommits_info_175_vecWen_cons;
    extern constraint default_io_diffCommits_info_175_v0Wen_cons;
    extern constraint default_io_diffCommits_info_175_vlWen_cons;
    extern constraint default_io_diffCommits_info_176_ldest_cons;
    extern constraint default_io_diffCommits_info_176_pdest_cons;
    extern constraint default_io_diffCommits_info_176_rfWen_cons;
    extern constraint default_io_diffCommits_info_176_fpWen_cons;
    extern constraint default_io_diffCommits_info_176_vecWen_cons;
    extern constraint default_io_diffCommits_info_176_v0Wen_cons;
    extern constraint default_io_diffCommits_info_176_vlWen_cons;
    extern constraint default_io_diffCommits_info_177_ldest_cons;
    extern constraint default_io_diffCommits_info_177_pdest_cons;
    extern constraint default_io_diffCommits_info_177_rfWen_cons;
    extern constraint default_io_diffCommits_info_177_fpWen_cons;
    extern constraint default_io_diffCommits_info_177_vecWen_cons;
    extern constraint default_io_diffCommits_info_177_v0Wen_cons;
    extern constraint default_io_diffCommits_info_177_vlWen_cons;
    extern constraint default_io_diffCommits_info_178_ldest_cons;
    extern constraint default_io_diffCommits_info_178_pdest_cons;
    extern constraint default_io_diffCommits_info_178_rfWen_cons;
    extern constraint default_io_diffCommits_info_178_fpWen_cons;
    extern constraint default_io_diffCommits_info_178_vecWen_cons;
    extern constraint default_io_diffCommits_info_178_v0Wen_cons;
    extern constraint default_io_diffCommits_info_178_vlWen_cons;
    extern constraint default_io_diffCommits_info_179_ldest_cons;
    extern constraint default_io_diffCommits_info_179_pdest_cons;
    extern constraint default_io_diffCommits_info_179_rfWen_cons;
    extern constraint default_io_diffCommits_info_179_fpWen_cons;
    extern constraint default_io_diffCommits_info_179_vecWen_cons;
    extern constraint default_io_diffCommits_info_179_v0Wen_cons;
    extern constraint default_io_diffCommits_info_179_vlWen_cons;
    extern constraint default_io_diffCommits_info_180_ldest_cons;
    extern constraint default_io_diffCommits_info_180_pdest_cons;
    extern constraint default_io_diffCommits_info_180_rfWen_cons;
    extern constraint default_io_diffCommits_info_180_fpWen_cons;
    extern constraint default_io_diffCommits_info_180_vecWen_cons;
    extern constraint default_io_diffCommits_info_180_v0Wen_cons;
    extern constraint default_io_diffCommits_info_180_vlWen_cons;
    extern constraint default_io_diffCommits_info_181_ldest_cons;
    extern constraint default_io_diffCommits_info_181_pdest_cons;
    extern constraint default_io_diffCommits_info_181_rfWen_cons;
    extern constraint default_io_diffCommits_info_181_fpWen_cons;
    extern constraint default_io_diffCommits_info_181_vecWen_cons;
    extern constraint default_io_diffCommits_info_181_v0Wen_cons;
    extern constraint default_io_diffCommits_info_181_vlWen_cons;
    extern constraint default_io_diffCommits_info_182_ldest_cons;
    extern constraint default_io_diffCommits_info_182_pdest_cons;
    extern constraint default_io_diffCommits_info_182_rfWen_cons;
    extern constraint default_io_diffCommits_info_182_fpWen_cons;
    extern constraint default_io_diffCommits_info_182_vecWen_cons;
    extern constraint default_io_diffCommits_info_182_v0Wen_cons;
    extern constraint default_io_diffCommits_info_182_vlWen_cons;
    extern constraint default_io_diffCommits_info_183_ldest_cons;
    extern constraint default_io_diffCommits_info_183_pdest_cons;
    extern constraint default_io_diffCommits_info_183_rfWen_cons;
    extern constraint default_io_diffCommits_info_183_fpWen_cons;
    extern constraint default_io_diffCommits_info_183_vecWen_cons;
    extern constraint default_io_diffCommits_info_183_v0Wen_cons;
    extern constraint default_io_diffCommits_info_183_vlWen_cons;
    extern constraint default_io_diffCommits_info_184_ldest_cons;
    extern constraint default_io_diffCommits_info_184_pdest_cons;
    extern constraint default_io_diffCommits_info_184_rfWen_cons;
    extern constraint default_io_diffCommits_info_184_fpWen_cons;
    extern constraint default_io_diffCommits_info_184_vecWen_cons;
    extern constraint default_io_diffCommits_info_184_v0Wen_cons;
    extern constraint default_io_diffCommits_info_184_vlWen_cons;
    extern constraint default_io_diffCommits_info_185_ldest_cons;
    extern constraint default_io_diffCommits_info_185_pdest_cons;
    extern constraint default_io_diffCommits_info_185_rfWen_cons;
    extern constraint default_io_diffCommits_info_185_fpWen_cons;
    extern constraint default_io_diffCommits_info_185_vecWen_cons;
    extern constraint default_io_diffCommits_info_185_v0Wen_cons;
    extern constraint default_io_diffCommits_info_185_vlWen_cons;
    extern constraint default_io_diffCommits_info_186_ldest_cons;
    extern constraint default_io_diffCommits_info_186_pdest_cons;
    extern constraint default_io_diffCommits_info_186_rfWen_cons;
    extern constraint default_io_diffCommits_info_186_fpWen_cons;
    extern constraint default_io_diffCommits_info_186_vecWen_cons;
    extern constraint default_io_diffCommits_info_186_v0Wen_cons;
    extern constraint default_io_diffCommits_info_186_vlWen_cons;
    extern constraint default_io_diffCommits_info_187_ldest_cons;
    extern constraint default_io_diffCommits_info_187_pdest_cons;
    extern constraint default_io_diffCommits_info_187_rfWen_cons;
    extern constraint default_io_diffCommits_info_187_fpWen_cons;
    extern constraint default_io_diffCommits_info_187_vecWen_cons;
    extern constraint default_io_diffCommits_info_187_v0Wen_cons;
    extern constraint default_io_diffCommits_info_187_vlWen_cons;
    extern constraint default_io_diffCommits_info_188_ldest_cons;
    extern constraint default_io_diffCommits_info_188_pdest_cons;
    extern constraint default_io_diffCommits_info_188_rfWen_cons;
    extern constraint default_io_diffCommits_info_188_fpWen_cons;
    extern constraint default_io_diffCommits_info_188_vecWen_cons;
    extern constraint default_io_diffCommits_info_188_v0Wen_cons;
    extern constraint default_io_diffCommits_info_188_vlWen_cons;
    extern constraint default_io_diffCommits_info_189_ldest_cons;
    extern constraint default_io_diffCommits_info_189_pdest_cons;
    extern constraint default_io_diffCommits_info_189_rfWen_cons;
    extern constraint default_io_diffCommits_info_189_fpWen_cons;
    extern constraint default_io_diffCommits_info_189_vecWen_cons;
    extern constraint default_io_diffCommits_info_189_v0Wen_cons;
    extern constraint default_io_diffCommits_info_189_vlWen_cons;
    extern constraint default_io_diffCommits_info_190_ldest_cons;
    extern constraint default_io_diffCommits_info_190_pdest_cons;
    extern constraint default_io_diffCommits_info_190_rfWen_cons;
    extern constraint default_io_diffCommits_info_190_fpWen_cons;
    extern constraint default_io_diffCommits_info_190_vecWen_cons;
    extern constraint default_io_diffCommits_info_190_v0Wen_cons;
    extern constraint default_io_diffCommits_info_190_vlWen_cons;
    extern constraint default_io_diffCommits_info_191_ldest_cons;
    extern constraint default_io_diffCommits_info_191_pdest_cons;
    extern constraint default_io_diffCommits_info_191_rfWen_cons;
    extern constraint default_io_diffCommits_info_191_fpWen_cons;
    extern constraint default_io_diffCommits_info_191_vecWen_cons;
    extern constraint default_io_diffCommits_info_191_v0Wen_cons;
    extern constraint default_io_diffCommits_info_191_vlWen_cons;
    extern constraint default_io_diffCommits_info_192_ldest_cons;
    extern constraint default_io_diffCommits_info_192_pdest_cons;
    extern constraint default_io_diffCommits_info_192_rfWen_cons;
    extern constraint default_io_diffCommits_info_192_fpWen_cons;
    extern constraint default_io_diffCommits_info_192_vecWen_cons;
    extern constraint default_io_diffCommits_info_192_v0Wen_cons;
    extern constraint default_io_diffCommits_info_192_vlWen_cons;
    extern constraint default_io_diffCommits_info_193_ldest_cons;
    extern constraint default_io_diffCommits_info_193_pdest_cons;
    extern constraint default_io_diffCommits_info_193_rfWen_cons;
    extern constraint default_io_diffCommits_info_193_fpWen_cons;
    extern constraint default_io_diffCommits_info_193_vecWen_cons;
    extern constraint default_io_diffCommits_info_193_v0Wen_cons;
    extern constraint default_io_diffCommits_info_193_vlWen_cons;
    extern constraint default_io_diffCommits_info_194_ldest_cons;
    extern constraint default_io_diffCommits_info_194_pdest_cons;
    extern constraint default_io_diffCommits_info_194_rfWen_cons;
    extern constraint default_io_diffCommits_info_194_fpWen_cons;
    extern constraint default_io_diffCommits_info_194_vecWen_cons;
    extern constraint default_io_diffCommits_info_194_v0Wen_cons;
    extern constraint default_io_diffCommits_info_194_vlWen_cons;
    extern constraint default_io_diffCommits_info_195_ldest_cons;
    extern constraint default_io_diffCommits_info_195_pdest_cons;
    extern constraint default_io_diffCommits_info_195_rfWen_cons;
    extern constraint default_io_diffCommits_info_195_fpWen_cons;
    extern constraint default_io_diffCommits_info_195_vecWen_cons;
    extern constraint default_io_diffCommits_info_195_v0Wen_cons;
    extern constraint default_io_diffCommits_info_195_vlWen_cons;
    extern constraint default_io_diffCommits_info_196_ldest_cons;
    extern constraint default_io_diffCommits_info_196_pdest_cons;
    extern constraint default_io_diffCommits_info_196_rfWen_cons;
    extern constraint default_io_diffCommits_info_196_fpWen_cons;
    extern constraint default_io_diffCommits_info_196_vecWen_cons;
    extern constraint default_io_diffCommits_info_196_v0Wen_cons;
    extern constraint default_io_diffCommits_info_196_vlWen_cons;
    extern constraint default_io_diffCommits_info_197_ldest_cons;
    extern constraint default_io_diffCommits_info_197_pdest_cons;
    extern constraint default_io_diffCommits_info_197_rfWen_cons;
    extern constraint default_io_diffCommits_info_197_fpWen_cons;
    extern constraint default_io_diffCommits_info_197_vecWen_cons;
    extern constraint default_io_diffCommits_info_197_v0Wen_cons;
    extern constraint default_io_diffCommits_info_197_vlWen_cons;
    extern constraint default_io_diffCommits_info_198_ldest_cons;
    extern constraint default_io_diffCommits_info_198_pdest_cons;
    extern constraint default_io_diffCommits_info_198_rfWen_cons;
    extern constraint default_io_diffCommits_info_198_fpWen_cons;
    extern constraint default_io_diffCommits_info_198_vecWen_cons;
    extern constraint default_io_diffCommits_info_198_v0Wen_cons;
    extern constraint default_io_diffCommits_info_198_vlWen_cons;
    extern constraint default_io_diffCommits_info_199_ldest_cons;
    extern constraint default_io_diffCommits_info_199_pdest_cons;
    extern constraint default_io_diffCommits_info_199_rfWen_cons;
    extern constraint default_io_diffCommits_info_199_fpWen_cons;
    extern constraint default_io_diffCommits_info_199_vecWen_cons;
    extern constraint default_io_diffCommits_info_199_v0Wen_cons;
    extern constraint default_io_diffCommits_info_199_vlWen_cons;
    extern constraint default_io_diffCommits_info_200_ldest_cons;
    extern constraint default_io_diffCommits_info_200_pdest_cons;
    extern constraint default_io_diffCommits_info_200_rfWen_cons;
    extern constraint default_io_diffCommits_info_200_fpWen_cons;
    extern constraint default_io_diffCommits_info_200_vecWen_cons;
    extern constraint default_io_diffCommits_info_200_v0Wen_cons;
    extern constraint default_io_diffCommits_info_200_vlWen_cons;
    extern constraint default_io_diffCommits_info_201_ldest_cons;
    extern constraint default_io_diffCommits_info_201_pdest_cons;
    extern constraint default_io_diffCommits_info_201_rfWen_cons;
    extern constraint default_io_diffCommits_info_201_fpWen_cons;
    extern constraint default_io_diffCommits_info_201_vecWen_cons;
    extern constraint default_io_diffCommits_info_201_v0Wen_cons;
    extern constraint default_io_diffCommits_info_201_vlWen_cons;
    extern constraint default_io_diffCommits_info_202_ldest_cons;
    extern constraint default_io_diffCommits_info_202_pdest_cons;
    extern constraint default_io_diffCommits_info_202_rfWen_cons;
    extern constraint default_io_diffCommits_info_202_fpWen_cons;
    extern constraint default_io_diffCommits_info_202_vecWen_cons;
    extern constraint default_io_diffCommits_info_202_v0Wen_cons;
    extern constraint default_io_diffCommits_info_202_vlWen_cons;
    extern constraint default_io_diffCommits_info_203_ldest_cons;
    extern constraint default_io_diffCommits_info_203_pdest_cons;
    extern constraint default_io_diffCommits_info_203_rfWen_cons;
    extern constraint default_io_diffCommits_info_203_fpWen_cons;
    extern constraint default_io_diffCommits_info_203_vecWen_cons;
    extern constraint default_io_diffCommits_info_203_v0Wen_cons;
    extern constraint default_io_diffCommits_info_203_vlWen_cons;
    extern constraint default_io_diffCommits_info_204_ldest_cons;
    extern constraint default_io_diffCommits_info_204_pdest_cons;
    extern constraint default_io_diffCommits_info_204_rfWen_cons;
    extern constraint default_io_diffCommits_info_204_fpWen_cons;
    extern constraint default_io_diffCommits_info_204_vecWen_cons;
    extern constraint default_io_diffCommits_info_204_v0Wen_cons;
    extern constraint default_io_diffCommits_info_204_vlWen_cons;
    extern constraint default_io_diffCommits_info_205_ldest_cons;
    extern constraint default_io_diffCommits_info_205_pdest_cons;
    extern constraint default_io_diffCommits_info_205_rfWen_cons;
    extern constraint default_io_diffCommits_info_205_fpWen_cons;
    extern constraint default_io_diffCommits_info_205_vecWen_cons;
    extern constraint default_io_diffCommits_info_205_v0Wen_cons;
    extern constraint default_io_diffCommits_info_205_vlWen_cons;
    extern constraint default_io_diffCommits_info_206_ldest_cons;
    extern constraint default_io_diffCommits_info_206_pdest_cons;
    extern constraint default_io_diffCommits_info_206_rfWen_cons;
    extern constraint default_io_diffCommits_info_206_fpWen_cons;
    extern constraint default_io_diffCommits_info_206_vecWen_cons;
    extern constraint default_io_diffCommits_info_206_v0Wen_cons;
    extern constraint default_io_diffCommits_info_206_vlWen_cons;
    extern constraint default_io_diffCommits_info_207_ldest_cons;
    extern constraint default_io_diffCommits_info_207_pdest_cons;
    extern constraint default_io_diffCommits_info_207_rfWen_cons;
    extern constraint default_io_diffCommits_info_207_fpWen_cons;
    extern constraint default_io_diffCommits_info_207_vecWen_cons;
    extern constraint default_io_diffCommits_info_207_v0Wen_cons;
    extern constraint default_io_diffCommits_info_207_vlWen_cons;
    extern constraint default_io_diffCommits_info_208_ldest_cons;
    extern constraint default_io_diffCommits_info_208_pdest_cons;
    extern constraint default_io_diffCommits_info_208_rfWen_cons;
    extern constraint default_io_diffCommits_info_208_fpWen_cons;
    extern constraint default_io_diffCommits_info_208_vecWen_cons;
    extern constraint default_io_diffCommits_info_208_v0Wen_cons;
    extern constraint default_io_diffCommits_info_208_vlWen_cons;
    extern constraint default_io_diffCommits_info_209_ldest_cons;
    extern constraint default_io_diffCommits_info_209_pdest_cons;
    extern constraint default_io_diffCommits_info_209_rfWen_cons;
    extern constraint default_io_diffCommits_info_209_fpWen_cons;
    extern constraint default_io_diffCommits_info_209_vecWen_cons;
    extern constraint default_io_diffCommits_info_209_v0Wen_cons;
    extern constraint default_io_diffCommits_info_209_vlWen_cons;
    extern constraint default_io_diffCommits_info_210_ldest_cons;
    extern constraint default_io_diffCommits_info_210_pdest_cons;
    extern constraint default_io_diffCommits_info_210_rfWen_cons;
    extern constraint default_io_diffCommits_info_210_fpWen_cons;
    extern constraint default_io_diffCommits_info_210_vecWen_cons;
    extern constraint default_io_diffCommits_info_210_v0Wen_cons;
    extern constraint default_io_diffCommits_info_210_vlWen_cons;
    extern constraint default_io_diffCommits_info_211_ldest_cons;
    extern constraint default_io_diffCommits_info_211_pdest_cons;
    extern constraint default_io_diffCommits_info_211_rfWen_cons;
    extern constraint default_io_diffCommits_info_211_fpWen_cons;
    extern constraint default_io_diffCommits_info_211_vecWen_cons;
    extern constraint default_io_diffCommits_info_211_v0Wen_cons;
    extern constraint default_io_diffCommits_info_211_vlWen_cons;
    extern constraint default_io_diffCommits_info_212_ldest_cons;
    extern constraint default_io_diffCommits_info_212_pdest_cons;
    extern constraint default_io_diffCommits_info_212_rfWen_cons;
    extern constraint default_io_diffCommits_info_212_fpWen_cons;
    extern constraint default_io_diffCommits_info_212_vecWen_cons;
    extern constraint default_io_diffCommits_info_212_v0Wen_cons;
    extern constraint default_io_diffCommits_info_212_vlWen_cons;
    extern constraint default_io_diffCommits_info_213_ldest_cons;
    extern constraint default_io_diffCommits_info_213_pdest_cons;
    extern constraint default_io_diffCommits_info_213_rfWen_cons;
    extern constraint default_io_diffCommits_info_213_fpWen_cons;
    extern constraint default_io_diffCommits_info_213_vecWen_cons;
    extern constraint default_io_diffCommits_info_213_v0Wen_cons;
    extern constraint default_io_diffCommits_info_213_vlWen_cons;
    extern constraint default_io_diffCommits_info_214_ldest_cons;
    extern constraint default_io_diffCommits_info_214_pdest_cons;
    extern constraint default_io_diffCommits_info_214_rfWen_cons;
    extern constraint default_io_diffCommits_info_214_fpWen_cons;
    extern constraint default_io_diffCommits_info_214_vecWen_cons;
    extern constraint default_io_diffCommits_info_214_v0Wen_cons;
    extern constraint default_io_diffCommits_info_214_vlWen_cons;
    extern constraint default_io_diffCommits_info_215_ldest_cons;
    extern constraint default_io_diffCommits_info_215_pdest_cons;
    extern constraint default_io_diffCommits_info_215_rfWen_cons;
    extern constraint default_io_diffCommits_info_215_fpWen_cons;
    extern constraint default_io_diffCommits_info_215_vecWen_cons;
    extern constraint default_io_diffCommits_info_215_v0Wen_cons;
    extern constraint default_io_diffCommits_info_215_vlWen_cons;
    extern constraint default_io_diffCommits_info_216_ldest_cons;
    extern constraint default_io_diffCommits_info_216_pdest_cons;
    extern constraint default_io_diffCommits_info_216_rfWen_cons;
    extern constraint default_io_diffCommits_info_216_fpWen_cons;
    extern constraint default_io_diffCommits_info_216_vecWen_cons;
    extern constraint default_io_diffCommits_info_216_v0Wen_cons;
    extern constraint default_io_diffCommits_info_216_vlWen_cons;
    extern constraint default_io_diffCommits_info_217_ldest_cons;
    extern constraint default_io_diffCommits_info_217_pdest_cons;
    extern constraint default_io_diffCommits_info_217_rfWen_cons;
    extern constraint default_io_diffCommits_info_217_fpWen_cons;
    extern constraint default_io_diffCommits_info_217_vecWen_cons;
    extern constraint default_io_diffCommits_info_217_v0Wen_cons;
    extern constraint default_io_diffCommits_info_217_vlWen_cons;
    extern constraint default_io_diffCommits_info_218_ldest_cons;
    extern constraint default_io_diffCommits_info_218_pdest_cons;
    extern constraint default_io_diffCommits_info_218_rfWen_cons;
    extern constraint default_io_diffCommits_info_218_fpWen_cons;
    extern constraint default_io_diffCommits_info_218_vecWen_cons;
    extern constraint default_io_diffCommits_info_218_v0Wen_cons;
    extern constraint default_io_diffCommits_info_218_vlWen_cons;
    extern constraint default_io_diffCommits_info_219_ldest_cons;
    extern constraint default_io_diffCommits_info_219_pdest_cons;
    extern constraint default_io_diffCommits_info_219_rfWen_cons;
    extern constraint default_io_diffCommits_info_219_fpWen_cons;
    extern constraint default_io_diffCommits_info_219_vecWen_cons;
    extern constraint default_io_diffCommits_info_219_v0Wen_cons;
    extern constraint default_io_diffCommits_info_219_vlWen_cons;
    extern constraint default_io_diffCommits_info_220_ldest_cons;
    extern constraint default_io_diffCommits_info_220_pdest_cons;
    extern constraint default_io_diffCommits_info_220_rfWen_cons;
    extern constraint default_io_diffCommits_info_220_fpWen_cons;
    extern constraint default_io_diffCommits_info_220_vecWen_cons;
    extern constraint default_io_diffCommits_info_220_v0Wen_cons;
    extern constraint default_io_diffCommits_info_220_vlWen_cons;
    extern constraint default_io_diffCommits_info_221_ldest_cons;
    extern constraint default_io_diffCommits_info_221_pdest_cons;
    extern constraint default_io_diffCommits_info_221_rfWen_cons;
    extern constraint default_io_diffCommits_info_221_fpWen_cons;
    extern constraint default_io_diffCommits_info_221_vecWen_cons;
    extern constraint default_io_diffCommits_info_221_v0Wen_cons;
    extern constraint default_io_diffCommits_info_221_vlWen_cons;
    extern constraint default_io_diffCommits_info_222_ldest_cons;
    extern constraint default_io_diffCommits_info_222_pdest_cons;
    extern constraint default_io_diffCommits_info_222_rfWen_cons;
    extern constraint default_io_diffCommits_info_222_fpWen_cons;
    extern constraint default_io_diffCommits_info_222_vecWen_cons;
    extern constraint default_io_diffCommits_info_222_v0Wen_cons;
    extern constraint default_io_diffCommits_info_222_vlWen_cons;
    extern constraint default_io_diffCommits_info_223_ldest_cons;
    extern constraint default_io_diffCommits_info_223_pdest_cons;
    extern constraint default_io_diffCommits_info_223_rfWen_cons;
    extern constraint default_io_diffCommits_info_223_fpWen_cons;
    extern constraint default_io_diffCommits_info_223_vecWen_cons;
    extern constraint default_io_diffCommits_info_223_v0Wen_cons;
    extern constraint default_io_diffCommits_info_223_vlWen_cons;
    extern constraint default_io_diffCommits_info_224_ldest_cons;
    extern constraint default_io_diffCommits_info_224_pdest_cons;
    extern constraint default_io_diffCommits_info_224_rfWen_cons;
    extern constraint default_io_diffCommits_info_224_fpWen_cons;
    extern constraint default_io_diffCommits_info_224_vecWen_cons;
    extern constraint default_io_diffCommits_info_224_v0Wen_cons;
    extern constraint default_io_diffCommits_info_224_vlWen_cons;
    extern constraint default_io_diffCommits_info_225_ldest_cons;
    extern constraint default_io_diffCommits_info_225_pdest_cons;
    extern constraint default_io_diffCommits_info_225_rfWen_cons;
    extern constraint default_io_diffCommits_info_225_fpWen_cons;
    extern constraint default_io_diffCommits_info_225_vecWen_cons;
    extern constraint default_io_diffCommits_info_225_v0Wen_cons;
    extern constraint default_io_diffCommits_info_225_vlWen_cons;
    extern constraint default_io_diffCommits_info_226_ldest_cons;
    extern constraint default_io_diffCommits_info_226_pdest_cons;
    extern constraint default_io_diffCommits_info_226_rfWen_cons;
    extern constraint default_io_diffCommits_info_226_fpWen_cons;
    extern constraint default_io_diffCommits_info_226_vecWen_cons;
    extern constraint default_io_diffCommits_info_226_v0Wen_cons;
    extern constraint default_io_diffCommits_info_226_vlWen_cons;
    extern constraint default_io_diffCommits_info_227_ldest_cons;
    extern constraint default_io_diffCommits_info_227_pdest_cons;
    extern constraint default_io_diffCommits_info_227_rfWen_cons;
    extern constraint default_io_diffCommits_info_227_fpWen_cons;
    extern constraint default_io_diffCommits_info_227_vecWen_cons;
    extern constraint default_io_diffCommits_info_227_v0Wen_cons;
    extern constraint default_io_diffCommits_info_227_vlWen_cons;
    extern constraint default_io_diffCommits_info_228_ldest_cons;
    extern constraint default_io_diffCommits_info_228_pdest_cons;
    extern constraint default_io_diffCommits_info_228_rfWen_cons;
    extern constraint default_io_diffCommits_info_228_fpWen_cons;
    extern constraint default_io_diffCommits_info_228_vecWen_cons;
    extern constraint default_io_diffCommits_info_228_v0Wen_cons;
    extern constraint default_io_diffCommits_info_228_vlWen_cons;
    extern constraint default_io_diffCommits_info_229_ldest_cons;
    extern constraint default_io_diffCommits_info_229_pdest_cons;
    extern constraint default_io_diffCommits_info_229_rfWen_cons;
    extern constraint default_io_diffCommits_info_229_fpWen_cons;
    extern constraint default_io_diffCommits_info_229_vecWen_cons;
    extern constraint default_io_diffCommits_info_229_v0Wen_cons;
    extern constraint default_io_diffCommits_info_229_vlWen_cons;
    extern constraint default_io_diffCommits_info_230_ldest_cons;
    extern constraint default_io_diffCommits_info_230_pdest_cons;
    extern constraint default_io_diffCommits_info_230_rfWen_cons;
    extern constraint default_io_diffCommits_info_230_fpWen_cons;
    extern constraint default_io_diffCommits_info_230_vecWen_cons;
    extern constraint default_io_diffCommits_info_230_v0Wen_cons;
    extern constraint default_io_diffCommits_info_230_vlWen_cons;
    extern constraint default_io_diffCommits_info_231_ldest_cons;
    extern constraint default_io_diffCommits_info_231_pdest_cons;
    extern constraint default_io_diffCommits_info_231_rfWen_cons;
    extern constraint default_io_diffCommits_info_231_fpWen_cons;
    extern constraint default_io_diffCommits_info_231_vecWen_cons;
    extern constraint default_io_diffCommits_info_231_v0Wen_cons;
    extern constraint default_io_diffCommits_info_231_vlWen_cons;
    extern constraint default_io_diffCommits_info_232_ldest_cons;
    extern constraint default_io_diffCommits_info_232_pdest_cons;
    extern constraint default_io_diffCommits_info_232_rfWen_cons;
    extern constraint default_io_diffCommits_info_232_fpWen_cons;
    extern constraint default_io_diffCommits_info_232_vecWen_cons;
    extern constraint default_io_diffCommits_info_232_v0Wen_cons;
    extern constraint default_io_diffCommits_info_232_vlWen_cons;
    extern constraint default_io_diffCommits_info_233_ldest_cons;
    extern constraint default_io_diffCommits_info_233_pdest_cons;
    extern constraint default_io_diffCommits_info_233_rfWen_cons;
    extern constraint default_io_diffCommits_info_233_fpWen_cons;
    extern constraint default_io_diffCommits_info_233_vecWen_cons;
    extern constraint default_io_diffCommits_info_233_v0Wen_cons;
    extern constraint default_io_diffCommits_info_233_vlWen_cons;
    extern constraint default_io_diffCommits_info_234_ldest_cons;
    extern constraint default_io_diffCommits_info_234_pdest_cons;
    extern constraint default_io_diffCommits_info_234_rfWen_cons;
    extern constraint default_io_diffCommits_info_234_fpWen_cons;
    extern constraint default_io_diffCommits_info_234_vecWen_cons;
    extern constraint default_io_diffCommits_info_234_v0Wen_cons;
    extern constraint default_io_diffCommits_info_234_vlWen_cons;
    extern constraint default_io_diffCommits_info_235_ldest_cons;
    extern constraint default_io_diffCommits_info_235_pdest_cons;
    extern constraint default_io_diffCommits_info_235_rfWen_cons;
    extern constraint default_io_diffCommits_info_235_fpWen_cons;
    extern constraint default_io_diffCommits_info_235_vecWen_cons;
    extern constraint default_io_diffCommits_info_235_v0Wen_cons;
    extern constraint default_io_diffCommits_info_235_vlWen_cons;
    extern constraint default_io_diffCommits_info_236_ldest_cons;
    extern constraint default_io_diffCommits_info_236_pdest_cons;
    extern constraint default_io_diffCommits_info_236_rfWen_cons;
    extern constraint default_io_diffCommits_info_236_fpWen_cons;
    extern constraint default_io_diffCommits_info_236_vecWen_cons;
    extern constraint default_io_diffCommits_info_236_v0Wen_cons;
    extern constraint default_io_diffCommits_info_236_vlWen_cons;
    extern constraint default_io_diffCommits_info_237_ldest_cons;
    extern constraint default_io_diffCommits_info_237_pdest_cons;
    extern constraint default_io_diffCommits_info_237_rfWen_cons;
    extern constraint default_io_diffCommits_info_237_fpWen_cons;
    extern constraint default_io_diffCommits_info_237_vecWen_cons;
    extern constraint default_io_diffCommits_info_237_v0Wen_cons;
    extern constraint default_io_diffCommits_info_237_vlWen_cons;
    extern constraint default_io_diffCommits_info_238_ldest_cons;
    extern constraint default_io_diffCommits_info_238_pdest_cons;
    extern constraint default_io_diffCommits_info_238_rfWen_cons;
    extern constraint default_io_diffCommits_info_238_fpWen_cons;
    extern constraint default_io_diffCommits_info_238_vecWen_cons;
    extern constraint default_io_diffCommits_info_238_v0Wen_cons;
    extern constraint default_io_diffCommits_info_238_vlWen_cons;
    extern constraint default_io_diffCommits_info_239_ldest_cons;
    extern constraint default_io_diffCommits_info_239_pdest_cons;
    extern constraint default_io_diffCommits_info_239_rfWen_cons;
    extern constraint default_io_diffCommits_info_239_fpWen_cons;
    extern constraint default_io_diffCommits_info_239_vecWen_cons;
    extern constraint default_io_diffCommits_info_239_v0Wen_cons;
    extern constraint default_io_diffCommits_info_239_vlWen_cons;
    extern constraint default_io_diffCommits_info_240_ldest_cons;
    extern constraint default_io_diffCommits_info_240_pdest_cons;
    extern constraint default_io_diffCommits_info_240_rfWen_cons;
    extern constraint default_io_diffCommits_info_240_fpWen_cons;
    extern constraint default_io_diffCommits_info_240_vecWen_cons;
    extern constraint default_io_diffCommits_info_240_v0Wen_cons;
    extern constraint default_io_diffCommits_info_240_vlWen_cons;
    extern constraint default_io_diffCommits_info_241_ldest_cons;
    extern constraint default_io_diffCommits_info_241_pdest_cons;
    extern constraint default_io_diffCommits_info_241_rfWen_cons;
    extern constraint default_io_diffCommits_info_241_fpWen_cons;
    extern constraint default_io_diffCommits_info_241_vecWen_cons;
    extern constraint default_io_diffCommits_info_241_v0Wen_cons;
    extern constraint default_io_diffCommits_info_241_vlWen_cons;
    extern constraint default_io_diffCommits_info_242_ldest_cons;
    extern constraint default_io_diffCommits_info_242_pdest_cons;
    extern constraint default_io_diffCommits_info_242_rfWen_cons;
    extern constraint default_io_diffCommits_info_242_fpWen_cons;
    extern constraint default_io_diffCommits_info_242_vecWen_cons;
    extern constraint default_io_diffCommits_info_242_v0Wen_cons;
    extern constraint default_io_diffCommits_info_242_vlWen_cons;
    extern constraint default_io_diffCommits_info_243_ldest_cons;
    extern constraint default_io_diffCommits_info_243_pdest_cons;
    extern constraint default_io_diffCommits_info_243_rfWen_cons;
    extern constraint default_io_diffCommits_info_243_fpWen_cons;
    extern constraint default_io_diffCommits_info_243_vecWen_cons;
    extern constraint default_io_diffCommits_info_243_v0Wen_cons;
    extern constraint default_io_diffCommits_info_243_vlWen_cons;
    extern constraint default_io_diffCommits_info_244_ldest_cons;
    extern constraint default_io_diffCommits_info_244_pdest_cons;
    extern constraint default_io_diffCommits_info_244_rfWen_cons;
    extern constraint default_io_diffCommits_info_244_fpWen_cons;
    extern constraint default_io_diffCommits_info_244_vecWen_cons;
    extern constraint default_io_diffCommits_info_244_v0Wen_cons;
    extern constraint default_io_diffCommits_info_244_vlWen_cons;
    extern constraint default_io_diffCommits_info_245_ldest_cons;
    extern constraint default_io_diffCommits_info_245_pdest_cons;
    extern constraint default_io_diffCommits_info_245_rfWen_cons;
    extern constraint default_io_diffCommits_info_245_fpWen_cons;
    extern constraint default_io_diffCommits_info_245_vecWen_cons;
    extern constraint default_io_diffCommits_info_245_v0Wen_cons;
    extern constraint default_io_diffCommits_info_245_vlWen_cons;
    extern constraint default_io_diffCommits_info_246_ldest_cons;
    extern constraint default_io_diffCommits_info_246_pdest_cons;
    extern constraint default_io_diffCommits_info_246_rfWen_cons;
    extern constraint default_io_diffCommits_info_246_fpWen_cons;
    extern constraint default_io_diffCommits_info_246_vecWen_cons;
    extern constraint default_io_diffCommits_info_246_v0Wen_cons;
    extern constraint default_io_diffCommits_info_246_vlWen_cons;
    extern constraint default_io_diffCommits_info_247_ldest_cons;
    extern constraint default_io_diffCommits_info_247_pdest_cons;
    extern constraint default_io_diffCommits_info_247_rfWen_cons;
    extern constraint default_io_diffCommits_info_247_fpWen_cons;
    extern constraint default_io_diffCommits_info_247_vecWen_cons;
    extern constraint default_io_diffCommits_info_247_v0Wen_cons;
    extern constraint default_io_diffCommits_info_247_vlWen_cons;
    extern constraint default_io_diffCommits_info_248_ldest_cons;
    extern constraint default_io_diffCommits_info_248_pdest_cons;
    extern constraint default_io_diffCommits_info_248_rfWen_cons;
    extern constraint default_io_diffCommits_info_248_fpWen_cons;
    extern constraint default_io_diffCommits_info_248_vecWen_cons;
    extern constraint default_io_diffCommits_info_248_v0Wen_cons;
    extern constraint default_io_diffCommits_info_248_vlWen_cons;
    extern constraint default_io_diffCommits_info_249_ldest_cons;
    extern constraint default_io_diffCommits_info_249_pdest_cons;
    extern constraint default_io_diffCommits_info_249_rfWen_cons;
    extern constraint default_io_diffCommits_info_249_fpWen_cons;
    extern constraint default_io_diffCommits_info_249_vecWen_cons;
    extern constraint default_io_diffCommits_info_249_v0Wen_cons;
    extern constraint default_io_diffCommits_info_249_vlWen_cons;
    extern constraint default_io_diffCommits_info_250_ldest_cons;
    extern constraint default_io_diffCommits_info_250_pdest_cons;
    extern constraint default_io_diffCommits_info_250_rfWen_cons;
    extern constraint default_io_diffCommits_info_250_fpWen_cons;
    extern constraint default_io_diffCommits_info_250_vecWen_cons;
    extern constraint default_io_diffCommits_info_250_v0Wen_cons;
    extern constraint default_io_diffCommits_info_250_vlWen_cons;
    extern constraint default_io_diffCommits_info_251_ldest_cons;
    extern constraint default_io_diffCommits_info_251_pdest_cons;
    extern constraint default_io_diffCommits_info_251_rfWen_cons;
    extern constraint default_io_diffCommits_info_251_fpWen_cons;
    extern constraint default_io_diffCommits_info_251_vecWen_cons;
    extern constraint default_io_diffCommits_info_251_v0Wen_cons;
    extern constraint default_io_diffCommits_info_251_vlWen_cons;
    extern constraint default_io_diffCommits_info_252_ldest_cons;
    extern constraint default_io_diffCommits_info_252_pdest_cons;
    extern constraint default_io_diffCommits_info_252_rfWen_cons;
    extern constraint default_io_diffCommits_info_252_fpWen_cons;
    extern constraint default_io_diffCommits_info_252_vecWen_cons;
    extern constraint default_io_diffCommits_info_252_v0Wen_cons;
    extern constraint default_io_diffCommits_info_252_vlWen_cons;
    extern constraint default_io_diffCommits_info_253_ldest_cons;
    extern constraint default_io_diffCommits_info_253_pdest_cons;
    extern constraint default_io_diffCommits_info_253_rfWen_cons;
    extern constraint default_io_diffCommits_info_253_fpWen_cons;
    extern constraint default_io_diffCommits_info_253_vecWen_cons;
    extern constraint default_io_diffCommits_info_253_v0Wen_cons;
    extern constraint default_io_diffCommits_info_253_vlWen_cons;
    extern constraint default_io_diffCommits_info_254_ldest_cons;
    extern constraint default_io_diffCommits_info_254_pdest_cons;
    extern constraint default_io_diffCommits_info_254_rfWen_cons;
    extern constraint default_io_diffCommits_info_254_fpWen_cons;
    extern constraint default_io_diffCommits_info_254_vecWen_cons;
    extern constraint default_io_diffCommits_info_254_v0Wen_cons;
    extern constraint default_io_diffCommits_info_254_vlWen_cons;
    extern constraint default_io_diffCommits_info_255_ldest_cons;
    extern constraint default_io_diffCommits_info_255_pdest_cons;
    extern constraint default_io_diffCommits_info_256_ldest_cons;
    extern constraint default_io_diffCommits_info_256_pdest_cons;
    extern constraint default_io_diffCommits_info_257_ldest_cons;
    extern constraint default_io_diffCommits_info_257_pdest_cons;
    extern constraint default_io_diffCommits_info_258_ldest_cons;
    extern constraint default_io_diffCommits_info_258_pdest_cons;
    extern constraint default_io_diffCommits_info_259_ldest_cons;
    extern constraint default_io_diffCommits_info_259_pdest_cons;
    extern constraint default_io_diffCommits_info_260_ldest_cons;
    extern constraint default_io_diffCommits_info_260_pdest_cons;
    extern constraint default_io_diffCommits_info_261_ldest_cons;
    extern constraint default_io_diffCommits_info_261_pdest_cons;
    extern constraint default_io_diffCommits_info_262_ldest_cons;
    extern constraint default_io_diffCommits_info_262_pdest_cons;
    extern constraint default_io_diffCommits_info_263_ldest_cons;
    extern constraint default_io_diffCommits_info_263_pdest_cons;
    extern constraint default_io_diffCommits_info_264_ldest_cons;
    extern constraint default_io_diffCommits_info_264_pdest_cons;
    extern constraint default_io_diffCommits_info_265_ldest_cons;
    extern constraint default_io_diffCommits_info_265_pdest_cons;
    extern constraint default_io_diffCommits_info_266_ldest_cons;
    extern constraint default_io_diffCommits_info_266_pdest_cons;
    extern constraint default_io_diffCommits_info_267_ldest_cons;
    extern constraint default_io_diffCommits_info_267_pdest_cons;
    extern constraint default_io_diffCommits_info_268_ldest_cons;
    extern constraint default_io_diffCommits_info_268_pdest_cons;
    extern constraint default_io_diffCommits_info_269_ldest_cons;
    extern constraint default_io_diffCommits_info_269_pdest_cons;
    extern constraint default_io_diffCommits_info_270_ldest_cons;
    extern constraint default_io_diffCommits_info_270_pdest_cons;
    extern constraint default_io_diffCommits_info_271_ldest_cons;
    extern constraint default_io_diffCommits_info_271_pdest_cons;
    extern constraint default_io_diffCommits_info_272_ldest_cons;
    extern constraint default_io_diffCommits_info_272_pdest_cons;
    extern constraint default_io_diffCommits_info_273_ldest_cons;
    extern constraint default_io_diffCommits_info_273_pdest_cons;
    extern constraint default_io_diffCommits_info_274_ldest_cons;
    extern constraint default_io_diffCommits_info_274_pdest_cons;
    extern constraint default_io_diffCommits_info_275_ldest_cons;
    extern constraint default_io_diffCommits_info_275_pdest_cons;
    extern constraint default_io_diffCommits_info_276_ldest_cons;
    extern constraint default_io_diffCommits_info_276_pdest_cons;
    extern constraint default_io_diffCommits_info_277_ldest_cons;
    extern constraint default_io_diffCommits_info_277_pdest_cons;
    extern constraint default_io_diffCommits_info_278_ldest_cons;
    extern constraint default_io_diffCommits_info_278_pdest_cons;
    extern constraint default_io_diffCommits_info_279_ldest_cons;
    extern constraint default_io_diffCommits_info_279_pdest_cons;
    extern constraint default_io_diffCommits_info_280_ldest_cons;
    extern constraint default_io_diffCommits_info_280_pdest_cons;
    extern constraint default_io_diffCommits_info_281_ldest_cons;
    extern constraint default_io_diffCommits_info_281_pdest_cons;
    extern constraint default_io_diffCommits_info_282_ldest_cons;
    extern constraint default_io_diffCommits_info_282_pdest_cons;
    extern constraint default_io_diffCommits_info_283_ldest_cons;
    extern constraint default_io_diffCommits_info_283_pdest_cons;
    extern constraint default_io_diffCommits_info_284_ldest_cons;
    extern constraint default_io_diffCommits_info_284_pdest_cons;
    extern constraint default_io_diffCommits_info_285_ldest_cons;
    extern constraint default_io_diffCommits_info_285_pdest_cons;
    extern constraint default_io_diffCommits_info_286_ldest_cons;
    extern constraint default_io_diffCommits_info_286_pdest_cons;
    extern constraint default_io_diffCommits_info_287_ldest_cons;
    extern constraint default_io_diffCommits_info_287_pdest_cons;
    extern constraint default_io_diffCommits_info_288_ldest_cons;
    extern constraint default_io_diffCommits_info_288_pdest_cons;
    extern constraint default_io_diffCommits_info_289_ldest_cons;
    extern constraint default_io_diffCommits_info_289_pdest_cons;
    extern constraint default_io_diffCommits_info_290_ldest_cons;
    extern constraint default_io_diffCommits_info_290_pdest_cons;
    extern constraint default_io_diffCommits_info_291_ldest_cons;
    extern constraint default_io_diffCommits_info_291_pdest_cons;
    extern constraint default_io_diffCommits_info_292_ldest_cons;
    extern constraint default_io_diffCommits_info_292_pdest_cons;
    extern constraint default_io_diffCommits_info_293_ldest_cons;
    extern constraint default_io_diffCommits_info_293_pdest_cons;
    extern constraint default_io_diffCommits_info_294_ldest_cons;
    extern constraint default_io_diffCommits_info_294_pdest_cons;
    extern constraint default_io_diffCommits_info_295_ldest_cons;
    extern constraint default_io_diffCommits_info_295_pdest_cons;
    extern constraint default_io_diffCommits_info_296_ldest_cons;
    extern constraint default_io_diffCommits_info_296_pdest_cons;
    extern constraint default_io_diffCommits_info_297_ldest_cons;
    extern constraint default_io_diffCommits_info_297_pdest_cons;
    extern constraint default_io_diffCommits_info_298_ldest_cons;
    extern constraint default_io_diffCommits_info_298_pdest_cons;
    extern constraint default_io_diffCommits_info_299_ldest_cons;
    extern constraint default_io_diffCommits_info_299_pdest_cons;
    extern constraint default_io_diffCommits_info_300_ldest_cons;
    extern constraint default_io_diffCommits_info_300_pdest_cons;
    extern constraint default_io_diffCommits_info_301_ldest_cons;
    extern constraint default_io_diffCommits_info_301_pdest_cons;
    extern constraint default_io_diffCommits_info_302_ldest_cons;
    extern constraint default_io_diffCommits_info_302_pdest_cons;
    extern constraint default_io_diffCommits_info_303_ldest_cons;
    extern constraint default_io_diffCommits_info_303_pdest_cons;
    extern constraint default_io_diffCommits_info_304_ldest_cons;
    extern constraint default_io_diffCommits_info_304_pdest_cons;
    extern constraint default_io_diffCommits_info_305_ldest_cons;
    extern constraint default_io_diffCommits_info_305_pdest_cons;
    extern constraint default_io_diffCommits_info_306_ldest_cons;
    extern constraint default_io_diffCommits_info_306_pdest_cons;
    extern constraint default_io_diffCommits_info_307_ldest_cons;
    extern constraint default_io_diffCommits_info_307_pdest_cons;
    extern constraint default_io_diffCommits_info_308_ldest_cons;
    extern constraint default_io_diffCommits_info_308_pdest_cons;
    extern constraint default_io_diffCommits_info_309_ldest_cons;
    extern constraint default_io_diffCommits_info_309_pdest_cons;
    extern constraint default_io_diffCommits_info_310_ldest_cons;
    extern constraint default_io_diffCommits_info_310_pdest_cons;
    extern constraint default_io_diffCommits_info_311_ldest_cons;
    extern constraint default_io_diffCommits_info_311_pdest_cons;
    extern constraint default_io_diffCommits_info_312_ldest_cons;
    extern constraint default_io_diffCommits_info_312_pdest_cons;
    extern constraint default_io_diffCommits_info_313_ldest_cons;
    extern constraint default_io_diffCommits_info_313_pdest_cons;
    extern constraint default_io_diffCommits_info_314_ldest_cons;
    extern constraint default_io_diffCommits_info_314_pdest_cons;
    extern constraint default_io_diffCommits_info_315_ldest_cons;
    extern constraint default_io_diffCommits_info_315_pdest_cons;
    extern constraint default_io_diffCommits_info_316_ldest_cons;
    extern constraint default_io_diffCommits_info_316_pdest_cons;
    extern constraint default_io_diffCommits_info_317_ldest_cons;
    extern constraint default_io_diffCommits_info_317_pdest_cons;
    extern constraint default_io_diffCommits_info_318_ldest_cons;
    extern constraint default_io_diffCommits_info_318_pdest_cons;
    extern constraint default_io_diffCommits_info_319_ldest_cons;
    extern constraint default_io_diffCommits_info_319_pdest_cons;
    extern constraint default_io_diffCommits_info_320_ldest_cons;
    extern constraint default_io_diffCommits_info_320_pdest_cons;
    extern constraint default_io_diffCommits_info_321_ldest_cons;
    extern constraint default_io_diffCommits_info_321_pdest_cons;
    extern constraint default_io_diffCommits_info_322_ldest_cons;
    extern constraint default_io_diffCommits_info_322_pdest_cons;
    extern constraint default_io_diffCommits_info_323_ldest_cons;
    extern constraint default_io_diffCommits_info_323_pdest_cons;
    extern constraint default_io_diffCommits_info_324_ldest_cons;
    extern constraint default_io_diffCommits_info_324_pdest_cons;
    extern constraint default_io_diffCommits_info_325_ldest_cons;
    extern constraint default_io_diffCommits_info_325_pdest_cons;
    extern constraint default_io_diffCommits_info_326_ldest_cons;
    extern constraint default_io_diffCommits_info_326_pdest_cons;
    extern constraint default_io_diffCommits_info_327_ldest_cons;
    extern constraint default_io_diffCommits_info_327_pdest_cons;
    extern constraint default_io_diffCommits_info_328_ldest_cons;
    extern constraint default_io_diffCommits_info_328_pdest_cons;
    extern constraint default_io_diffCommits_info_329_ldest_cons;
    extern constraint default_io_diffCommits_info_329_pdest_cons;
    extern constraint default_io_diffCommits_info_330_ldest_cons;
    extern constraint default_io_diffCommits_info_330_pdest_cons;
    extern constraint default_io_diffCommits_info_331_ldest_cons;
    extern constraint default_io_diffCommits_info_331_pdest_cons;
    extern constraint default_io_diffCommits_info_332_ldest_cons;
    extern constraint default_io_diffCommits_info_332_pdest_cons;
    extern constraint default_io_diffCommits_info_333_ldest_cons;
    extern constraint default_io_diffCommits_info_333_pdest_cons;
    extern constraint default_io_diffCommits_info_334_ldest_cons;
    extern constraint default_io_diffCommits_info_334_pdest_cons;
    extern constraint default_io_diffCommits_info_335_ldest_cons;
    extern constraint default_io_diffCommits_info_335_pdest_cons;
    extern constraint default_io_diffCommits_info_336_ldest_cons;
    extern constraint default_io_diffCommits_info_336_pdest_cons;
    extern constraint default_io_diffCommits_info_337_ldest_cons;
    extern constraint default_io_diffCommits_info_337_pdest_cons;
    extern constraint default_io_diffCommits_info_338_ldest_cons;
    extern constraint default_io_diffCommits_info_338_pdest_cons;
    extern constraint default_io_diffCommits_info_339_ldest_cons;
    extern constraint default_io_diffCommits_info_339_pdest_cons;
    extern constraint default_io_diffCommits_info_340_ldest_cons;
    extern constraint default_io_diffCommits_info_340_pdest_cons;
    extern constraint default_io_diffCommits_info_341_ldest_cons;
    extern constraint default_io_diffCommits_info_341_pdest_cons;
    extern constraint default_io_diffCommits_info_342_ldest_cons;
    extern constraint default_io_diffCommits_info_342_pdest_cons;
    extern constraint default_io_diffCommits_info_343_ldest_cons;
    extern constraint default_io_diffCommits_info_343_pdest_cons;
    extern constraint default_io_diffCommits_info_344_ldest_cons;
    extern constraint default_io_diffCommits_info_344_pdest_cons;
    extern constraint default_io_diffCommits_info_345_ldest_cons;
    extern constraint default_io_diffCommits_info_345_pdest_cons;
    extern constraint default_io_diffCommits_info_346_ldest_cons;
    extern constraint default_io_diffCommits_info_346_pdest_cons;
    extern constraint default_io_diffCommits_info_347_ldest_cons;
    extern constraint default_io_diffCommits_info_347_pdest_cons;
    extern constraint default_io_diffCommits_info_348_ldest_cons;
    extern constraint default_io_diffCommits_info_348_pdest_cons;
    extern constraint default_io_diffCommits_info_349_ldest_cons;
    extern constraint default_io_diffCommits_info_349_pdest_cons;
    extern constraint default_io_diffCommits_info_350_ldest_cons;
    extern constraint default_io_diffCommits_info_350_pdest_cons;
    extern constraint default_io_diffCommits_info_351_ldest_cons;
    extern constraint default_io_diffCommits_info_351_pdest_cons;
    extern constraint default_io_diffCommits_info_352_ldest_cons;
    extern constraint default_io_diffCommits_info_352_pdest_cons;
    extern constraint default_io_diffCommits_info_353_ldest_cons;
    extern constraint default_io_diffCommits_info_353_pdest_cons;
    extern constraint default_io_diffCommits_info_354_ldest_cons;
    extern constraint default_io_diffCommits_info_354_pdest_cons;
    extern constraint default_io_diffCommits_info_355_ldest_cons;
    extern constraint default_io_diffCommits_info_355_pdest_cons;
    extern constraint default_io_diffCommits_info_356_ldest_cons;
    extern constraint default_io_diffCommits_info_356_pdest_cons;
    extern constraint default_io_diffCommits_info_357_ldest_cons;
    extern constraint default_io_diffCommits_info_357_pdest_cons;
    extern constraint default_io_diffCommits_info_358_ldest_cons;
    extern constraint default_io_diffCommits_info_358_pdest_cons;
    extern constraint default_io_diffCommits_info_359_ldest_cons;
    extern constraint default_io_diffCommits_info_359_pdest_cons;
    extern constraint default_io_diffCommits_info_360_ldest_cons;
    extern constraint default_io_diffCommits_info_360_pdest_cons;
    extern constraint default_io_diffCommits_info_361_ldest_cons;
    extern constraint default_io_diffCommits_info_361_pdest_cons;
    extern constraint default_io_diffCommits_info_362_ldest_cons;
    extern constraint default_io_diffCommits_info_362_pdest_cons;
    extern constraint default_io_diffCommits_info_363_ldest_cons;
    extern constraint default_io_diffCommits_info_363_pdest_cons;
    extern constraint default_io_diffCommits_info_364_ldest_cons;
    extern constraint default_io_diffCommits_info_364_pdest_cons;
    extern constraint default_io_diffCommits_info_365_ldest_cons;
    extern constraint default_io_diffCommits_info_365_pdest_cons;
    extern constraint default_io_diffCommits_info_366_ldest_cons;
    extern constraint default_io_diffCommits_info_366_pdest_cons;
    extern constraint default_io_diffCommits_info_367_ldest_cons;
    extern constraint default_io_diffCommits_info_367_pdest_cons;
    extern constraint default_io_diffCommits_info_368_ldest_cons;
    extern constraint default_io_diffCommits_info_368_pdest_cons;
    extern constraint default_io_diffCommits_info_369_ldest_cons;
    extern constraint default_io_diffCommits_info_369_pdest_cons;
    extern constraint default_io_diffCommits_info_370_ldest_cons;
    extern constraint default_io_diffCommits_info_370_pdest_cons;
    extern constraint default_io_diffCommits_info_371_ldest_cons;
    extern constraint default_io_diffCommits_info_371_pdest_cons;
    extern constraint default_io_diffCommits_info_372_ldest_cons;
    extern constraint default_io_diffCommits_info_372_pdest_cons;
    extern constraint default_io_diffCommits_info_373_ldest_cons;
    extern constraint default_io_diffCommits_info_373_pdest_cons;
    extern constraint default_io_diffCommits_info_374_ldest_cons;
    extern constraint default_io_diffCommits_info_374_pdest_cons;
    extern constraint default_io_diffCommits_info_375_ldest_cons;
    extern constraint default_io_diffCommits_info_375_pdest_cons;
    extern constraint default_io_diffCommits_info_376_ldest_cons;
    extern constraint default_io_diffCommits_info_376_pdest_cons;
    extern constraint default_io_diffCommits_info_377_ldest_cons;
    extern constraint default_io_diffCommits_info_377_pdest_cons;
    extern constraint default_io_diffCommits_info_378_ldest_cons;
    extern constraint default_io_diffCommits_info_378_pdest_cons;
    extern constraint default_io_diffCommits_info_379_ldest_cons;
    extern constraint default_io_diffCommits_info_379_pdest_cons;
    extern constraint default_io_diffCommits_info_380_ldest_cons;
    extern constraint default_io_diffCommits_info_380_pdest_cons;
    extern constraint default_io_diffCommits_info_381_ldest_cons;
    extern constraint default_io_diffCommits_info_381_pdest_cons;
    extern constraint default_io_diffCommits_info_382_ldest_cons;
    extern constraint default_io_diffCommits_info_382_pdest_cons;
    extern constraint default_io_diffCommits_info_383_ldest_cons;
    extern constraint default_io_diffCommits_info_383_pdest_cons;
    extern constraint default_io_diffCommits_info_384_ldest_cons;
    extern constraint default_io_diffCommits_info_384_pdest_cons;
    extern constraint default_io_diffCommits_info_385_ldest_cons;
    extern constraint default_io_diffCommits_info_385_pdest_cons;
    extern constraint default_io_diffCommits_info_386_ldest_cons;
    extern constraint default_io_diffCommits_info_386_pdest_cons;
    extern constraint default_io_diffCommits_info_387_ldest_cons;
    extern constraint default_io_diffCommits_info_387_pdest_cons;
    extern constraint default_io_diffCommits_info_388_ldest_cons;
    extern constraint default_io_diffCommits_info_388_pdest_cons;
    extern constraint default_io_diffCommits_info_389_ldest_cons;
    extern constraint default_io_diffCommits_info_389_pdest_cons;
    extern constraint default_io_lsq_scommit_cons;
    extern constraint default_io_lsq_pendingMMIOld_cons;
    extern constraint default_io_lsq_pendingst_cons;
    extern constraint default_io_lsq_pendingPtr_flag_cons;
    extern constraint default_io_lsq_pendingPtr_value_cons;
    extern constraint default_io_robDeqPtr_flag_cons;
    extern constraint default_io_robDeqPtr_value_cons;
    extern constraint default_io_csr_fflags_valid_cons;
    extern constraint default_io_csr_fflags_bits_cons;
    extern constraint default_io_csr_vxsat_valid_cons;
    extern constraint default_io_csr_vxsat_bits_cons;
    extern constraint default_io_csr_vstart_valid_cons;
    extern constraint default_io_csr_vstart_bits_cons;
    extern constraint default_io_csr_dirty_fs_cons;
    extern constraint default_io_csr_dirty_vs_cons;
    extern constraint default_io_csr_perfinfo_retiredInstr_cons;
    extern constraint default_io_cpu_halt_cons;
    extern constraint default_io_wfi_wfiReq_cons;
    extern constraint default_io_toDecode_isResumeVType_cons;
    extern constraint default_io_toDecode_walkToArchVType_cons;
    extern constraint default_io_toDecode_walkVType_valid_cons;
    extern constraint default_io_toDecode_walkVType_bits_illegal_cons;
    extern constraint default_io_toDecode_walkVType_bits_vma_cons;
    extern constraint default_io_toDecode_walkVType_bits_vta_cons;
    extern constraint default_io_toDecode_walkVType_bits_vsew_cons;
    extern constraint default_io_toDecode_walkVType_bits_vlmul_cons;
    extern constraint default_io_toDecode_commitVType_vtype_valid_cons;
    extern constraint default_io_toDecode_commitVType_vtype_bits_illegal_cons;
    extern constraint default_io_toDecode_commitVType_vtype_bits_vma_cons;
    extern constraint default_io_toDecode_commitVType_vtype_bits_vta_cons;
    extern constraint default_io_toDecode_commitVType_vtype_bits_vsew_cons;
    extern constraint default_io_toDecode_commitVType_vtype_bits_vlmul_cons;
    extern constraint default_io_toDecode_commitVType_hasVsetvl_cons;
    extern constraint default_io_readGPAMemAddr_valid_cons;
    extern constraint default_io_readGPAMemAddr_bits_ftqPtr_value_cons;
    extern constraint default_io_readGPAMemAddr_bits_ftqOffset_cons;
    extern constraint default_io_toVecExcpMod_logicPhyRegMap_0_valid_cons;
    extern constraint default_io_toVecExcpMod_logicPhyRegMap_0_bits_lreg_cons;
    extern constraint default_io_toVecExcpMod_logicPhyRegMap_0_bits_preg_cons;
    extern constraint default_io_toVecExcpMod_logicPhyRegMap_1_valid_cons;
    extern constraint default_io_toVecExcpMod_logicPhyRegMap_1_bits_lreg_cons;
    extern constraint default_io_toVecExcpMod_logicPhyRegMap_1_bits_preg_cons;
    extern constraint default_io_toVecExcpMod_logicPhyRegMap_2_valid_cons;
    extern constraint default_io_toVecExcpMod_logicPhyRegMap_2_bits_lreg_cons;
    extern constraint default_io_toVecExcpMod_logicPhyRegMap_2_bits_preg_cons;
    extern constraint default_io_toVecExcpMod_logicPhyRegMap_3_valid_cons;
    extern constraint default_io_toVecExcpMod_logicPhyRegMap_3_bits_lreg_cons;
    extern constraint default_io_toVecExcpMod_logicPhyRegMap_3_bits_preg_cons;
    extern constraint default_io_toVecExcpMod_logicPhyRegMap_4_valid_cons;
    extern constraint default_io_toVecExcpMod_logicPhyRegMap_4_bits_lreg_cons;
    extern constraint default_io_toVecExcpMod_logicPhyRegMap_4_bits_preg_cons;
    extern constraint default_io_toVecExcpMod_logicPhyRegMap_5_valid_cons;
    extern constraint default_io_toVecExcpMod_logicPhyRegMap_5_bits_lreg_cons;
    extern constraint default_io_toVecExcpMod_logicPhyRegMap_5_bits_preg_cons;
    extern constraint default_io_toVecExcpMod_excpInfo_valid_cons;
    extern constraint default_io_toVecExcpMod_excpInfo_bits_vstart_cons;
    extern constraint default_io_toVecExcpMod_excpInfo_bits_vsew_cons;
    extern constraint default_io_toVecExcpMod_excpInfo_bits_veew_cons;
    extern constraint default_io_toVecExcpMod_excpInfo_bits_vlmul_cons;
    extern constraint default_io_toVecExcpMod_excpInfo_bits_nf_cons;
    extern constraint default_io_toVecExcpMod_excpInfo_bits_isStride_cons;
    extern constraint default_io_toVecExcpMod_excpInfo_bits_isIndexed_cons;
    extern constraint default_io_toVecExcpMod_excpInfo_bits_isWhole_cons;
    extern constraint default_io_toVecExcpMod_excpInfo_bits_isVlm_cons;
    extern constraint default_io_storeDebugInfo_1_pc_cons;
    extern constraint default_io_perf_0_value_cons;
    extern constraint default_io_perf_1_value_cons;
    extern constraint default_io_perf_2_value_cons;
    extern constraint default_io_perf_3_value_cons;
    extern constraint default_io_perf_4_value_cons;
    extern constraint default_io_perf_5_value_cons;
    extern constraint default_io_perf_6_value_cons;
    extern constraint default_io_perf_7_value_cons;
    extern constraint default_io_perf_8_value_cons;
    extern constraint default_io_perf_9_value_cons;
    extern constraint default_io_perf_10_value_cons;
    extern constraint default_io_perf_11_value_cons;
    extern constraint default_io_perf_12_value_cons;
    extern constraint default_io_perf_13_value_cons;
    extern constraint default_io_perf_14_value_cons;
    extern constraint default_io_perf_15_value_cons;
    extern constraint default_io_perf_16_value_cons;
    extern constraint default_io_perf_17_value_cons;
    extern constraint default_io_error_0_cons;

    extern function new(string name="Rob_output_agent_xaction");
    extern function void pack();
    extern function void unpack();
    extern function void pre_randomize();
    extern function void post_randomize();
    extern function string psdisplay(string prefix = "");
    extern function bit compare(uvm_object rhs, uvm_comparer comparer=null);

    `uvm_object_utils_begin(Rob_output_agent_xaction)
        `uvm_field_int(io_enq_canAccept, UVM_ALL_ON);
        `uvm_field_int(io_enq_canAcceptForDispatch, UVM_ALL_ON);
        `uvm_field_int(io_enq_isEmpty, UVM_ALL_ON);
        `uvm_field_int(io_flushOut_valid, UVM_ALL_ON);
        `uvm_field_int(io_flushOut_bits_isRVC, UVM_ALL_ON);
        `uvm_field_int(io_flushOut_bits_robIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_flushOut_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_flushOut_bits_ftqIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_flushOut_bits_ftqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_flushOut_bits_ftqOffset, UVM_ALL_ON);
        `uvm_field_int(io_flushOut_bits_level, UVM_ALL_ON);
        `uvm_field_int(io_exception_valid, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_instr, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_commitType, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_exceptionVec_0, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_exceptionVec_1, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_exceptionVec_2, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_exceptionVec_3, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_exceptionVec_4, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_exceptionVec_5, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_exceptionVec_6, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_exceptionVec_7, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_exceptionVec_8, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_exceptionVec_9, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_exceptionVec_10, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_exceptionVec_11, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_exceptionVec_12, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_exceptionVec_13, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_exceptionVec_14, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_exceptionVec_15, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_exceptionVec_16, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_exceptionVec_17, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_exceptionVec_18, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_exceptionVec_19, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_exceptionVec_20, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_exceptionVec_21, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_exceptionVec_22, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_exceptionVec_23, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_isPcBkpt, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_isFetchMalAddr, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_gpaddr, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_singleStep, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_crossPageIPFFix, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_isInterrupt, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_isHls, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_trigger, UVM_ALL_ON);
        `uvm_field_int(io_exception_bits_isForVSnonLeafPTE, UVM_ALL_ON);
        `uvm_field_int(io_commits_isCommit, UVM_ALL_ON);
        `uvm_field_int(io_commits_commitValid_0, UVM_ALL_ON);
        `uvm_field_int(io_commits_commitValid_1, UVM_ALL_ON);
        `uvm_field_int(io_commits_commitValid_2, UVM_ALL_ON);
        `uvm_field_int(io_commits_commitValid_3, UVM_ALL_ON);
        `uvm_field_int(io_commits_commitValid_4, UVM_ALL_ON);
        `uvm_field_int(io_commits_commitValid_5, UVM_ALL_ON);
        `uvm_field_int(io_commits_commitValid_6, UVM_ALL_ON);
        `uvm_field_int(io_commits_commitValid_7, UVM_ALL_ON);
        `uvm_field_int(io_commits_isWalk, UVM_ALL_ON);
        `uvm_field_int(io_commits_walkValid_0, UVM_ALL_ON);
        `uvm_field_int(io_commits_walkValid_1, UVM_ALL_ON);
        `uvm_field_int(io_commits_walkValid_2, UVM_ALL_ON);
        `uvm_field_int(io_commits_walkValid_3, UVM_ALL_ON);
        `uvm_field_int(io_commits_walkValid_4, UVM_ALL_ON);
        `uvm_field_int(io_commits_walkValid_5, UVM_ALL_ON);
        `uvm_field_int(io_commits_walkValid_6, UVM_ALL_ON);
        `uvm_field_int(io_commits_walkValid_7, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_walk_v, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_commit_v, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_commit_w, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_realDestSize, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_interrupt_safe, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_wflags, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_fflags, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_vxsat, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_isRVC, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_isVset, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_isHls, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_isVls, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_vls, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_mmio, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_commitType, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_ftqIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_ftqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_ftqOffset, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_instrSize, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_needFlush, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_traceBlockInPipe_itype, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_traceBlockInPipe_iretire, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_traceBlockInPipe_ilastsize, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_debug_pc, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_debug_instr, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_debug_ldest, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_debug_pdest, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_debug_otherPdest_0, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_debug_otherPdest_1, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_debug_otherPdest_2, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_debug_otherPdest_3, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_debug_otherPdest_4, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_debug_otherPdest_5, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_debug_otherPdest_6, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_debug_fuType, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_dirtyFs, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_0_dirtyVs, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_walk_v, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_commit_v, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_commit_w, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_realDestSize, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_interrupt_safe, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_wflags, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_fflags, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_vxsat, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_isRVC, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_isVset, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_isHls, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_isVls, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_vls, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_mmio, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_commitType, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_ftqIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_ftqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_ftqOffset, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_instrSize, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_needFlush, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_traceBlockInPipe_itype, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_traceBlockInPipe_iretire, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_traceBlockInPipe_ilastsize, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_debug_pc, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_debug_instr, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_debug_ldest, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_debug_pdest, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_debug_otherPdest_0, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_debug_otherPdest_1, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_debug_otherPdest_2, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_debug_otherPdest_3, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_debug_otherPdest_4, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_debug_otherPdest_5, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_debug_otherPdest_6, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_debug_fuType, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_dirtyFs, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_1_dirtyVs, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_walk_v, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_commit_v, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_commit_w, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_realDestSize, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_interrupt_safe, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_wflags, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_fflags, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_vxsat, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_isRVC, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_isVset, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_isHls, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_isVls, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_vls, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_mmio, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_commitType, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_ftqIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_ftqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_ftqOffset, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_instrSize, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_needFlush, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_traceBlockInPipe_itype, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_traceBlockInPipe_iretire, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_traceBlockInPipe_ilastsize, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_debug_pc, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_debug_instr, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_debug_ldest, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_debug_pdest, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_debug_otherPdest_0, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_debug_otherPdest_1, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_debug_otherPdest_2, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_debug_otherPdest_3, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_debug_otherPdest_4, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_debug_otherPdest_5, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_debug_otherPdest_6, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_debug_fuType, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_dirtyFs, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_2_dirtyVs, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_walk_v, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_commit_v, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_commit_w, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_realDestSize, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_interrupt_safe, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_wflags, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_fflags, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_vxsat, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_isRVC, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_isVset, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_isHls, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_isVls, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_vls, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_mmio, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_commitType, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_ftqIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_ftqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_ftqOffset, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_instrSize, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_needFlush, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_traceBlockInPipe_itype, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_traceBlockInPipe_iretire, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_traceBlockInPipe_ilastsize, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_debug_pc, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_debug_instr, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_debug_ldest, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_debug_pdest, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_debug_otherPdest_0, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_debug_otherPdest_1, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_debug_otherPdest_2, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_debug_otherPdest_3, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_debug_otherPdest_4, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_debug_otherPdest_5, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_debug_otherPdest_6, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_debug_fuType, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_dirtyFs, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_3_dirtyVs, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_walk_v, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_commit_v, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_commit_w, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_realDestSize, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_interrupt_safe, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_wflags, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_fflags, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_vxsat, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_isRVC, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_isVset, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_isHls, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_isVls, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_vls, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_mmio, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_commitType, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_ftqIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_ftqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_ftqOffset, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_instrSize, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_needFlush, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_traceBlockInPipe_itype, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_traceBlockInPipe_iretire, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_traceBlockInPipe_ilastsize, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_debug_pc, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_debug_instr, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_debug_ldest, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_debug_pdest, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_debug_otherPdest_0, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_debug_otherPdest_1, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_debug_otherPdest_2, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_debug_otherPdest_3, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_debug_otherPdest_4, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_debug_otherPdest_5, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_debug_otherPdest_6, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_debug_fuType, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_dirtyFs, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_4_dirtyVs, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_walk_v, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_commit_v, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_commit_w, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_realDestSize, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_interrupt_safe, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_wflags, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_fflags, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_vxsat, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_isRVC, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_isVset, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_isHls, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_isVls, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_vls, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_mmio, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_commitType, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_ftqIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_ftqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_ftqOffset, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_instrSize, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_needFlush, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_traceBlockInPipe_itype, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_traceBlockInPipe_iretire, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_traceBlockInPipe_ilastsize, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_debug_pc, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_debug_instr, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_debug_ldest, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_debug_pdest, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_debug_otherPdest_0, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_debug_otherPdest_1, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_debug_otherPdest_2, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_debug_otherPdest_3, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_debug_otherPdest_4, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_debug_otherPdest_5, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_debug_otherPdest_6, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_debug_fuType, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_dirtyFs, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_5_dirtyVs, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_walk_v, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_commit_v, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_commit_w, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_realDestSize, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_interrupt_safe, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_wflags, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_fflags, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_vxsat, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_isRVC, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_isVset, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_isHls, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_isVls, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_vls, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_mmio, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_commitType, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_ftqIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_ftqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_ftqOffset, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_instrSize, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_needFlush, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_traceBlockInPipe_itype, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_traceBlockInPipe_iretire, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_traceBlockInPipe_ilastsize, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_debug_pc, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_debug_instr, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_debug_ldest, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_debug_pdest, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_debug_otherPdest_0, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_debug_otherPdest_1, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_debug_otherPdest_2, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_debug_otherPdest_3, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_debug_otherPdest_4, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_debug_otherPdest_5, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_debug_otherPdest_6, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_debug_fuType, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_dirtyFs, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_6_dirtyVs, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_walk_v, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_commit_v, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_commit_w, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_realDestSize, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_interrupt_safe, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_wflags, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_fflags, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_vxsat, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_isRVC, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_isVset, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_isHls, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_isVls, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_vls, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_mmio, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_commitType, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_ftqIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_ftqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_ftqOffset, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_instrSize, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_needFlush, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_traceBlockInPipe_itype, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_traceBlockInPipe_iretire, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_traceBlockInPipe_ilastsize, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_debug_pc, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_debug_instr, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_debug_ldest, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_debug_pdest, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_debug_otherPdest_0, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_debug_otherPdest_1, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_debug_otherPdest_2, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_debug_otherPdest_3, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_debug_otherPdest_4, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_debug_otherPdest_5, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_debug_otherPdest_6, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_debug_fuType, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_dirtyFs, UVM_ALL_ON);
        `uvm_field_int(io_commits_info_7_dirtyVs, UVM_ALL_ON);
        `uvm_field_int(io_commits_robIdx_0_flag, UVM_ALL_ON);
        `uvm_field_int(io_commits_robIdx_0_value, UVM_ALL_ON);
        `uvm_field_int(io_commits_robIdx_1_flag, UVM_ALL_ON);
        `uvm_field_int(io_commits_robIdx_1_value, UVM_ALL_ON);
        `uvm_field_int(io_commits_robIdx_2_flag, UVM_ALL_ON);
        `uvm_field_int(io_commits_robIdx_2_value, UVM_ALL_ON);
        `uvm_field_int(io_commits_robIdx_3_flag, UVM_ALL_ON);
        `uvm_field_int(io_commits_robIdx_3_value, UVM_ALL_ON);
        `uvm_field_int(io_commits_robIdx_4_flag, UVM_ALL_ON);
        `uvm_field_int(io_commits_robIdx_4_value, UVM_ALL_ON);
        `uvm_field_int(io_commits_robIdx_5_flag, UVM_ALL_ON);
        `uvm_field_int(io_commits_robIdx_5_value, UVM_ALL_ON);
        `uvm_field_int(io_commits_robIdx_6_flag, UVM_ALL_ON);
        `uvm_field_int(io_commits_robIdx_6_value, UVM_ALL_ON);
        `uvm_field_int(io_commits_robIdx_7_flag, UVM_ALL_ON);
        `uvm_field_int(io_commits_robIdx_7_value, UVM_ALL_ON);
        `uvm_field_int(io_trace_blockCommit, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_0_valid, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_0_bits_ftqOffset, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_1_valid, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_1_bits_ftqOffset, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_2_valid, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_2_bits_ftqOffset, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_3_valid, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_3_bits_ftqOffset, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_4_valid, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_4_bits_ftqOffset, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_5_valid, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_5_bits_ftqOffset, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_6_valid, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_6_bits_ftqOffset, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_7_valid, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_7_bits_ftqOffset, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire, UVM_ALL_ON);
        `uvm_field_int(io_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_isCommit, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_commitValid_0, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_commitValid_1, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_commitValid_2, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_commitValid_3, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_commitValid_4, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_commitValid_5, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_isWalk, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_walkValid_0, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_walkValid_1, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_walkValid_2, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_walkValid_3, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_walkValid_4, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_walkValid_5, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_0_ldest, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_0_pdest, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_0_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_0_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_0_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_0_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_0_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_0_isMove, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_1_ldest, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_1_pdest, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_1_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_1_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_1_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_1_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_1_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_1_isMove, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_2_ldest, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_2_pdest, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_2_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_2_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_2_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_2_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_2_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_2_isMove, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_3_ldest, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_3_pdest, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_3_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_3_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_3_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_3_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_3_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_3_isMove, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_4_ldest, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_4_pdest, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_4_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_4_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_4_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_4_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_4_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_4_isMove, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_5_ldest, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_5_pdest, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_5_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_5_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_5_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_5_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_5_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_rabCommits_info_5_isMove, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_0, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_1, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_2, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_3, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_4, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_5, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_6, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_7, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_8, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_9, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_10, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_11, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_12, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_13, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_14, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_15, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_16, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_17, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_18, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_19, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_20, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_21, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_22, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_23, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_24, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_25, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_26, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_27, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_28, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_29, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_30, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_31, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_32, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_33, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_34, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_35, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_36, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_37, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_38, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_39, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_40, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_41, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_42, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_43, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_44, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_45, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_46, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_47, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_48, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_49, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_50, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_51, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_52, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_53, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_54, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_55, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_56, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_57, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_58, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_59, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_60, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_61, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_62, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_63, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_64, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_65, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_66, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_67, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_68, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_69, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_70, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_71, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_72, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_73, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_74, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_75, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_76, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_77, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_78, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_79, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_80, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_81, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_82, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_83, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_84, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_85, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_86, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_87, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_88, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_89, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_90, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_91, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_92, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_93, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_94, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_95, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_96, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_97, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_98, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_99, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_100, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_101, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_102, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_103, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_104, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_105, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_106, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_107, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_108, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_109, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_110, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_111, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_112, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_113, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_114, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_115, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_116, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_117, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_118, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_119, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_120, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_121, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_122, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_123, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_124, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_125, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_126, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_127, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_128, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_129, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_130, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_131, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_132, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_133, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_134, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_135, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_136, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_137, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_138, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_139, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_140, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_141, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_142, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_143, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_144, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_145, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_146, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_147, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_148, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_149, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_150, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_151, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_152, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_153, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_154, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_155, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_156, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_157, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_158, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_159, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_160, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_161, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_162, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_163, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_164, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_165, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_166, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_167, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_168, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_169, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_170, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_171, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_172, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_173, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_174, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_175, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_176, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_177, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_178, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_179, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_180, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_181, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_182, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_183, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_184, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_185, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_186, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_187, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_188, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_189, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_190, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_191, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_192, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_193, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_194, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_195, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_196, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_197, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_198, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_199, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_200, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_201, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_202, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_203, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_204, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_205, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_206, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_207, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_208, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_209, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_210, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_211, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_212, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_213, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_214, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_215, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_216, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_217, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_218, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_219, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_220, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_221, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_222, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_223, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_224, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_225, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_226, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_227, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_228, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_229, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_230, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_231, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_232, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_233, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_234, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_235, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_236, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_237, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_238, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_239, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_240, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_241, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_242, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_243, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_244, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_245, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_246, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_247, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_248, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_249, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_250, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_251, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_252, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_253, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_commitValid_254, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_0_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_0_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_0_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_0_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_0_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_0_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_0_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_1_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_1_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_1_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_1_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_1_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_1_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_1_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_2_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_2_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_2_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_2_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_2_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_2_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_2_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_3_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_3_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_3_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_3_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_3_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_3_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_3_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_4_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_4_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_4_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_4_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_4_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_4_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_4_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_5_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_5_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_5_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_5_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_5_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_5_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_5_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_6_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_6_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_6_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_6_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_6_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_6_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_6_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_7_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_7_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_7_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_7_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_7_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_7_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_7_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_8_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_8_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_8_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_8_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_8_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_8_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_8_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_9_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_9_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_9_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_9_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_9_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_9_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_9_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_10_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_10_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_10_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_10_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_10_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_10_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_10_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_11_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_11_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_11_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_11_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_11_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_11_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_11_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_12_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_12_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_12_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_12_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_12_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_12_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_12_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_13_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_13_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_13_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_13_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_13_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_13_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_13_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_14_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_14_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_14_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_14_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_14_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_14_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_14_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_15_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_15_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_15_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_15_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_15_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_15_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_15_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_16_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_16_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_16_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_16_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_16_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_16_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_16_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_17_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_17_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_17_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_17_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_17_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_17_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_17_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_18_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_18_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_18_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_18_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_18_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_18_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_18_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_19_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_19_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_19_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_19_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_19_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_19_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_19_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_20_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_20_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_20_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_20_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_20_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_20_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_20_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_21_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_21_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_21_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_21_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_21_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_21_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_21_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_22_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_22_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_22_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_22_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_22_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_22_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_22_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_23_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_23_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_23_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_23_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_23_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_23_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_23_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_24_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_24_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_24_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_24_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_24_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_24_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_24_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_25_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_25_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_25_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_25_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_25_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_25_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_25_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_26_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_26_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_26_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_26_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_26_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_26_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_26_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_27_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_27_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_27_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_27_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_27_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_27_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_27_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_28_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_28_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_28_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_28_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_28_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_28_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_28_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_29_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_29_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_29_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_29_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_29_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_29_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_29_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_30_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_30_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_30_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_30_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_30_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_30_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_30_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_31_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_31_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_31_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_31_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_31_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_31_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_31_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_32_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_32_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_32_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_32_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_32_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_32_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_32_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_33_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_33_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_33_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_33_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_33_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_33_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_33_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_34_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_34_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_34_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_34_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_34_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_34_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_34_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_35_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_35_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_35_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_35_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_35_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_35_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_35_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_36_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_36_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_36_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_36_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_36_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_36_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_36_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_37_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_37_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_37_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_37_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_37_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_37_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_37_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_38_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_38_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_38_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_38_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_38_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_38_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_38_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_39_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_39_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_39_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_39_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_39_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_39_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_39_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_40_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_40_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_40_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_40_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_40_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_40_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_40_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_41_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_41_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_41_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_41_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_41_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_41_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_41_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_42_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_42_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_42_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_42_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_42_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_42_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_42_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_43_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_43_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_43_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_43_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_43_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_43_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_43_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_44_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_44_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_44_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_44_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_44_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_44_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_44_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_45_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_45_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_45_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_45_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_45_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_45_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_45_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_46_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_46_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_46_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_46_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_46_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_46_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_46_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_47_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_47_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_47_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_47_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_47_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_47_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_47_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_48_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_48_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_48_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_48_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_48_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_48_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_48_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_49_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_49_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_49_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_49_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_49_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_49_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_49_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_50_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_50_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_50_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_50_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_50_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_50_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_50_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_51_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_51_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_51_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_51_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_51_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_51_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_51_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_52_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_52_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_52_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_52_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_52_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_52_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_52_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_53_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_53_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_53_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_53_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_53_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_53_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_53_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_54_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_54_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_54_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_54_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_54_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_54_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_54_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_55_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_55_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_55_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_55_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_55_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_55_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_55_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_56_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_56_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_56_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_56_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_56_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_56_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_56_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_57_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_57_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_57_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_57_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_57_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_57_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_57_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_58_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_58_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_58_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_58_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_58_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_58_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_58_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_59_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_59_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_59_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_59_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_59_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_59_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_59_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_60_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_60_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_60_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_60_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_60_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_60_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_60_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_61_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_61_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_61_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_61_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_61_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_61_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_61_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_62_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_62_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_62_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_62_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_62_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_62_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_62_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_63_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_63_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_63_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_63_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_63_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_63_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_63_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_64_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_64_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_64_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_64_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_64_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_64_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_64_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_65_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_65_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_65_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_65_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_65_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_65_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_65_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_66_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_66_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_66_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_66_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_66_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_66_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_66_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_67_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_67_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_67_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_67_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_67_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_67_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_67_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_68_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_68_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_68_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_68_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_68_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_68_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_68_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_69_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_69_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_69_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_69_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_69_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_69_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_69_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_70_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_70_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_70_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_70_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_70_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_70_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_70_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_71_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_71_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_71_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_71_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_71_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_71_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_71_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_72_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_72_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_72_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_72_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_72_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_72_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_72_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_73_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_73_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_73_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_73_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_73_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_73_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_73_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_74_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_74_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_74_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_74_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_74_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_74_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_74_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_75_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_75_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_75_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_75_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_75_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_75_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_75_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_76_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_76_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_76_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_76_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_76_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_76_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_76_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_77_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_77_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_77_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_77_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_77_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_77_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_77_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_78_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_78_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_78_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_78_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_78_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_78_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_78_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_79_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_79_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_79_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_79_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_79_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_79_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_79_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_80_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_80_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_80_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_80_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_80_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_80_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_80_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_81_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_81_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_81_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_81_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_81_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_81_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_81_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_82_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_82_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_82_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_82_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_82_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_82_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_82_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_83_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_83_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_83_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_83_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_83_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_83_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_83_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_84_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_84_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_84_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_84_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_84_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_84_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_84_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_85_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_85_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_85_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_85_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_85_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_85_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_85_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_86_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_86_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_86_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_86_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_86_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_86_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_86_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_87_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_87_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_87_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_87_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_87_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_87_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_87_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_88_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_88_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_88_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_88_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_88_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_88_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_88_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_89_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_89_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_89_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_89_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_89_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_89_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_89_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_90_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_90_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_90_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_90_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_90_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_90_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_90_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_91_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_91_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_91_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_91_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_91_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_91_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_91_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_92_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_92_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_92_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_92_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_92_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_92_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_92_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_93_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_93_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_93_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_93_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_93_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_93_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_93_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_94_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_94_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_94_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_94_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_94_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_94_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_94_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_95_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_95_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_95_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_95_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_95_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_95_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_95_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_96_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_96_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_96_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_96_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_96_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_96_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_96_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_97_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_97_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_97_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_97_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_97_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_97_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_97_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_98_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_98_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_98_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_98_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_98_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_98_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_98_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_99_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_99_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_99_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_99_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_99_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_99_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_99_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_100_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_100_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_100_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_100_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_100_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_100_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_100_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_101_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_101_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_101_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_101_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_101_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_101_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_101_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_102_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_102_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_102_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_102_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_102_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_102_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_102_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_103_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_103_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_103_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_103_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_103_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_103_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_103_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_104_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_104_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_104_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_104_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_104_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_104_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_104_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_105_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_105_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_105_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_105_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_105_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_105_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_105_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_106_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_106_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_106_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_106_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_106_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_106_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_106_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_107_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_107_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_107_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_107_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_107_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_107_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_107_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_108_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_108_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_108_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_108_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_108_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_108_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_108_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_109_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_109_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_109_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_109_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_109_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_109_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_109_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_110_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_110_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_110_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_110_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_110_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_110_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_110_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_111_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_111_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_111_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_111_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_111_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_111_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_111_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_112_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_112_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_112_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_112_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_112_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_112_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_112_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_113_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_113_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_113_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_113_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_113_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_113_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_113_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_114_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_114_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_114_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_114_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_114_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_114_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_114_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_115_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_115_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_115_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_115_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_115_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_115_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_115_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_116_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_116_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_116_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_116_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_116_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_116_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_116_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_117_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_117_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_117_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_117_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_117_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_117_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_117_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_118_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_118_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_118_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_118_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_118_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_118_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_118_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_119_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_119_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_119_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_119_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_119_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_119_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_119_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_120_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_120_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_120_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_120_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_120_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_120_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_120_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_121_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_121_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_121_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_121_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_121_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_121_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_121_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_122_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_122_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_122_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_122_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_122_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_122_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_122_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_123_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_123_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_123_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_123_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_123_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_123_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_123_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_124_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_124_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_124_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_124_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_124_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_124_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_124_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_125_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_125_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_125_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_125_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_125_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_125_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_125_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_126_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_126_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_126_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_126_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_126_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_126_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_126_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_127_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_127_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_127_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_127_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_127_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_127_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_127_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_128_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_128_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_128_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_128_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_128_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_128_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_128_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_129_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_129_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_129_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_129_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_129_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_129_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_129_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_130_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_130_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_130_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_130_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_130_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_130_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_130_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_131_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_131_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_131_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_131_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_131_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_131_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_131_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_132_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_132_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_132_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_132_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_132_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_132_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_132_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_133_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_133_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_133_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_133_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_133_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_133_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_133_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_134_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_134_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_134_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_134_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_134_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_134_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_134_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_135_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_135_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_135_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_135_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_135_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_135_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_135_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_136_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_136_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_136_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_136_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_136_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_136_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_136_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_137_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_137_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_137_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_137_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_137_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_137_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_137_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_138_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_138_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_138_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_138_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_138_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_138_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_138_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_139_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_139_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_139_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_139_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_139_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_139_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_139_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_140_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_140_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_140_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_140_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_140_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_140_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_140_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_141_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_141_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_141_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_141_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_141_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_141_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_141_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_142_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_142_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_142_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_142_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_142_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_142_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_142_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_143_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_143_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_143_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_143_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_143_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_143_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_143_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_144_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_144_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_144_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_144_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_144_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_144_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_144_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_145_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_145_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_145_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_145_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_145_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_145_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_145_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_146_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_146_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_146_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_146_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_146_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_146_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_146_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_147_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_147_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_147_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_147_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_147_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_147_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_147_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_148_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_148_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_148_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_148_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_148_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_148_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_148_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_149_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_149_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_149_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_149_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_149_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_149_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_149_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_150_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_150_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_150_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_150_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_150_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_150_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_150_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_151_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_151_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_151_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_151_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_151_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_151_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_151_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_152_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_152_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_152_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_152_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_152_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_152_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_152_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_153_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_153_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_153_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_153_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_153_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_153_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_153_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_154_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_154_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_154_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_154_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_154_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_154_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_154_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_155_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_155_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_155_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_155_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_155_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_155_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_155_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_156_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_156_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_156_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_156_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_156_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_156_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_156_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_157_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_157_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_157_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_157_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_157_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_157_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_157_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_158_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_158_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_158_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_158_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_158_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_158_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_158_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_159_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_159_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_159_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_159_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_159_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_159_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_159_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_160_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_160_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_160_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_160_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_160_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_160_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_160_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_161_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_161_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_161_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_161_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_161_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_161_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_161_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_162_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_162_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_162_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_162_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_162_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_162_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_162_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_163_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_163_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_163_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_163_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_163_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_163_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_163_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_164_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_164_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_164_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_164_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_164_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_164_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_164_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_165_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_165_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_165_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_165_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_165_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_165_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_165_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_166_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_166_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_166_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_166_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_166_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_166_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_166_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_167_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_167_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_167_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_167_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_167_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_167_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_167_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_168_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_168_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_168_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_168_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_168_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_168_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_168_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_169_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_169_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_169_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_169_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_169_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_169_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_169_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_170_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_170_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_170_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_170_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_170_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_170_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_170_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_171_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_171_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_171_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_171_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_171_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_171_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_171_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_172_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_172_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_172_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_172_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_172_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_172_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_172_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_173_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_173_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_173_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_173_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_173_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_173_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_173_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_174_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_174_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_174_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_174_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_174_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_174_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_174_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_175_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_175_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_175_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_175_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_175_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_175_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_175_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_176_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_176_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_176_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_176_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_176_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_176_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_176_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_177_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_177_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_177_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_177_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_177_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_177_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_177_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_178_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_178_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_178_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_178_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_178_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_178_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_178_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_179_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_179_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_179_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_179_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_179_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_179_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_179_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_180_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_180_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_180_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_180_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_180_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_180_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_180_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_181_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_181_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_181_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_181_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_181_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_181_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_181_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_182_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_182_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_182_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_182_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_182_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_182_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_182_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_183_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_183_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_183_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_183_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_183_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_183_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_183_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_184_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_184_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_184_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_184_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_184_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_184_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_184_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_185_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_185_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_185_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_185_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_185_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_185_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_185_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_186_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_186_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_186_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_186_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_186_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_186_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_186_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_187_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_187_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_187_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_187_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_187_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_187_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_187_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_188_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_188_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_188_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_188_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_188_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_188_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_188_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_189_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_189_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_189_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_189_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_189_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_189_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_189_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_190_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_190_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_190_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_190_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_190_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_190_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_190_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_191_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_191_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_191_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_191_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_191_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_191_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_191_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_192_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_192_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_192_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_192_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_192_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_192_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_192_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_193_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_193_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_193_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_193_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_193_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_193_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_193_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_194_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_194_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_194_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_194_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_194_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_194_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_194_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_195_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_195_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_195_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_195_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_195_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_195_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_195_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_196_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_196_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_196_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_196_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_196_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_196_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_196_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_197_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_197_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_197_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_197_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_197_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_197_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_197_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_198_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_198_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_198_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_198_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_198_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_198_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_198_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_199_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_199_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_199_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_199_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_199_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_199_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_199_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_200_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_200_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_200_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_200_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_200_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_200_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_200_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_201_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_201_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_201_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_201_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_201_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_201_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_201_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_202_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_202_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_202_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_202_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_202_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_202_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_202_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_203_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_203_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_203_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_203_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_203_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_203_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_203_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_204_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_204_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_204_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_204_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_204_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_204_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_204_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_205_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_205_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_205_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_205_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_205_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_205_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_205_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_206_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_206_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_206_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_206_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_206_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_206_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_206_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_207_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_207_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_207_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_207_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_207_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_207_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_207_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_208_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_208_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_208_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_208_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_208_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_208_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_208_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_209_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_209_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_209_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_209_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_209_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_209_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_209_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_210_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_210_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_210_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_210_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_210_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_210_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_210_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_211_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_211_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_211_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_211_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_211_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_211_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_211_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_212_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_212_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_212_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_212_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_212_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_212_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_212_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_213_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_213_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_213_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_213_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_213_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_213_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_213_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_214_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_214_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_214_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_214_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_214_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_214_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_214_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_215_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_215_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_215_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_215_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_215_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_215_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_215_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_216_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_216_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_216_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_216_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_216_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_216_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_216_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_217_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_217_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_217_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_217_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_217_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_217_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_217_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_218_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_218_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_218_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_218_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_218_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_218_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_218_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_219_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_219_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_219_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_219_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_219_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_219_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_219_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_220_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_220_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_220_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_220_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_220_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_220_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_220_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_221_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_221_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_221_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_221_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_221_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_221_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_221_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_222_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_222_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_222_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_222_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_222_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_222_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_222_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_223_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_223_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_223_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_223_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_223_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_223_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_223_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_224_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_224_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_224_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_224_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_224_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_224_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_224_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_225_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_225_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_225_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_225_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_225_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_225_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_225_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_226_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_226_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_226_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_226_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_226_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_226_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_226_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_227_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_227_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_227_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_227_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_227_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_227_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_227_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_228_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_228_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_228_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_228_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_228_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_228_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_228_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_229_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_229_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_229_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_229_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_229_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_229_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_229_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_230_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_230_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_230_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_230_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_230_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_230_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_230_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_231_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_231_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_231_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_231_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_231_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_231_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_231_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_232_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_232_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_232_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_232_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_232_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_232_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_232_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_233_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_233_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_233_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_233_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_233_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_233_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_233_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_234_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_234_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_234_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_234_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_234_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_234_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_234_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_235_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_235_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_235_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_235_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_235_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_235_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_235_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_236_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_236_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_236_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_236_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_236_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_236_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_236_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_237_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_237_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_237_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_237_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_237_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_237_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_237_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_238_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_238_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_238_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_238_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_238_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_238_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_238_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_239_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_239_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_239_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_239_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_239_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_239_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_239_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_240_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_240_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_240_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_240_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_240_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_240_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_240_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_241_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_241_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_241_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_241_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_241_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_241_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_241_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_242_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_242_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_242_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_242_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_242_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_242_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_242_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_243_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_243_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_243_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_243_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_243_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_243_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_243_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_244_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_244_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_244_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_244_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_244_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_244_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_244_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_245_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_245_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_245_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_245_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_245_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_245_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_245_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_246_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_246_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_246_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_246_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_246_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_246_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_246_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_247_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_247_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_247_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_247_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_247_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_247_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_247_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_248_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_248_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_248_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_248_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_248_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_248_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_248_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_249_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_249_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_249_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_249_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_249_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_249_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_249_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_250_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_250_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_250_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_250_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_250_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_250_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_250_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_251_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_251_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_251_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_251_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_251_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_251_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_251_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_252_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_252_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_252_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_252_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_252_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_252_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_252_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_253_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_253_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_253_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_253_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_253_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_253_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_253_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_254_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_254_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_254_rfWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_254_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_254_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_254_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_254_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_255_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_255_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_256_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_256_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_257_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_257_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_258_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_258_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_259_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_259_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_260_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_260_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_261_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_261_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_262_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_262_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_263_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_263_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_264_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_264_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_265_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_265_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_266_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_266_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_267_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_267_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_268_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_268_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_269_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_269_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_270_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_270_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_271_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_271_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_272_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_272_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_273_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_273_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_274_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_274_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_275_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_275_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_276_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_276_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_277_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_277_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_278_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_278_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_279_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_279_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_280_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_280_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_281_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_281_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_282_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_282_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_283_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_283_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_284_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_284_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_285_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_285_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_286_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_286_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_287_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_287_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_288_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_288_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_289_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_289_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_290_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_290_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_291_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_291_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_292_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_292_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_293_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_293_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_294_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_294_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_295_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_295_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_296_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_296_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_297_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_297_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_298_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_298_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_299_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_299_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_300_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_300_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_301_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_301_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_302_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_302_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_303_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_303_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_304_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_304_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_305_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_305_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_306_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_306_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_307_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_307_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_308_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_308_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_309_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_309_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_310_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_310_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_311_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_311_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_312_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_312_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_313_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_313_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_314_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_314_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_315_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_315_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_316_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_316_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_317_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_317_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_318_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_318_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_319_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_319_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_320_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_320_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_321_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_321_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_322_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_322_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_323_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_323_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_324_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_324_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_325_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_325_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_326_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_326_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_327_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_327_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_328_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_328_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_329_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_329_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_330_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_330_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_331_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_331_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_332_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_332_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_333_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_333_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_334_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_334_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_335_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_335_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_336_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_336_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_337_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_337_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_338_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_338_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_339_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_339_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_340_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_340_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_341_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_341_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_342_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_342_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_343_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_343_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_344_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_344_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_345_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_345_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_346_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_346_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_347_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_347_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_348_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_348_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_349_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_349_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_350_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_350_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_351_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_351_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_352_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_352_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_353_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_353_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_354_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_354_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_355_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_355_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_356_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_356_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_357_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_357_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_358_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_358_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_359_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_359_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_360_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_360_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_361_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_361_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_362_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_362_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_363_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_363_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_364_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_364_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_365_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_365_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_366_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_366_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_367_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_367_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_368_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_368_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_369_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_369_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_370_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_370_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_371_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_371_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_372_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_372_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_373_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_373_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_374_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_374_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_375_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_375_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_376_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_376_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_377_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_377_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_378_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_378_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_379_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_379_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_380_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_380_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_381_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_381_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_382_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_382_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_383_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_383_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_384_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_384_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_385_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_385_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_386_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_386_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_387_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_387_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_388_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_388_pdest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_389_ldest, UVM_ALL_ON);
        `uvm_field_int(io_diffCommits_info_389_pdest, UVM_ALL_ON);
        `uvm_field_int(io_lsq_scommit, UVM_ALL_ON);
        `uvm_field_int(io_lsq_pendingMMIOld, UVM_ALL_ON);
        `uvm_field_int(io_lsq_pendingst, UVM_ALL_ON);
        `uvm_field_int(io_lsq_pendingPtr_flag, UVM_ALL_ON);
        `uvm_field_int(io_lsq_pendingPtr_value, UVM_ALL_ON);
        `uvm_field_int(io_robDeqPtr_flag, UVM_ALL_ON);
        `uvm_field_int(io_robDeqPtr_value, UVM_ALL_ON);
        `uvm_field_int(io_csr_fflags_valid, UVM_ALL_ON);
        `uvm_field_int(io_csr_fflags_bits, UVM_ALL_ON);
        `uvm_field_int(io_csr_vxsat_valid, UVM_ALL_ON);
        `uvm_field_int(io_csr_vxsat_bits, UVM_ALL_ON);
        `uvm_field_int(io_csr_vstart_valid, UVM_ALL_ON);
        `uvm_field_int(io_csr_vstart_bits, UVM_ALL_ON);
        `uvm_field_int(io_csr_dirty_fs, UVM_ALL_ON);
        `uvm_field_int(io_csr_dirty_vs, UVM_ALL_ON);
        `uvm_field_int(io_csr_perfinfo_retiredInstr, UVM_ALL_ON);
        `uvm_field_int(io_cpu_halt, UVM_ALL_ON);
        `uvm_field_int(io_wfi_wfiReq, UVM_ALL_ON);
        `uvm_field_int(io_toDecode_isResumeVType, UVM_ALL_ON);
        `uvm_field_int(io_toDecode_walkToArchVType, UVM_ALL_ON);
        `uvm_field_int(io_toDecode_walkVType_valid, UVM_ALL_ON);
        `uvm_field_int(io_toDecode_walkVType_bits_illegal, UVM_ALL_ON);
        `uvm_field_int(io_toDecode_walkVType_bits_vma, UVM_ALL_ON);
        `uvm_field_int(io_toDecode_walkVType_bits_vta, UVM_ALL_ON);
        `uvm_field_int(io_toDecode_walkVType_bits_vsew, UVM_ALL_ON);
        `uvm_field_int(io_toDecode_walkVType_bits_vlmul, UVM_ALL_ON);
        `uvm_field_int(io_toDecode_commitVType_vtype_valid, UVM_ALL_ON);
        `uvm_field_int(io_toDecode_commitVType_vtype_bits_illegal, UVM_ALL_ON);
        `uvm_field_int(io_toDecode_commitVType_vtype_bits_vma, UVM_ALL_ON);
        `uvm_field_int(io_toDecode_commitVType_vtype_bits_vta, UVM_ALL_ON);
        `uvm_field_int(io_toDecode_commitVType_vtype_bits_vsew, UVM_ALL_ON);
        `uvm_field_int(io_toDecode_commitVType_vtype_bits_vlmul, UVM_ALL_ON);
        `uvm_field_int(io_toDecode_commitVType_hasVsetvl, UVM_ALL_ON);
        `uvm_field_int(io_readGPAMemAddr_valid, UVM_ALL_ON);
        `uvm_field_int(io_readGPAMemAddr_bits_ftqPtr_value, UVM_ALL_ON);
        `uvm_field_int(io_readGPAMemAddr_bits_ftqOffset, UVM_ALL_ON);
        `uvm_field_int(io_toVecExcpMod_logicPhyRegMap_0_valid, UVM_ALL_ON);
        `uvm_field_int(io_toVecExcpMod_logicPhyRegMap_0_bits_lreg, UVM_ALL_ON);
        `uvm_field_int(io_toVecExcpMod_logicPhyRegMap_0_bits_preg, UVM_ALL_ON);
        `uvm_field_int(io_toVecExcpMod_logicPhyRegMap_1_valid, UVM_ALL_ON);
        `uvm_field_int(io_toVecExcpMod_logicPhyRegMap_1_bits_lreg, UVM_ALL_ON);
        `uvm_field_int(io_toVecExcpMod_logicPhyRegMap_1_bits_preg, UVM_ALL_ON);
        `uvm_field_int(io_toVecExcpMod_logicPhyRegMap_2_valid, UVM_ALL_ON);
        `uvm_field_int(io_toVecExcpMod_logicPhyRegMap_2_bits_lreg, UVM_ALL_ON);
        `uvm_field_int(io_toVecExcpMod_logicPhyRegMap_2_bits_preg, UVM_ALL_ON);
        `uvm_field_int(io_toVecExcpMod_logicPhyRegMap_3_valid, UVM_ALL_ON);
        `uvm_field_int(io_toVecExcpMod_logicPhyRegMap_3_bits_lreg, UVM_ALL_ON);
        `uvm_field_int(io_toVecExcpMod_logicPhyRegMap_3_bits_preg, UVM_ALL_ON);
        `uvm_field_int(io_toVecExcpMod_logicPhyRegMap_4_valid, UVM_ALL_ON);
        `uvm_field_int(io_toVecExcpMod_logicPhyRegMap_4_bits_lreg, UVM_ALL_ON);
        `uvm_field_int(io_toVecExcpMod_logicPhyRegMap_4_bits_preg, UVM_ALL_ON);
        `uvm_field_int(io_toVecExcpMod_logicPhyRegMap_5_valid, UVM_ALL_ON);
        `uvm_field_int(io_toVecExcpMod_logicPhyRegMap_5_bits_lreg, UVM_ALL_ON);
        `uvm_field_int(io_toVecExcpMod_logicPhyRegMap_5_bits_preg, UVM_ALL_ON);
        `uvm_field_int(io_toVecExcpMod_excpInfo_valid, UVM_ALL_ON);
        `uvm_field_int(io_toVecExcpMod_excpInfo_bits_vstart, UVM_ALL_ON);
        `uvm_field_int(io_toVecExcpMod_excpInfo_bits_vsew, UVM_ALL_ON);
        `uvm_field_int(io_toVecExcpMod_excpInfo_bits_veew, UVM_ALL_ON);
        `uvm_field_int(io_toVecExcpMod_excpInfo_bits_vlmul, UVM_ALL_ON);
        `uvm_field_int(io_toVecExcpMod_excpInfo_bits_nf, UVM_ALL_ON);
        `uvm_field_int(io_toVecExcpMod_excpInfo_bits_isStride, UVM_ALL_ON);
        `uvm_field_int(io_toVecExcpMod_excpInfo_bits_isIndexed, UVM_ALL_ON);
        `uvm_field_int(io_toVecExcpMod_excpInfo_bits_isWhole, UVM_ALL_ON);
        `uvm_field_int(io_toVecExcpMod_excpInfo_bits_isVlm, UVM_ALL_ON);
        `uvm_field_int(io_storeDebugInfo_1_pc, UVM_ALL_ON);
        `uvm_field_int(io_perf_0_value, UVM_ALL_ON);
        `uvm_field_int(io_perf_1_value, UVM_ALL_ON);
        `uvm_field_int(io_perf_2_value, UVM_ALL_ON);
        `uvm_field_int(io_perf_3_value, UVM_ALL_ON);
        `uvm_field_int(io_perf_4_value, UVM_ALL_ON);
        `uvm_field_int(io_perf_5_value, UVM_ALL_ON);
        `uvm_field_int(io_perf_6_value, UVM_ALL_ON);
        `uvm_field_int(io_perf_7_value, UVM_ALL_ON);
        `uvm_field_int(io_perf_8_value, UVM_ALL_ON);
        `uvm_field_int(io_perf_9_value, UVM_ALL_ON);
        `uvm_field_int(io_perf_10_value, UVM_ALL_ON);
        `uvm_field_int(io_perf_11_value, UVM_ALL_ON);
        `uvm_field_int(io_perf_12_value, UVM_ALL_ON);
        `uvm_field_int(io_perf_13_value, UVM_ALL_ON);
        `uvm_field_int(io_perf_14_value, UVM_ALL_ON);
        `uvm_field_int(io_perf_15_value, UVM_ALL_ON);
        `uvm_field_int(io_perf_16_value, UVM_ALL_ON);
        `uvm_field_int(io_perf_17_value, UVM_ALL_ON);
        `uvm_field_int(io_error_0, UVM_ALL_ON);

    `uvm_object_utils_end

endclass:Rob_output_agent_xaction

constraint Rob_output_agent_xaction::default_io_enq_canAccept_cons{

}

constraint Rob_output_agent_xaction::default_io_enq_canAcceptForDispatch_cons{

}

constraint Rob_output_agent_xaction::default_io_enq_isEmpty_cons{

}

constraint Rob_output_agent_xaction::default_io_flushOut_valid_cons{

}

constraint Rob_output_agent_xaction::default_io_flushOut_bits_isRVC_cons{

}

constraint Rob_output_agent_xaction::default_io_flushOut_bits_robIdx_flag_cons{

}

constraint Rob_output_agent_xaction::default_io_flushOut_bits_robIdx_value_cons{

}

constraint Rob_output_agent_xaction::default_io_flushOut_bits_ftqIdx_flag_cons{

}

constraint Rob_output_agent_xaction::default_io_flushOut_bits_ftqIdx_value_cons{

}

constraint Rob_output_agent_xaction::default_io_flushOut_bits_ftqOffset_cons{

}

constraint Rob_output_agent_xaction::default_io_flushOut_bits_level_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_valid_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_instr_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_commitType_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_exceptionVec_0_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_exceptionVec_1_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_exceptionVec_2_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_exceptionVec_3_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_exceptionVec_4_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_exceptionVec_5_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_exceptionVec_6_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_exceptionVec_7_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_exceptionVec_8_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_exceptionVec_9_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_exceptionVec_10_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_exceptionVec_11_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_exceptionVec_12_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_exceptionVec_13_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_exceptionVec_14_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_exceptionVec_15_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_exceptionVec_16_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_exceptionVec_17_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_exceptionVec_18_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_exceptionVec_19_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_exceptionVec_20_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_exceptionVec_21_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_exceptionVec_22_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_exceptionVec_23_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_isPcBkpt_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_isFetchMalAddr_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_gpaddr_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_singleStep_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_crossPageIPFFix_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_isInterrupt_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_isHls_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_trigger_cons{

}

constraint Rob_output_agent_xaction::default_io_exception_bits_isForVSnonLeafPTE_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_isCommit_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_commitValid_0_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_commitValid_1_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_commitValid_2_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_commitValid_3_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_commitValid_4_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_commitValid_5_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_commitValid_6_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_commitValid_7_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_isWalk_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_walkValid_0_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_walkValid_1_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_walkValid_2_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_walkValid_3_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_walkValid_4_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_walkValid_5_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_walkValid_6_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_walkValid_7_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_walk_v_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_commit_v_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_commit_w_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_realDestSize_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_interrupt_safe_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_wflags_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_fflags_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_vxsat_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_isRVC_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_isVset_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_isHls_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_isVls_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_vls_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_mmio_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_commitType_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_ftqIdx_flag_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_ftqIdx_value_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_ftqOffset_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_instrSize_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_needFlush_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_traceBlockInPipe_itype_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_traceBlockInPipe_iretire_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_traceBlockInPipe_ilastsize_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_debug_pc_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_debug_instr_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_debug_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_debug_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_debug_otherPdest_0_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_debug_otherPdest_1_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_debug_otherPdest_2_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_debug_otherPdest_3_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_debug_otherPdest_4_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_debug_otherPdest_5_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_debug_otherPdest_6_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_debug_fuType_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_dirtyFs_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_0_dirtyVs_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_walk_v_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_commit_v_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_commit_w_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_realDestSize_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_interrupt_safe_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_wflags_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_fflags_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_vxsat_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_isRVC_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_isVset_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_isHls_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_isVls_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_vls_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_mmio_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_commitType_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_ftqIdx_flag_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_ftqIdx_value_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_ftqOffset_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_instrSize_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_needFlush_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_traceBlockInPipe_itype_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_traceBlockInPipe_iretire_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_traceBlockInPipe_ilastsize_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_debug_pc_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_debug_instr_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_debug_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_debug_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_debug_otherPdest_0_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_debug_otherPdest_1_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_debug_otherPdest_2_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_debug_otherPdest_3_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_debug_otherPdest_4_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_debug_otherPdest_5_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_debug_otherPdest_6_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_debug_fuType_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_dirtyFs_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_1_dirtyVs_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_walk_v_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_commit_v_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_commit_w_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_realDestSize_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_interrupt_safe_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_wflags_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_fflags_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_vxsat_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_isRVC_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_isVset_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_isHls_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_isVls_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_vls_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_mmio_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_commitType_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_ftqIdx_flag_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_ftqIdx_value_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_ftqOffset_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_instrSize_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_needFlush_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_traceBlockInPipe_itype_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_traceBlockInPipe_iretire_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_traceBlockInPipe_ilastsize_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_debug_pc_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_debug_instr_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_debug_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_debug_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_debug_otherPdest_0_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_debug_otherPdest_1_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_debug_otherPdest_2_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_debug_otherPdest_3_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_debug_otherPdest_4_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_debug_otherPdest_5_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_debug_otherPdest_6_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_debug_fuType_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_dirtyFs_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_2_dirtyVs_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_walk_v_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_commit_v_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_commit_w_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_realDestSize_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_interrupt_safe_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_wflags_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_fflags_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_vxsat_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_isRVC_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_isVset_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_isHls_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_isVls_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_vls_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_mmio_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_commitType_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_ftqIdx_flag_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_ftqIdx_value_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_ftqOffset_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_instrSize_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_needFlush_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_traceBlockInPipe_itype_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_traceBlockInPipe_iretire_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_traceBlockInPipe_ilastsize_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_debug_pc_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_debug_instr_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_debug_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_debug_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_debug_otherPdest_0_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_debug_otherPdest_1_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_debug_otherPdest_2_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_debug_otherPdest_3_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_debug_otherPdest_4_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_debug_otherPdest_5_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_debug_otherPdest_6_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_debug_fuType_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_dirtyFs_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_3_dirtyVs_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_walk_v_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_commit_v_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_commit_w_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_realDestSize_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_interrupt_safe_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_wflags_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_fflags_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_vxsat_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_isRVC_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_isVset_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_isHls_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_isVls_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_vls_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_mmio_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_commitType_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_ftqIdx_flag_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_ftqIdx_value_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_ftqOffset_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_instrSize_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_needFlush_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_traceBlockInPipe_itype_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_traceBlockInPipe_iretire_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_traceBlockInPipe_ilastsize_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_debug_pc_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_debug_instr_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_debug_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_debug_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_debug_otherPdest_0_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_debug_otherPdest_1_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_debug_otherPdest_2_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_debug_otherPdest_3_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_debug_otherPdest_4_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_debug_otherPdest_5_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_debug_otherPdest_6_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_debug_fuType_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_dirtyFs_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_4_dirtyVs_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_walk_v_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_commit_v_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_commit_w_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_realDestSize_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_interrupt_safe_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_wflags_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_fflags_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_vxsat_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_isRVC_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_isVset_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_isHls_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_isVls_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_vls_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_mmio_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_commitType_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_ftqIdx_flag_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_ftqIdx_value_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_ftqOffset_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_instrSize_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_needFlush_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_traceBlockInPipe_itype_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_traceBlockInPipe_iretire_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_traceBlockInPipe_ilastsize_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_debug_pc_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_debug_instr_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_debug_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_debug_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_debug_otherPdest_0_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_debug_otherPdest_1_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_debug_otherPdest_2_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_debug_otherPdest_3_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_debug_otherPdest_4_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_debug_otherPdest_5_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_debug_otherPdest_6_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_debug_fuType_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_dirtyFs_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_5_dirtyVs_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_walk_v_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_commit_v_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_commit_w_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_realDestSize_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_interrupt_safe_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_wflags_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_fflags_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_vxsat_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_isRVC_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_isVset_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_isHls_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_isVls_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_vls_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_mmio_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_commitType_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_ftqIdx_flag_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_ftqIdx_value_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_ftqOffset_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_instrSize_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_needFlush_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_traceBlockInPipe_itype_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_traceBlockInPipe_iretire_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_traceBlockInPipe_ilastsize_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_debug_pc_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_debug_instr_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_debug_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_debug_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_debug_otherPdest_0_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_debug_otherPdest_1_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_debug_otherPdest_2_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_debug_otherPdest_3_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_debug_otherPdest_4_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_debug_otherPdest_5_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_debug_otherPdest_6_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_debug_fuType_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_dirtyFs_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_6_dirtyVs_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_walk_v_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_commit_v_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_commit_w_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_realDestSize_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_interrupt_safe_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_wflags_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_fflags_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_vxsat_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_isRVC_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_isVset_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_isHls_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_isVls_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_vls_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_mmio_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_commitType_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_ftqIdx_flag_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_ftqIdx_value_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_ftqOffset_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_instrSize_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_needFlush_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_traceBlockInPipe_itype_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_traceBlockInPipe_iretire_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_traceBlockInPipe_ilastsize_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_debug_pc_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_debug_instr_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_debug_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_debug_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_debug_otherPdest_0_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_debug_otherPdest_1_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_debug_otherPdest_2_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_debug_otherPdest_3_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_debug_otherPdest_4_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_debug_otherPdest_5_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_debug_otherPdest_6_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_debug_fuType_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_dirtyFs_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_info_7_dirtyVs_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_robIdx_0_flag_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_robIdx_0_value_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_robIdx_1_flag_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_robIdx_1_value_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_robIdx_2_flag_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_robIdx_2_value_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_robIdx_3_flag_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_robIdx_3_value_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_robIdx_4_flag_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_robIdx_4_value_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_robIdx_5_flag_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_robIdx_5_value_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_robIdx_6_flag_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_robIdx_6_value_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_robIdx_7_flag_cons{

}

constraint Rob_output_agent_xaction::default_io_commits_robIdx_7_value_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_blockCommit_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_0_valid_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_0_bits_ftqOffset_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_1_valid_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_1_bits_ftqOffset_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_2_valid_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_2_bits_ftqOffset_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_3_valid_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_3_bits_ftqOffset_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_4_valid_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_4_bits_ftqOffset_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_5_valid_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_5_bits_ftqOffset_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_6_valid_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_6_bits_ftqOffset_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_7_valid_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_7_bits_ftqOffset_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire_cons{

}

constraint Rob_output_agent_xaction::default_io_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_isCommit_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_commitValid_0_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_commitValid_1_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_commitValid_2_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_commitValid_3_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_commitValid_4_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_commitValid_5_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_isWalk_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_walkValid_0_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_walkValid_1_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_walkValid_2_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_walkValid_3_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_walkValid_4_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_walkValid_5_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_0_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_0_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_0_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_0_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_0_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_0_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_0_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_0_isMove_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_1_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_1_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_1_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_1_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_1_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_1_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_1_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_1_isMove_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_2_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_2_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_2_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_2_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_2_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_2_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_2_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_2_isMove_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_3_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_3_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_3_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_3_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_3_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_3_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_3_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_3_isMove_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_4_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_4_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_4_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_4_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_4_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_4_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_4_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_4_isMove_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_5_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_5_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_5_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_5_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_5_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_5_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_5_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_rabCommits_info_5_isMove_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_0_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_1_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_2_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_3_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_4_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_5_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_6_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_7_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_8_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_9_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_10_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_11_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_12_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_13_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_14_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_15_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_16_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_17_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_18_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_19_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_20_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_21_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_22_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_23_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_24_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_25_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_26_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_27_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_28_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_29_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_30_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_31_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_32_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_33_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_34_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_35_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_36_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_37_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_38_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_39_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_40_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_41_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_42_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_43_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_44_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_45_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_46_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_47_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_48_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_49_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_50_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_51_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_52_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_53_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_54_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_55_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_56_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_57_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_58_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_59_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_60_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_61_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_62_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_63_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_64_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_65_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_66_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_67_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_68_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_69_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_70_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_71_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_72_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_73_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_74_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_75_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_76_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_77_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_78_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_79_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_80_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_81_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_82_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_83_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_84_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_85_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_86_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_87_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_88_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_89_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_90_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_91_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_92_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_93_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_94_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_95_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_96_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_97_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_98_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_99_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_100_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_101_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_102_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_103_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_104_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_105_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_106_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_107_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_108_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_109_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_110_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_111_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_112_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_113_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_114_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_115_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_116_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_117_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_118_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_119_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_120_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_121_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_122_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_123_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_124_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_125_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_126_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_127_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_128_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_129_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_130_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_131_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_132_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_133_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_134_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_135_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_136_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_137_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_138_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_139_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_140_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_141_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_142_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_143_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_144_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_145_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_146_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_147_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_148_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_149_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_150_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_151_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_152_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_153_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_154_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_155_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_156_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_157_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_158_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_159_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_160_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_161_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_162_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_163_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_164_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_165_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_166_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_167_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_168_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_169_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_170_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_171_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_172_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_173_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_174_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_175_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_176_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_177_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_178_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_179_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_180_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_181_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_182_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_183_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_184_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_185_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_186_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_187_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_188_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_189_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_190_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_191_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_192_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_193_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_194_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_195_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_196_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_197_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_198_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_199_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_200_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_201_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_202_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_203_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_204_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_205_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_206_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_207_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_208_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_209_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_210_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_211_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_212_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_213_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_214_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_215_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_216_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_217_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_218_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_219_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_220_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_221_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_222_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_223_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_224_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_225_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_226_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_227_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_228_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_229_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_230_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_231_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_232_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_233_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_234_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_235_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_236_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_237_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_238_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_239_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_240_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_241_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_242_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_243_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_244_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_245_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_246_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_247_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_248_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_249_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_250_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_251_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_252_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_253_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_commitValid_254_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_0_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_0_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_0_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_0_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_0_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_0_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_0_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_1_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_1_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_1_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_1_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_1_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_1_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_1_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_2_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_2_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_2_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_2_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_2_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_2_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_2_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_3_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_3_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_3_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_3_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_3_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_3_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_3_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_4_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_4_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_4_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_4_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_4_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_4_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_4_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_5_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_5_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_5_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_5_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_5_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_5_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_5_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_6_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_6_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_6_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_6_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_6_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_6_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_6_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_7_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_7_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_7_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_7_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_7_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_7_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_7_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_8_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_8_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_8_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_8_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_8_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_8_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_8_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_9_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_9_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_9_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_9_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_9_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_9_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_9_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_10_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_10_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_10_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_10_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_10_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_10_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_10_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_11_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_11_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_11_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_11_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_11_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_11_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_11_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_12_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_12_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_12_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_12_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_12_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_12_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_12_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_13_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_13_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_13_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_13_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_13_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_13_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_13_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_14_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_14_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_14_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_14_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_14_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_14_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_14_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_15_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_15_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_15_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_15_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_15_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_15_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_15_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_16_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_16_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_16_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_16_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_16_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_16_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_16_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_17_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_17_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_17_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_17_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_17_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_17_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_17_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_18_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_18_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_18_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_18_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_18_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_18_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_18_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_19_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_19_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_19_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_19_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_19_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_19_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_19_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_20_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_20_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_20_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_20_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_20_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_20_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_20_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_21_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_21_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_21_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_21_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_21_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_21_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_21_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_22_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_22_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_22_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_22_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_22_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_22_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_22_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_23_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_23_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_23_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_23_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_23_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_23_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_23_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_24_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_24_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_24_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_24_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_24_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_24_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_24_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_25_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_25_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_25_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_25_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_25_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_25_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_25_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_26_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_26_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_26_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_26_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_26_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_26_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_26_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_27_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_27_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_27_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_27_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_27_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_27_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_27_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_28_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_28_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_28_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_28_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_28_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_28_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_28_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_29_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_29_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_29_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_29_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_29_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_29_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_29_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_30_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_30_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_30_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_30_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_30_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_30_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_30_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_31_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_31_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_31_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_31_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_31_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_31_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_31_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_32_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_32_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_32_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_32_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_32_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_32_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_32_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_33_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_33_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_33_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_33_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_33_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_33_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_33_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_34_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_34_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_34_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_34_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_34_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_34_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_34_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_35_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_35_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_35_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_35_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_35_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_35_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_35_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_36_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_36_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_36_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_36_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_36_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_36_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_36_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_37_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_37_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_37_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_37_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_37_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_37_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_37_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_38_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_38_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_38_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_38_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_38_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_38_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_38_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_39_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_39_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_39_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_39_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_39_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_39_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_39_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_40_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_40_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_40_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_40_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_40_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_40_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_40_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_41_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_41_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_41_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_41_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_41_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_41_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_41_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_42_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_42_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_42_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_42_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_42_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_42_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_42_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_43_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_43_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_43_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_43_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_43_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_43_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_43_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_44_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_44_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_44_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_44_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_44_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_44_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_44_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_45_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_45_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_45_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_45_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_45_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_45_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_45_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_46_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_46_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_46_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_46_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_46_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_46_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_46_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_47_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_47_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_47_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_47_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_47_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_47_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_47_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_48_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_48_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_48_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_48_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_48_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_48_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_48_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_49_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_49_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_49_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_49_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_49_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_49_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_49_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_50_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_50_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_50_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_50_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_50_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_50_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_50_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_51_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_51_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_51_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_51_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_51_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_51_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_51_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_52_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_52_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_52_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_52_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_52_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_52_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_52_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_53_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_53_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_53_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_53_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_53_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_53_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_53_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_54_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_54_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_54_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_54_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_54_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_54_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_54_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_55_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_55_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_55_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_55_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_55_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_55_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_55_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_56_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_56_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_56_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_56_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_56_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_56_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_56_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_57_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_57_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_57_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_57_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_57_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_57_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_57_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_58_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_58_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_58_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_58_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_58_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_58_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_58_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_59_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_59_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_59_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_59_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_59_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_59_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_59_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_60_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_60_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_60_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_60_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_60_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_60_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_60_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_61_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_61_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_61_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_61_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_61_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_61_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_61_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_62_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_62_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_62_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_62_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_62_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_62_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_62_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_63_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_63_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_63_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_63_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_63_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_63_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_63_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_64_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_64_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_64_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_64_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_64_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_64_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_64_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_65_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_65_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_65_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_65_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_65_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_65_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_65_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_66_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_66_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_66_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_66_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_66_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_66_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_66_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_67_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_67_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_67_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_67_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_67_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_67_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_67_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_68_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_68_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_68_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_68_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_68_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_68_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_68_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_69_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_69_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_69_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_69_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_69_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_69_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_69_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_70_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_70_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_70_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_70_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_70_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_70_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_70_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_71_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_71_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_71_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_71_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_71_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_71_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_71_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_72_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_72_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_72_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_72_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_72_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_72_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_72_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_73_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_73_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_73_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_73_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_73_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_73_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_73_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_74_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_74_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_74_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_74_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_74_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_74_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_74_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_75_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_75_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_75_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_75_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_75_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_75_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_75_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_76_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_76_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_76_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_76_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_76_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_76_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_76_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_77_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_77_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_77_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_77_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_77_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_77_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_77_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_78_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_78_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_78_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_78_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_78_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_78_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_78_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_79_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_79_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_79_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_79_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_79_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_79_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_79_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_80_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_80_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_80_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_80_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_80_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_80_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_80_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_81_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_81_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_81_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_81_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_81_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_81_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_81_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_82_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_82_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_82_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_82_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_82_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_82_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_82_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_83_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_83_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_83_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_83_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_83_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_83_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_83_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_84_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_84_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_84_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_84_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_84_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_84_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_84_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_85_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_85_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_85_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_85_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_85_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_85_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_85_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_86_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_86_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_86_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_86_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_86_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_86_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_86_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_87_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_87_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_87_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_87_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_87_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_87_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_87_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_88_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_88_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_88_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_88_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_88_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_88_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_88_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_89_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_89_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_89_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_89_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_89_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_89_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_89_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_90_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_90_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_90_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_90_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_90_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_90_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_90_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_91_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_91_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_91_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_91_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_91_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_91_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_91_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_92_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_92_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_92_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_92_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_92_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_92_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_92_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_93_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_93_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_93_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_93_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_93_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_93_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_93_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_94_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_94_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_94_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_94_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_94_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_94_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_94_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_95_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_95_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_95_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_95_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_95_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_95_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_95_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_96_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_96_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_96_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_96_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_96_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_96_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_96_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_97_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_97_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_97_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_97_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_97_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_97_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_97_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_98_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_98_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_98_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_98_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_98_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_98_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_98_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_99_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_99_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_99_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_99_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_99_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_99_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_99_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_100_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_100_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_100_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_100_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_100_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_100_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_100_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_101_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_101_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_101_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_101_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_101_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_101_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_101_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_102_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_102_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_102_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_102_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_102_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_102_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_102_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_103_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_103_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_103_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_103_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_103_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_103_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_103_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_104_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_104_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_104_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_104_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_104_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_104_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_104_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_105_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_105_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_105_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_105_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_105_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_105_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_105_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_106_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_106_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_106_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_106_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_106_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_106_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_106_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_107_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_107_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_107_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_107_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_107_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_107_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_107_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_108_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_108_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_108_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_108_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_108_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_108_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_108_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_109_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_109_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_109_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_109_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_109_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_109_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_109_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_110_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_110_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_110_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_110_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_110_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_110_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_110_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_111_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_111_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_111_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_111_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_111_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_111_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_111_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_112_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_112_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_112_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_112_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_112_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_112_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_112_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_113_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_113_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_113_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_113_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_113_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_113_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_113_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_114_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_114_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_114_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_114_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_114_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_114_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_114_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_115_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_115_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_115_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_115_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_115_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_115_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_115_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_116_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_116_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_116_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_116_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_116_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_116_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_116_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_117_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_117_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_117_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_117_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_117_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_117_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_117_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_118_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_118_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_118_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_118_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_118_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_118_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_118_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_119_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_119_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_119_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_119_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_119_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_119_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_119_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_120_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_120_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_120_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_120_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_120_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_120_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_120_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_121_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_121_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_121_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_121_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_121_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_121_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_121_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_122_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_122_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_122_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_122_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_122_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_122_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_122_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_123_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_123_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_123_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_123_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_123_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_123_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_123_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_124_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_124_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_124_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_124_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_124_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_124_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_124_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_125_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_125_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_125_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_125_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_125_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_125_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_125_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_126_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_126_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_126_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_126_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_126_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_126_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_126_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_127_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_127_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_127_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_127_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_127_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_127_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_127_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_128_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_128_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_128_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_128_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_128_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_128_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_128_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_129_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_129_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_129_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_129_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_129_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_129_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_129_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_130_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_130_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_130_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_130_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_130_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_130_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_130_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_131_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_131_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_131_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_131_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_131_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_131_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_131_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_132_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_132_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_132_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_132_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_132_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_132_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_132_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_133_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_133_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_133_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_133_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_133_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_133_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_133_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_134_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_134_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_134_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_134_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_134_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_134_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_134_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_135_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_135_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_135_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_135_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_135_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_135_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_135_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_136_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_136_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_136_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_136_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_136_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_136_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_136_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_137_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_137_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_137_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_137_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_137_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_137_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_137_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_138_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_138_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_138_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_138_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_138_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_138_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_138_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_139_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_139_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_139_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_139_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_139_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_139_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_139_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_140_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_140_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_140_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_140_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_140_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_140_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_140_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_141_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_141_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_141_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_141_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_141_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_141_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_141_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_142_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_142_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_142_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_142_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_142_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_142_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_142_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_143_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_143_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_143_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_143_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_143_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_143_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_143_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_144_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_144_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_144_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_144_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_144_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_144_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_144_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_145_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_145_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_145_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_145_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_145_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_145_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_145_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_146_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_146_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_146_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_146_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_146_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_146_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_146_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_147_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_147_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_147_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_147_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_147_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_147_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_147_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_148_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_148_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_148_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_148_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_148_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_148_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_148_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_149_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_149_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_149_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_149_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_149_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_149_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_149_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_150_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_150_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_150_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_150_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_150_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_150_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_150_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_151_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_151_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_151_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_151_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_151_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_151_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_151_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_152_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_152_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_152_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_152_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_152_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_152_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_152_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_153_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_153_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_153_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_153_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_153_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_153_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_153_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_154_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_154_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_154_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_154_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_154_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_154_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_154_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_155_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_155_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_155_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_155_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_155_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_155_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_155_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_156_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_156_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_156_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_156_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_156_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_156_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_156_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_157_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_157_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_157_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_157_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_157_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_157_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_157_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_158_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_158_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_158_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_158_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_158_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_158_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_158_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_159_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_159_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_159_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_159_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_159_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_159_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_159_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_160_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_160_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_160_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_160_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_160_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_160_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_160_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_161_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_161_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_161_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_161_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_161_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_161_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_161_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_162_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_162_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_162_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_162_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_162_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_162_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_162_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_163_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_163_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_163_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_163_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_163_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_163_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_163_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_164_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_164_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_164_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_164_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_164_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_164_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_164_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_165_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_165_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_165_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_165_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_165_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_165_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_165_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_166_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_166_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_166_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_166_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_166_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_166_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_166_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_167_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_167_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_167_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_167_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_167_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_167_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_167_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_168_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_168_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_168_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_168_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_168_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_168_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_168_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_169_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_169_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_169_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_169_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_169_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_169_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_169_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_170_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_170_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_170_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_170_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_170_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_170_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_170_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_171_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_171_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_171_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_171_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_171_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_171_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_171_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_172_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_172_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_172_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_172_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_172_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_172_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_172_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_173_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_173_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_173_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_173_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_173_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_173_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_173_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_174_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_174_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_174_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_174_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_174_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_174_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_174_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_175_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_175_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_175_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_175_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_175_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_175_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_175_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_176_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_176_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_176_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_176_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_176_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_176_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_176_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_177_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_177_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_177_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_177_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_177_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_177_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_177_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_178_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_178_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_178_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_178_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_178_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_178_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_178_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_179_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_179_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_179_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_179_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_179_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_179_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_179_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_180_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_180_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_180_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_180_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_180_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_180_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_180_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_181_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_181_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_181_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_181_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_181_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_181_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_181_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_182_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_182_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_182_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_182_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_182_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_182_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_182_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_183_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_183_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_183_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_183_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_183_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_183_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_183_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_184_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_184_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_184_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_184_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_184_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_184_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_184_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_185_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_185_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_185_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_185_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_185_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_185_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_185_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_186_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_186_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_186_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_186_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_186_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_186_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_186_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_187_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_187_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_187_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_187_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_187_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_187_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_187_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_188_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_188_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_188_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_188_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_188_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_188_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_188_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_189_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_189_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_189_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_189_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_189_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_189_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_189_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_190_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_190_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_190_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_190_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_190_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_190_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_190_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_191_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_191_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_191_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_191_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_191_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_191_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_191_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_192_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_192_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_192_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_192_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_192_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_192_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_192_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_193_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_193_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_193_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_193_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_193_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_193_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_193_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_194_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_194_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_194_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_194_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_194_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_194_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_194_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_195_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_195_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_195_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_195_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_195_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_195_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_195_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_196_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_196_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_196_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_196_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_196_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_196_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_196_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_197_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_197_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_197_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_197_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_197_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_197_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_197_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_198_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_198_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_198_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_198_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_198_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_198_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_198_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_199_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_199_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_199_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_199_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_199_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_199_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_199_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_200_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_200_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_200_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_200_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_200_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_200_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_200_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_201_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_201_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_201_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_201_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_201_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_201_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_201_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_202_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_202_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_202_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_202_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_202_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_202_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_202_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_203_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_203_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_203_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_203_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_203_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_203_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_203_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_204_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_204_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_204_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_204_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_204_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_204_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_204_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_205_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_205_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_205_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_205_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_205_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_205_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_205_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_206_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_206_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_206_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_206_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_206_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_206_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_206_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_207_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_207_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_207_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_207_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_207_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_207_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_207_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_208_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_208_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_208_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_208_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_208_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_208_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_208_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_209_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_209_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_209_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_209_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_209_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_209_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_209_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_210_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_210_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_210_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_210_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_210_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_210_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_210_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_211_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_211_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_211_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_211_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_211_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_211_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_211_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_212_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_212_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_212_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_212_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_212_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_212_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_212_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_213_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_213_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_213_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_213_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_213_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_213_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_213_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_214_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_214_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_214_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_214_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_214_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_214_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_214_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_215_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_215_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_215_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_215_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_215_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_215_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_215_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_216_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_216_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_216_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_216_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_216_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_216_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_216_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_217_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_217_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_217_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_217_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_217_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_217_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_217_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_218_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_218_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_218_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_218_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_218_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_218_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_218_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_219_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_219_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_219_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_219_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_219_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_219_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_219_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_220_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_220_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_220_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_220_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_220_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_220_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_220_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_221_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_221_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_221_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_221_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_221_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_221_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_221_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_222_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_222_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_222_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_222_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_222_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_222_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_222_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_223_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_223_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_223_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_223_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_223_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_223_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_223_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_224_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_224_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_224_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_224_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_224_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_224_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_224_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_225_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_225_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_225_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_225_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_225_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_225_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_225_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_226_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_226_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_226_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_226_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_226_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_226_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_226_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_227_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_227_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_227_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_227_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_227_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_227_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_227_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_228_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_228_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_228_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_228_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_228_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_228_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_228_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_229_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_229_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_229_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_229_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_229_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_229_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_229_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_230_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_230_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_230_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_230_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_230_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_230_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_230_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_231_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_231_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_231_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_231_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_231_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_231_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_231_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_232_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_232_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_232_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_232_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_232_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_232_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_232_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_233_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_233_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_233_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_233_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_233_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_233_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_233_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_234_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_234_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_234_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_234_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_234_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_234_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_234_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_235_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_235_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_235_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_235_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_235_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_235_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_235_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_236_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_236_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_236_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_236_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_236_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_236_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_236_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_237_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_237_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_237_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_237_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_237_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_237_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_237_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_238_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_238_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_238_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_238_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_238_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_238_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_238_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_239_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_239_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_239_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_239_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_239_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_239_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_239_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_240_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_240_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_240_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_240_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_240_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_240_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_240_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_241_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_241_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_241_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_241_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_241_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_241_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_241_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_242_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_242_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_242_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_242_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_242_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_242_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_242_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_243_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_243_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_243_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_243_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_243_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_243_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_243_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_244_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_244_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_244_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_244_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_244_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_244_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_244_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_245_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_245_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_245_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_245_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_245_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_245_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_245_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_246_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_246_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_246_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_246_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_246_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_246_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_246_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_247_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_247_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_247_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_247_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_247_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_247_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_247_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_248_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_248_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_248_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_248_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_248_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_248_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_248_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_249_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_249_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_249_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_249_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_249_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_249_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_249_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_250_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_250_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_250_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_250_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_250_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_250_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_250_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_251_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_251_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_251_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_251_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_251_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_251_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_251_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_252_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_252_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_252_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_252_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_252_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_252_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_252_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_253_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_253_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_253_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_253_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_253_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_253_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_253_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_254_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_254_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_254_rfWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_254_fpWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_254_vecWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_254_v0Wen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_254_vlWen_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_255_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_255_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_256_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_256_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_257_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_257_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_258_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_258_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_259_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_259_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_260_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_260_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_261_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_261_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_262_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_262_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_263_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_263_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_264_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_264_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_265_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_265_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_266_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_266_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_267_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_267_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_268_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_268_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_269_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_269_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_270_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_270_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_271_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_271_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_272_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_272_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_273_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_273_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_274_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_274_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_275_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_275_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_276_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_276_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_277_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_277_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_278_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_278_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_279_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_279_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_280_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_280_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_281_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_281_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_282_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_282_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_283_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_283_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_284_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_284_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_285_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_285_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_286_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_286_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_287_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_287_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_288_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_288_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_289_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_289_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_290_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_290_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_291_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_291_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_292_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_292_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_293_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_293_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_294_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_294_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_295_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_295_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_296_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_296_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_297_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_297_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_298_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_298_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_299_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_299_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_300_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_300_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_301_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_301_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_302_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_302_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_303_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_303_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_304_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_304_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_305_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_305_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_306_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_306_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_307_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_307_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_308_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_308_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_309_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_309_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_310_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_310_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_311_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_311_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_312_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_312_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_313_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_313_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_314_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_314_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_315_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_315_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_316_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_316_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_317_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_317_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_318_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_318_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_319_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_319_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_320_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_320_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_321_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_321_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_322_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_322_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_323_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_323_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_324_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_324_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_325_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_325_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_326_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_326_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_327_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_327_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_328_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_328_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_329_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_329_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_330_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_330_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_331_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_331_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_332_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_332_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_333_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_333_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_334_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_334_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_335_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_335_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_336_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_336_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_337_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_337_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_338_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_338_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_339_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_339_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_340_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_340_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_341_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_341_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_342_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_342_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_343_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_343_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_344_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_344_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_345_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_345_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_346_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_346_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_347_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_347_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_348_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_348_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_349_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_349_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_350_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_350_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_351_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_351_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_352_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_352_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_353_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_353_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_354_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_354_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_355_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_355_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_356_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_356_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_357_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_357_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_358_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_358_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_359_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_359_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_360_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_360_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_361_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_361_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_362_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_362_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_363_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_363_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_364_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_364_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_365_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_365_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_366_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_366_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_367_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_367_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_368_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_368_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_369_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_369_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_370_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_370_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_371_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_371_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_372_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_372_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_373_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_373_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_374_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_374_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_375_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_375_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_376_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_376_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_377_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_377_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_378_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_378_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_379_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_379_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_380_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_380_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_381_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_381_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_382_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_382_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_383_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_383_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_384_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_384_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_385_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_385_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_386_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_386_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_387_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_387_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_388_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_388_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_389_ldest_cons{

}

constraint Rob_output_agent_xaction::default_io_diffCommits_info_389_pdest_cons{

}

constraint Rob_output_agent_xaction::default_io_lsq_scommit_cons{

}

constraint Rob_output_agent_xaction::default_io_lsq_pendingMMIOld_cons{

}

constraint Rob_output_agent_xaction::default_io_lsq_pendingst_cons{

}

constraint Rob_output_agent_xaction::default_io_lsq_pendingPtr_flag_cons{

}

constraint Rob_output_agent_xaction::default_io_lsq_pendingPtr_value_cons{

}

constraint Rob_output_agent_xaction::default_io_robDeqPtr_flag_cons{

}

constraint Rob_output_agent_xaction::default_io_robDeqPtr_value_cons{

}

constraint Rob_output_agent_xaction::default_io_csr_fflags_valid_cons{

}

constraint Rob_output_agent_xaction::default_io_csr_fflags_bits_cons{

}

constraint Rob_output_agent_xaction::default_io_csr_vxsat_valid_cons{

}

constraint Rob_output_agent_xaction::default_io_csr_vxsat_bits_cons{

}

constraint Rob_output_agent_xaction::default_io_csr_vstart_valid_cons{

}

constraint Rob_output_agent_xaction::default_io_csr_vstart_bits_cons{

}

constraint Rob_output_agent_xaction::default_io_csr_dirty_fs_cons{

}

constraint Rob_output_agent_xaction::default_io_csr_dirty_vs_cons{

}

constraint Rob_output_agent_xaction::default_io_csr_perfinfo_retiredInstr_cons{

}

constraint Rob_output_agent_xaction::default_io_cpu_halt_cons{

}

constraint Rob_output_agent_xaction::default_io_wfi_wfiReq_cons{

}

constraint Rob_output_agent_xaction::default_io_toDecode_isResumeVType_cons{

}

constraint Rob_output_agent_xaction::default_io_toDecode_walkToArchVType_cons{

}

constraint Rob_output_agent_xaction::default_io_toDecode_walkVType_valid_cons{

}

constraint Rob_output_agent_xaction::default_io_toDecode_walkVType_bits_illegal_cons{

}

constraint Rob_output_agent_xaction::default_io_toDecode_walkVType_bits_vma_cons{

}

constraint Rob_output_agent_xaction::default_io_toDecode_walkVType_bits_vta_cons{

}

constraint Rob_output_agent_xaction::default_io_toDecode_walkVType_bits_vsew_cons{

}

constraint Rob_output_agent_xaction::default_io_toDecode_walkVType_bits_vlmul_cons{

}

constraint Rob_output_agent_xaction::default_io_toDecode_commitVType_vtype_valid_cons{

}

constraint Rob_output_agent_xaction::default_io_toDecode_commitVType_vtype_bits_illegal_cons{

}

constraint Rob_output_agent_xaction::default_io_toDecode_commitVType_vtype_bits_vma_cons{

}

constraint Rob_output_agent_xaction::default_io_toDecode_commitVType_vtype_bits_vta_cons{

}

constraint Rob_output_agent_xaction::default_io_toDecode_commitVType_vtype_bits_vsew_cons{

}

constraint Rob_output_agent_xaction::default_io_toDecode_commitVType_vtype_bits_vlmul_cons{

}

constraint Rob_output_agent_xaction::default_io_toDecode_commitVType_hasVsetvl_cons{

}

constraint Rob_output_agent_xaction::default_io_readGPAMemAddr_valid_cons{

}

constraint Rob_output_agent_xaction::default_io_readGPAMemAddr_bits_ftqPtr_value_cons{

}

constraint Rob_output_agent_xaction::default_io_readGPAMemAddr_bits_ftqOffset_cons{

}

constraint Rob_output_agent_xaction::default_io_toVecExcpMod_logicPhyRegMap_0_valid_cons{

}

constraint Rob_output_agent_xaction::default_io_toVecExcpMod_logicPhyRegMap_0_bits_lreg_cons{

}

constraint Rob_output_agent_xaction::default_io_toVecExcpMod_logicPhyRegMap_0_bits_preg_cons{

}

constraint Rob_output_agent_xaction::default_io_toVecExcpMod_logicPhyRegMap_1_valid_cons{

}

constraint Rob_output_agent_xaction::default_io_toVecExcpMod_logicPhyRegMap_1_bits_lreg_cons{

}

constraint Rob_output_agent_xaction::default_io_toVecExcpMod_logicPhyRegMap_1_bits_preg_cons{

}

constraint Rob_output_agent_xaction::default_io_toVecExcpMod_logicPhyRegMap_2_valid_cons{

}

constraint Rob_output_agent_xaction::default_io_toVecExcpMod_logicPhyRegMap_2_bits_lreg_cons{

}

constraint Rob_output_agent_xaction::default_io_toVecExcpMod_logicPhyRegMap_2_bits_preg_cons{

}

constraint Rob_output_agent_xaction::default_io_toVecExcpMod_logicPhyRegMap_3_valid_cons{

}

constraint Rob_output_agent_xaction::default_io_toVecExcpMod_logicPhyRegMap_3_bits_lreg_cons{

}

constraint Rob_output_agent_xaction::default_io_toVecExcpMod_logicPhyRegMap_3_bits_preg_cons{

}

constraint Rob_output_agent_xaction::default_io_toVecExcpMod_logicPhyRegMap_4_valid_cons{

}

constraint Rob_output_agent_xaction::default_io_toVecExcpMod_logicPhyRegMap_4_bits_lreg_cons{

}

constraint Rob_output_agent_xaction::default_io_toVecExcpMod_logicPhyRegMap_4_bits_preg_cons{

}

constraint Rob_output_agent_xaction::default_io_toVecExcpMod_logicPhyRegMap_5_valid_cons{

}

constraint Rob_output_agent_xaction::default_io_toVecExcpMod_logicPhyRegMap_5_bits_lreg_cons{

}

constraint Rob_output_agent_xaction::default_io_toVecExcpMod_logicPhyRegMap_5_bits_preg_cons{

}

constraint Rob_output_agent_xaction::default_io_toVecExcpMod_excpInfo_valid_cons{

}

constraint Rob_output_agent_xaction::default_io_toVecExcpMod_excpInfo_bits_vstart_cons{

}

constraint Rob_output_agent_xaction::default_io_toVecExcpMod_excpInfo_bits_vsew_cons{

}

constraint Rob_output_agent_xaction::default_io_toVecExcpMod_excpInfo_bits_veew_cons{

}

constraint Rob_output_agent_xaction::default_io_toVecExcpMod_excpInfo_bits_vlmul_cons{

}

constraint Rob_output_agent_xaction::default_io_toVecExcpMod_excpInfo_bits_nf_cons{

}

constraint Rob_output_agent_xaction::default_io_toVecExcpMod_excpInfo_bits_isStride_cons{

}

constraint Rob_output_agent_xaction::default_io_toVecExcpMod_excpInfo_bits_isIndexed_cons{

}

constraint Rob_output_agent_xaction::default_io_toVecExcpMod_excpInfo_bits_isWhole_cons{

}

constraint Rob_output_agent_xaction::default_io_toVecExcpMod_excpInfo_bits_isVlm_cons{

}

constraint Rob_output_agent_xaction::default_io_storeDebugInfo_1_pc_cons{

}

constraint Rob_output_agent_xaction::default_io_perf_0_value_cons{

}

constraint Rob_output_agent_xaction::default_io_perf_1_value_cons{

}

constraint Rob_output_agent_xaction::default_io_perf_2_value_cons{

}

constraint Rob_output_agent_xaction::default_io_perf_3_value_cons{

}

constraint Rob_output_agent_xaction::default_io_perf_4_value_cons{

}

constraint Rob_output_agent_xaction::default_io_perf_5_value_cons{

}

constraint Rob_output_agent_xaction::default_io_perf_6_value_cons{

}

constraint Rob_output_agent_xaction::default_io_perf_7_value_cons{

}

constraint Rob_output_agent_xaction::default_io_perf_8_value_cons{

}

constraint Rob_output_agent_xaction::default_io_perf_9_value_cons{

}

constraint Rob_output_agent_xaction::default_io_perf_10_value_cons{

}

constraint Rob_output_agent_xaction::default_io_perf_11_value_cons{

}

constraint Rob_output_agent_xaction::default_io_perf_12_value_cons{

}

constraint Rob_output_agent_xaction::default_io_perf_13_value_cons{

}

constraint Rob_output_agent_xaction::default_io_perf_14_value_cons{

}

constraint Rob_output_agent_xaction::default_io_perf_15_value_cons{

}

constraint Rob_output_agent_xaction::default_io_perf_16_value_cons{

}

constraint Rob_output_agent_xaction::default_io_perf_17_value_cons{

}

constraint Rob_output_agent_xaction::default_io_error_0_cons{

}

function Rob_output_agent_xaction::new(string name = "Rob_output_agent_xaction");
    super.new();
endfunction:new

function void Rob_output_agent_xaction::pack();
    super.pack();
endfunction:pack
function void Rob_output_agent_xaction::unpack();
    super.unpack();
endfunction:unpack
function void Rob_output_agent_xaction::pre_randomize();
    super.pre_randomize();
endfunction:pre_randomize
function void Rob_output_agent_xaction::post_randomize();
    super.post_randomize();
    //this.pack();
endfunction:post_randomize

function string Rob_output_agent_xaction::psdisplay(string prefix = "");
    string pkt_str;
    pkt_str = $sformatf("%s for packet[%0d] >>>>",prefix,this.pkt_index);
    pkt_str = $sformatf("%schannel_id=%0d ",pkt_str,this.channel_id);
    pkt_str = $sformatf("%sstart=%0f finish=%0f >>>>\n",pkt_str,this.start,this.finish);
    //foreach(this.pload_q[i]) begin
    //    pkt_str = $sformatf("%spload_q[%0d]=0x%2h  ",pkt_str,i,this.pload_q[i]);
    //end
    pkt_str = $sformatf("%sio_enq_canAccept = 0x%0h ",pkt_str,this.io_enq_canAccept);
    pkt_str = $sformatf("%sio_enq_canAcceptForDispatch = 0x%0h ",pkt_str,this.io_enq_canAcceptForDispatch);
    pkt_str = $sformatf("%sio_enq_isEmpty = 0x%0h ",pkt_str,this.io_enq_isEmpty);
    pkt_str = $sformatf("%sio_flushOut_valid = 0x%0h ",pkt_str,this.io_flushOut_valid);
    pkt_str = $sformatf("%sio_flushOut_bits_isRVC = 0x%0h ",pkt_str,this.io_flushOut_bits_isRVC);
    pkt_str = $sformatf("%sio_flushOut_bits_robIdx_flag = 0x%0h ",pkt_str,this.io_flushOut_bits_robIdx_flag);
    pkt_str = $sformatf("%sio_flushOut_bits_robIdx_value = 0x%0h ",pkt_str,this.io_flushOut_bits_robIdx_value);
    pkt_str = $sformatf("%sio_flushOut_bits_ftqIdx_flag = 0x%0h ",pkt_str,this.io_flushOut_bits_ftqIdx_flag);
    pkt_str = $sformatf("%sio_flushOut_bits_ftqIdx_value = 0x%0h ",pkt_str,this.io_flushOut_bits_ftqIdx_value);
    pkt_str = $sformatf("%sio_flushOut_bits_ftqOffset = 0x%0h ",pkt_str,this.io_flushOut_bits_ftqOffset);
    pkt_str = $sformatf("%sio_flushOut_bits_level = 0x%0h ",pkt_str,this.io_flushOut_bits_level);
    pkt_str = $sformatf("%sio_exception_valid = 0x%0h ",pkt_str,this.io_exception_valid);
    pkt_str = $sformatf("%sio_exception_bits_instr = 0x%0h ",pkt_str,this.io_exception_bits_instr);
    pkt_str = $sformatf("%sio_exception_bits_commitType = 0x%0h ",pkt_str,this.io_exception_bits_commitType);
    pkt_str = $sformatf("%sio_exception_bits_exceptionVec_0 = 0x%0h ",pkt_str,this.io_exception_bits_exceptionVec_0);
    pkt_str = $sformatf("%sio_exception_bits_exceptionVec_1 = 0x%0h ",pkt_str,this.io_exception_bits_exceptionVec_1);
    pkt_str = $sformatf("%sio_exception_bits_exceptionVec_2 = 0x%0h ",pkt_str,this.io_exception_bits_exceptionVec_2);
    pkt_str = $sformatf("%sio_exception_bits_exceptionVec_3 = 0x%0h ",pkt_str,this.io_exception_bits_exceptionVec_3);
    pkt_str = $sformatf("%sio_exception_bits_exceptionVec_4 = 0x%0h ",pkt_str,this.io_exception_bits_exceptionVec_4);
    pkt_str = $sformatf("%sio_exception_bits_exceptionVec_5 = 0x%0h ",pkt_str,this.io_exception_bits_exceptionVec_5);
    pkt_str = $sformatf("%sio_exception_bits_exceptionVec_6 = 0x%0h ",pkt_str,this.io_exception_bits_exceptionVec_6);
    pkt_str = $sformatf("%sio_exception_bits_exceptionVec_7 = 0x%0h ",pkt_str,this.io_exception_bits_exceptionVec_7);
    pkt_str = $sformatf("%sio_exception_bits_exceptionVec_8 = 0x%0h ",pkt_str,this.io_exception_bits_exceptionVec_8);
    pkt_str = $sformatf("%sio_exception_bits_exceptionVec_9 = 0x%0h ",pkt_str,this.io_exception_bits_exceptionVec_9);
    pkt_str = $sformatf("%sio_exception_bits_exceptionVec_10 = 0x%0h ",pkt_str,this.io_exception_bits_exceptionVec_10);
    pkt_str = $sformatf("%sio_exception_bits_exceptionVec_11 = 0x%0h ",pkt_str,this.io_exception_bits_exceptionVec_11);
    pkt_str = $sformatf("%sio_exception_bits_exceptionVec_12 = 0x%0h ",pkt_str,this.io_exception_bits_exceptionVec_12);
    pkt_str = $sformatf("%sio_exception_bits_exceptionVec_13 = 0x%0h ",pkt_str,this.io_exception_bits_exceptionVec_13);
    pkt_str = $sformatf("%sio_exception_bits_exceptionVec_14 = 0x%0h ",pkt_str,this.io_exception_bits_exceptionVec_14);
    pkt_str = $sformatf("%sio_exception_bits_exceptionVec_15 = 0x%0h ",pkt_str,this.io_exception_bits_exceptionVec_15);
    pkt_str = $sformatf("%sio_exception_bits_exceptionVec_16 = 0x%0h ",pkt_str,this.io_exception_bits_exceptionVec_16);
    pkt_str = $sformatf("%sio_exception_bits_exceptionVec_17 = 0x%0h ",pkt_str,this.io_exception_bits_exceptionVec_17);
    pkt_str = $sformatf("%sio_exception_bits_exceptionVec_18 = 0x%0h ",pkt_str,this.io_exception_bits_exceptionVec_18);
    pkt_str = $sformatf("%sio_exception_bits_exceptionVec_19 = 0x%0h ",pkt_str,this.io_exception_bits_exceptionVec_19);
    pkt_str = $sformatf("%sio_exception_bits_exceptionVec_20 = 0x%0h ",pkt_str,this.io_exception_bits_exceptionVec_20);
    pkt_str = $sformatf("%sio_exception_bits_exceptionVec_21 = 0x%0h ",pkt_str,this.io_exception_bits_exceptionVec_21);
    pkt_str = $sformatf("%sio_exception_bits_exceptionVec_22 = 0x%0h ",pkt_str,this.io_exception_bits_exceptionVec_22);
    pkt_str = $sformatf("%sio_exception_bits_exceptionVec_23 = 0x%0h ",pkt_str,this.io_exception_bits_exceptionVec_23);
    pkt_str = $sformatf("%sio_exception_bits_isPcBkpt = 0x%0h ",pkt_str,this.io_exception_bits_isPcBkpt);
    pkt_str = $sformatf("%sio_exception_bits_isFetchMalAddr = 0x%0h ",pkt_str,this.io_exception_bits_isFetchMalAddr);
    pkt_str = $sformatf("%sio_exception_bits_gpaddr = 0x%0h ",pkt_str,this.io_exception_bits_gpaddr);
    pkt_str = $sformatf("%sio_exception_bits_singleStep = 0x%0h ",pkt_str,this.io_exception_bits_singleStep);
    pkt_str = $sformatf("%sio_exception_bits_crossPageIPFFix = 0x%0h ",pkt_str,this.io_exception_bits_crossPageIPFFix);
    pkt_str = $sformatf("%sio_exception_bits_isInterrupt = 0x%0h ",pkt_str,this.io_exception_bits_isInterrupt);
    pkt_str = $sformatf("%sio_exception_bits_isHls = 0x%0h ",pkt_str,this.io_exception_bits_isHls);
    pkt_str = $sformatf("%sio_exception_bits_trigger = 0x%0h ",pkt_str,this.io_exception_bits_trigger);
    pkt_str = $sformatf("%sio_exception_bits_isForVSnonLeafPTE = 0x%0h ",pkt_str,this.io_exception_bits_isForVSnonLeafPTE);
    pkt_str = $sformatf("%sio_commits_isCommit = 0x%0h ",pkt_str,this.io_commits_isCommit);
    pkt_str = $sformatf("%sio_commits_commitValid_0 = 0x%0h ",pkt_str,this.io_commits_commitValid_0);
    pkt_str = $sformatf("%sio_commits_commitValid_1 = 0x%0h ",pkt_str,this.io_commits_commitValid_1);
    pkt_str = $sformatf("%sio_commits_commitValid_2 = 0x%0h ",pkt_str,this.io_commits_commitValid_2);
    pkt_str = $sformatf("%sio_commits_commitValid_3 = 0x%0h ",pkt_str,this.io_commits_commitValid_3);
    pkt_str = $sformatf("%sio_commits_commitValid_4 = 0x%0h ",pkt_str,this.io_commits_commitValid_4);
    pkt_str = $sformatf("%sio_commits_commitValid_5 = 0x%0h ",pkt_str,this.io_commits_commitValid_5);
    pkt_str = $sformatf("%sio_commits_commitValid_6 = 0x%0h ",pkt_str,this.io_commits_commitValid_6);
    pkt_str = $sformatf("%sio_commits_commitValid_7 = 0x%0h ",pkt_str,this.io_commits_commitValid_7);
    pkt_str = $sformatf("%sio_commits_isWalk = 0x%0h ",pkt_str,this.io_commits_isWalk);
    pkt_str = $sformatf("%sio_commits_walkValid_0 = 0x%0h ",pkt_str,this.io_commits_walkValid_0);
    pkt_str = $sformatf("%sio_commits_walkValid_1 = 0x%0h ",pkt_str,this.io_commits_walkValid_1);
    pkt_str = $sformatf("%sio_commits_walkValid_2 = 0x%0h ",pkt_str,this.io_commits_walkValid_2);
    pkt_str = $sformatf("%sio_commits_walkValid_3 = 0x%0h ",pkt_str,this.io_commits_walkValid_3);
    pkt_str = $sformatf("%sio_commits_walkValid_4 = 0x%0h ",pkt_str,this.io_commits_walkValid_4);
    pkt_str = $sformatf("%sio_commits_walkValid_5 = 0x%0h ",pkt_str,this.io_commits_walkValid_5);
    pkt_str = $sformatf("%sio_commits_walkValid_6 = 0x%0h ",pkt_str,this.io_commits_walkValid_6);
    pkt_str = $sformatf("%sio_commits_walkValid_7 = 0x%0h ",pkt_str,this.io_commits_walkValid_7);
    pkt_str = $sformatf("%sio_commits_info_0_walk_v = 0x%0h ",pkt_str,this.io_commits_info_0_walk_v);
    pkt_str = $sformatf("%sio_commits_info_0_commit_v = 0x%0h ",pkt_str,this.io_commits_info_0_commit_v);
    pkt_str = $sformatf("%sio_commits_info_0_commit_w = 0x%0h ",pkt_str,this.io_commits_info_0_commit_w);
    pkt_str = $sformatf("%sio_commits_info_0_realDestSize = 0x%0h ",pkt_str,this.io_commits_info_0_realDestSize);
    pkt_str = $sformatf("%sio_commits_info_0_interrupt_safe = 0x%0h ",pkt_str,this.io_commits_info_0_interrupt_safe);
    pkt_str = $sformatf("%sio_commits_info_0_wflags = 0x%0h ",pkt_str,this.io_commits_info_0_wflags);
    pkt_str = $sformatf("%sio_commits_info_0_fflags = 0x%0h ",pkt_str,this.io_commits_info_0_fflags);
    pkt_str = $sformatf("%sio_commits_info_0_vxsat = 0x%0h ",pkt_str,this.io_commits_info_0_vxsat);
    pkt_str = $sformatf("%sio_commits_info_0_isRVC = 0x%0h ",pkt_str,this.io_commits_info_0_isRVC);
    pkt_str = $sformatf("%sio_commits_info_0_isVset = 0x%0h ",pkt_str,this.io_commits_info_0_isVset);
    pkt_str = $sformatf("%sio_commits_info_0_isHls = 0x%0h ",pkt_str,this.io_commits_info_0_isHls);
    pkt_str = $sformatf("%sio_commits_info_0_isVls = 0x%0h ",pkt_str,this.io_commits_info_0_isVls);
    pkt_str = $sformatf("%sio_commits_info_0_vls = 0x%0h ",pkt_str,this.io_commits_info_0_vls);
    pkt_str = $sformatf("%sio_commits_info_0_mmio = 0x%0h ",pkt_str,this.io_commits_info_0_mmio);
    pkt_str = $sformatf("%sio_commits_info_0_commitType = 0x%0h ",pkt_str,this.io_commits_info_0_commitType);
    pkt_str = $sformatf("%sio_commits_info_0_ftqIdx_flag = 0x%0h ",pkt_str,this.io_commits_info_0_ftqIdx_flag);
    pkt_str = $sformatf("%sio_commits_info_0_ftqIdx_value = 0x%0h ",pkt_str,this.io_commits_info_0_ftqIdx_value);
    pkt_str = $sformatf("%sio_commits_info_0_ftqOffset = 0x%0h ",pkt_str,this.io_commits_info_0_ftqOffset);
    pkt_str = $sformatf("%sio_commits_info_0_instrSize = 0x%0h ",pkt_str,this.io_commits_info_0_instrSize);
    pkt_str = $sformatf("%sio_commits_info_0_fpWen = 0x%0h ",pkt_str,this.io_commits_info_0_fpWen);
    pkt_str = $sformatf("%sio_commits_info_0_rfWen = 0x%0h ",pkt_str,this.io_commits_info_0_rfWen);
    pkt_str = $sformatf("%sio_commits_info_0_needFlush = 0x%0h ",pkt_str,this.io_commits_info_0_needFlush);
    pkt_str = $sformatf("%sio_commits_info_0_traceBlockInPipe_itype = 0x%0h ",pkt_str,this.io_commits_info_0_traceBlockInPipe_itype);
    pkt_str = $sformatf("%sio_commits_info_0_traceBlockInPipe_iretire = 0x%0h ",pkt_str,this.io_commits_info_0_traceBlockInPipe_iretire);
    pkt_str = $sformatf("%sio_commits_info_0_traceBlockInPipe_ilastsize = 0x%0h ",pkt_str,this.io_commits_info_0_traceBlockInPipe_ilastsize);
    pkt_str = $sformatf("%sio_commits_info_0_debug_pc = 0x%0h ",pkt_str,this.io_commits_info_0_debug_pc);
    pkt_str = $sformatf("%sio_commits_info_0_debug_instr = 0x%0h ",pkt_str,this.io_commits_info_0_debug_instr);
    pkt_str = $sformatf("%sio_commits_info_0_debug_ldest = 0x%0h ",pkt_str,this.io_commits_info_0_debug_ldest);
    pkt_str = $sformatf("%sio_commits_info_0_debug_pdest = 0x%0h ",pkt_str,this.io_commits_info_0_debug_pdest);
    pkt_str = $sformatf("%sio_commits_info_0_debug_otherPdest_0 = 0x%0h ",pkt_str,this.io_commits_info_0_debug_otherPdest_0);
    pkt_str = $sformatf("%sio_commits_info_0_debug_otherPdest_1 = 0x%0h ",pkt_str,this.io_commits_info_0_debug_otherPdest_1);
    pkt_str = $sformatf("%sio_commits_info_0_debug_otherPdest_2 = 0x%0h ",pkt_str,this.io_commits_info_0_debug_otherPdest_2);
    pkt_str = $sformatf("%sio_commits_info_0_debug_otherPdest_3 = 0x%0h ",pkt_str,this.io_commits_info_0_debug_otherPdest_3);
    pkt_str = $sformatf("%sio_commits_info_0_debug_otherPdest_4 = 0x%0h ",pkt_str,this.io_commits_info_0_debug_otherPdest_4);
    pkt_str = $sformatf("%sio_commits_info_0_debug_otherPdest_5 = 0x%0h ",pkt_str,this.io_commits_info_0_debug_otherPdest_5);
    pkt_str = $sformatf("%sio_commits_info_0_debug_otherPdest_6 = 0x%0h ",pkt_str,this.io_commits_info_0_debug_otherPdest_6);
    pkt_str = $sformatf("%sio_commits_info_0_debug_fuType = 0x%0h ",pkt_str,this.io_commits_info_0_debug_fuType);
    pkt_str = $sformatf("%sio_commits_info_0_dirtyFs = 0x%0h ",pkt_str,this.io_commits_info_0_dirtyFs);
    pkt_str = $sformatf("%sio_commits_info_0_dirtyVs = 0x%0h ",pkt_str,this.io_commits_info_0_dirtyVs);
    pkt_str = $sformatf("%sio_commits_info_1_walk_v = 0x%0h ",pkt_str,this.io_commits_info_1_walk_v);
    pkt_str = $sformatf("%sio_commits_info_1_commit_v = 0x%0h ",pkt_str,this.io_commits_info_1_commit_v);
    pkt_str = $sformatf("%sio_commits_info_1_commit_w = 0x%0h ",pkt_str,this.io_commits_info_1_commit_w);
    pkt_str = $sformatf("%sio_commits_info_1_realDestSize = 0x%0h ",pkt_str,this.io_commits_info_1_realDestSize);
    pkt_str = $sformatf("%sio_commits_info_1_interrupt_safe = 0x%0h ",pkt_str,this.io_commits_info_1_interrupt_safe);
    pkt_str = $sformatf("%sio_commits_info_1_wflags = 0x%0h ",pkt_str,this.io_commits_info_1_wflags);
    pkt_str = $sformatf("%sio_commits_info_1_fflags = 0x%0h ",pkt_str,this.io_commits_info_1_fflags);
    pkt_str = $sformatf("%sio_commits_info_1_vxsat = 0x%0h ",pkt_str,this.io_commits_info_1_vxsat);
    pkt_str = $sformatf("%sio_commits_info_1_isRVC = 0x%0h ",pkt_str,this.io_commits_info_1_isRVC);
    pkt_str = $sformatf("%sio_commits_info_1_isVset = 0x%0h ",pkt_str,this.io_commits_info_1_isVset);
    pkt_str = $sformatf("%sio_commits_info_1_isHls = 0x%0h ",pkt_str,this.io_commits_info_1_isHls);
    pkt_str = $sformatf("%sio_commits_info_1_isVls = 0x%0h ",pkt_str,this.io_commits_info_1_isVls);
    pkt_str = $sformatf("%sio_commits_info_1_vls = 0x%0h ",pkt_str,this.io_commits_info_1_vls);
    pkt_str = $sformatf("%sio_commits_info_1_mmio = 0x%0h ",pkt_str,this.io_commits_info_1_mmio);
    pkt_str = $sformatf("%sio_commits_info_1_commitType = 0x%0h ",pkt_str,this.io_commits_info_1_commitType);
    pkt_str = $sformatf("%sio_commits_info_1_ftqIdx_flag = 0x%0h ",pkt_str,this.io_commits_info_1_ftqIdx_flag);
    pkt_str = $sformatf("%sio_commits_info_1_ftqIdx_value = 0x%0h ",pkt_str,this.io_commits_info_1_ftqIdx_value);
    pkt_str = $sformatf("%sio_commits_info_1_ftqOffset = 0x%0h ",pkt_str,this.io_commits_info_1_ftqOffset);
    pkt_str = $sformatf("%sio_commits_info_1_instrSize = 0x%0h ",pkt_str,this.io_commits_info_1_instrSize);
    pkt_str = $sformatf("%sio_commits_info_1_fpWen = 0x%0h ",pkt_str,this.io_commits_info_1_fpWen);
    pkt_str = $sformatf("%sio_commits_info_1_rfWen = 0x%0h ",pkt_str,this.io_commits_info_1_rfWen);
    pkt_str = $sformatf("%sio_commits_info_1_needFlush = 0x%0h ",pkt_str,this.io_commits_info_1_needFlush);
    pkt_str = $sformatf("%sio_commits_info_1_traceBlockInPipe_itype = 0x%0h ",pkt_str,this.io_commits_info_1_traceBlockInPipe_itype);
    pkt_str = $sformatf("%sio_commits_info_1_traceBlockInPipe_iretire = 0x%0h ",pkt_str,this.io_commits_info_1_traceBlockInPipe_iretire);
    pkt_str = $sformatf("%sio_commits_info_1_traceBlockInPipe_ilastsize = 0x%0h ",pkt_str,this.io_commits_info_1_traceBlockInPipe_ilastsize);
    pkt_str = $sformatf("%sio_commits_info_1_debug_pc = 0x%0h ",pkt_str,this.io_commits_info_1_debug_pc);
    pkt_str = $sformatf("%sio_commits_info_1_debug_instr = 0x%0h ",pkt_str,this.io_commits_info_1_debug_instr);
    pkt_str = $sformatf("%sio_commits_info_1_debug_ldest = 0x%0h ",pkt_str,this.io_commits_info_1_debug_ldest);
    pkt_str = $sformatf("%sio_commits_info_1_debug_pdest = 0x%0h ",pkt_str,this.io_commits_info_1_debug_pdest);
    pkt_str = $sformatf("%sio_commits_info_1_debug_otherPdest_0 = 0x%0h ",pkt_str,this.io_commits_info_1_debug_otherPdest_0);
    pkt_str = $sformatf("%sio_commits_info_1_debug_otherPdest_1 = 0x%0h ",pkt_str,this.io_commits_info_1_debug_otherPdest_1);
    pkt_str = $sformatf("%sio_commits_info_1_debug_otherPdest_2 = 0x%0h ",pkt_str,this.io_commits_info_1_debug_otherPdest_2);
    pkt_str = $sformatf("%sio_commits_info_1_debug_otherPdest_3 = 0x%0h ",pkt_str,this.io_commits_info_1_debug_otherPdest_3);
    pkt_str = $sformatf("%sio_commits_info_1_debug_otherPdest_4 = 0x%0h ",pkt_str,this.io_commits_info_1_debug_otherPdest_4);
    pkt_str = $sformatf("%sio_commits_info_1_debug_otherPdest_5 = 0x%0h ",pkt_str,this.io_commits_info_1_debug_otherPdest_5);
    pkt_str = $sformatf("%sio_commits_info_1_debug_otherPdest_6 = 0x%0h ",pkt_str,this.io_commits_info_1_debug_otherPdest_6);
    pkt_str = $sformatf("%sio_commits_info_1_debug_fuType = 0x%0h ",pkt_str,this.io_commits_info_1_debug_fuType);
    pkt_str = $sformatf("%sio_commits_info_1_dirtyFs = 0x%0h ",pkt_str,this.io_commits_info_1_dirtyFs);
    pkt_str = $sformatf("%sio_commits_info_1_dirtyVs = 0x%0h ",pkt_str,this.io_commits_info_1_dirtyVs);
    pkt_str = $sformatf("%sio_commits_info_2_walk_v = 0x%0h ",pkt_str,this.io_commits_info_2_walk_v);
    pkt_str = $sformatf("%sio_commits_info_2_commit_v = 0x%0h ",pkt_str,this.io_commits_info_2_commit_v);
    pkt_str = $sformatf("%sio_commits_info_2_commit_w = 0x%0h ",pkt_str,this.io_commits_info_2_commit_w);
    pkt_str = $sformatf("%sio_commits_info_2_realDestSize = 0x%0h ",pkt_str,this.io_commits_info_2_realDestSize);
    pkt_str = $sformatf("%sio_commits_info_2_interrupt_safe = 0x%0h ",pkt_str,this.io_commits_info_2_interrupt_safe);
    pkt_str = $sformatf("%sio_commits_info_2_wflags = 0x%0h ",pkt_str,this.io_commits_info_2_wflags);
    pkt_str = $sformatf("%sio_commits_info_2_fflags = 0x%0h ",pkt_str,this.io_commits_info_2_fflags);
    pkt_str = $sformatf("%sio_commits_info_2_vxsat = 0x%0h ",pkt_str,this.io_commits_info_2_vxsat);
    pkt_str = $sformatf("%sio_commits_info_2_isRVC = 0x%0h ",pkt_str,this.io_commits_info_2_isRVC);
    pkt_str = $sformatf("%sio_commits_info_2_isVset = 0x%0h ",pkt_str,this.io_commits_info_2_isVset);
    pkt_str = $sformatf("%sio_commits_info_2_isHls = 0x%0h ",pkt_str,this.io_commits_info_2_isHls);
    pkt_str = $sformatf("%sio_commits_info_2_isVls = 0x%0h ",pkt_str,this.io_commits_info_2_isVls);
    pkt_str = $sformatf("%sio_commits_info_2_vls = 0x%0h ",pkt_str,this.io_commits_info_2_vls);
    pkt_str = $sformatf("%sio_commits_info_2_mmio = 0x%0h ",pkt_str,this.io_commits_info_2_mmio);
    pkt_str = $sformatf("%sio_commits_info_2_commitType = 0x%0h ",pkt_str,this.io_commits_info_2_commitType);
    pkt_str = $sformatf("%sio_commits_info_2_ftqIdx_flag = 0x%0h ",pkt_str,this.io_commits_info_2_ftqIdx_flag);
    pkt_str = $sformatf("%sio_commits_info_2_ftqIdx_value = 0x%0h ",pkt_str,this.io_commits_info_2_ftqIdx_value);
    pkt_str = $sformatf("%sio_commits_info_2_ftqOffset = 0x%0h ",pkt_str,this.io_commits_info_2_ftqOffset);
    pkt_str = $sformatf("%sio_commits_info_2_instrSize = 0x%0h ",pkt_str,this.io_commits_info_2_instrSize);
    pkt_str = $sformatf("%sio_commits_info_2_fpWen = 0x%0h ",pkt_str,this.io_commits_info_2_fpWen);
    pkt_str = $sformatf("%sio_commits_info_2_rfWen = 0x%0h ",pkt_str,this.io_commits_info_2_rfWen);
    pkt_str = $sformatf("%sio_commits_info_2_needFlush = 0x%0h ",pkt_str,this.io_commits_info_2_needFlush);
    pkt_str = $sformatf("%sio_commits_info_2_traceBlockInPipe_itype = 0x%0h ",pkt_str,this.io_commits_info_2_traceBlockInPipe_itype);
    pkt_str = $sformatf("%sio_commits_info_2_traceBlockInPipe_iretire = 0x%0h ",pkt_str,this.io_commits_info_2_traceBlockInPipe_iretire);
    pkt_str = $sformatf("%sio_commits_info_2_traceBlockInPipe_ilastsize = 0x%0h ",pkt_str,this.io_commits_info_2_traceBlockInPipe_ilastsize);
    pkt_str = $sformatf("%sio_commits_info_2_debug_pc = 0x%0h ",pkt_str,this.io_commits_info_2_debug_pc);
    pkt_str = $sformatf("%sio_commits_info_2_debug_instr = 0x%0h ",pkt_str,this.io_commits_info_2_debug_instr);
    pkt_str = $sformatf("%sio_commits_info_2_debug_ldest = 0x%0h ",pkt_str,this.io_commits_info_2_debug_ldest);
    pkt_str = $sformatf("%sio_commits_info_2_debug_pdest = 0x%0h ",pkt_str,this.io_commits_info_2_debug_pdest);
    pkt_str = $sformatf("%sio_commits_info_2_debug_otherPdest_0 = 0x%0h ",pkt_str,this.io_commits_info_2_debug_otherPdest_0);
    pkt_str = $sformatf("%sio_commits_info_2_debug_otherPdest_1 = 0x%0h ",pkt_str,this.io_commits_info_2_debug_otherPdest_1);
    pkt_str = $sformatf("%sio_commits_info_2_debug_otherPdest_2 = 0x%0h ",pkt_str,this.io_commits_info_2_debug_otherPdest_2);
    pkt_str = $sformatf("%sio_commits_info_2_debug_otherPdest_3 = 0x%0h ",pkt_str,this.io_commits_info_2_debug_otherPdest_3);
    pkt_str = $sformatf("%sio_commits_info_2_debug_otherPdest_4 = 0x%0h ",pkt_str,this.io_commits_info_2_debug_otherPdest_4);
    pkt_str = $sformatf("%sio_commits_info_2_debug_otherPdest_5 = 0x%0h ",pkt_str,this.io_commits_info_2_debug_otherPdest_5);
    pkt_str = $sformatf("%sio_commits_info_2_debug_otherPdest_6 = 0x%0h ",pkt_str,this.io_commits_info_2_debug_otherPdest_6);
    pkt_str = $sformatf("%sio_commits_info_2_debug_fuType = 0x%0h ",pkt_str,this.io_commits_info_2_debug_fuType);
    pkt_str = $sformatf("%sio_commits_info_2_dirtyFs = 0x%0h ",pkt_str,this.io_commits_info_2_dirtyFs);
    pkt_str = $sformatf("%sio_commits_info_2_dirtyVs = 0x%0h ",pkt_str,this.io_commits_info_2_dirtyVs);
    pkt_str = $sformatf("%sio_commits_info_3_walk_v = 0x%0h ",pkt_str,this.io_commits_info_3_walk_v);
    pkt_str = $sformatf("%sio_commits_info_3_commit_v = 0x%0h ",pkt_str,this.io_commits_info_3_commit_v);
    pkt_str = $sformatf("%sio_commits_info_3_commit_w = 0x%0h ",pkt_str,this.io_commits_info_3_commit_w);
    pkt_str = $sformatf("%sio_commits_info_3_realDestSize = 0x%0h ",pkt_str,this.io_commits_info_3_realDestSize);
    pkt_str = $sformatf("%sio_commits_info_3_interrupt_safe = 0x%0h ",pkt_str,this.io_commits_info_3_interrupt_safe);
    pkt_str = $sformatf("%sio_commits_info_3_wflags = 0x%0h ",pkt_str,this.io_commits_info_3_wflags);
    pkt_str = $sformatf("%sio_commits_info_3_fflags = 0x%0h ",pkt_str,this.io_commits_info_3_fflags);
    pkt_str = $sformatf("%sio_commits_info_3_vxsat = 0x%0h ",pkt_str,this.io_commits_info_3_vxsat);
    pkt_str = $sformatf("%sio_commits_info_3_isRVC = 0x%0h ",pkt_str,this.io_commits_info_3_isRVC);
    pkt_str = $sformatf("%sio_commits_info_3_isVset = 0x%0h ",pkt_str,this.io_commits_info_3_isVset);
    pkt_str = $sformatf("%sio_commits_info_3_isHls = 0x%0h ",pkt_str,this.io_commits_info_3_isHls);
    pkt_str = $sformatf("%sio_commits_info_3_isVls = 0x%0h ",pkt_str,this.io_commits_info_3_isVls);
    pkt_str = $sformatf("%sio_commits_info_3_vls = 0x%0h ",pkt_str,this.io_commits_info_3_vls);
    pkt_str = $sformatf("%sio_commits_info_3_mmio = 0x%0h ",pkt_str,this.io_commits_info_3_mmio);
    pkt_str = $sformatf("%sio_commits_info_3_commitType = 0x%0h ",pkt_str,this.io_commits_info_3_commitType);
    pkt_str = $sformatf("%sio_commits_info_3_ftqIdx_flag = 0x%0h ",pkt_str,this.io_commits_info_3_ftqIdx_flag);
    pkt_str = $sformatf("%sio_commits_info_3_ftqIdx_value = 0x%0h ",pkt_str,this.io_commits_info_3_ftqIdx_value);
    pkt_str = $sformatf("%sio_commits_info_3_ftqOffset = 0x%0h ",pkt_str,this.io_commits_info_3_ftqOffset);
    pkt_str = $sformatf("%sio_commits_info_3_instrSize = 0x%0h ",pkt_str,this.io_commits_info_3_instrSize);
    pkt_str = $sformatf("%sio_commits_info_3_fpWen = 0x%0h ",pkt_str,this.io_commits_info_3_fpWen);
    pkt_str = $sformatf("%sio_commits_info_3_rfWen = 0x%0h ",pkt_str,this.io_commits_info_3_rfWen);
    pkt_str = $sformatf("%sio_commits_info_3_needFlush = 0x%0h ",pkt_str,this.io_commits_info_3_needFlush);
    pkt_str = $sformatf("%sio_commits_info_3_traceBlockInPipe_itype = 0x%0h ",pkt_str,this.io_commits_info_3_traceBlockInPipe_itype);
    pkt_str = $sformatf("%sio_commits_info_3_traceBlockInPipe_iretire = 0x%0h ",pkt_str,this.io_commits_info_3_traceBlockInPipe_iretire);
    pkt_str = $sformatf("%sio_commits_info_3_traceBlockInPipe_ilastsize = 0x%0h ",pkt_str,this.io_commits_info_3_traceBlockInPipe_ilastsize);
    pkt_str = $sformatf("%sio_commits_info_3_debug_pc = 0x%0h ",pkt_str,this.io_commits_info_3_debug_pc);
    pkt_str = $sformatf("%sio_commits_info_3_debug_instr = 0x%0h ",pkt_str,this.io_commits_info_3_debug_instr);
    pkt_str = $sformatf("%sio_commits_info_3_debug_ldest = 0x%0h ",pkt_str,this.io_commits_info_3_debug_ldest);
    pkt_str = $sformatf("%sio_commits_info_3_debug_pdest = 0x%0h ",pkt_str,this.io_commits_info_3_debug_pdest);
    pkt_str = $sformatf("%sio_commits_info_3_debug_otherPdest_0 = 0x%0h ",pkt_str,this.io_commits_info_3_debug_otherPdest_0);
    pkt_str = $sformatf("%sio_commits_info_3_debug_otherPdest_1 = 0x%0h ",pkt_str,this.io_commits_info_3_debug_otherPdest_1);
    pkt_str = $sformatf("%sio_commits_info_3_debug_otherPdest_2 = 0x%0h ",pkt_str,this.io_commits_info_3_debug_otherPdest_2);
    pkt_str = $sformatf("%sio_commits_info_3_debug_otherPdest_3 = 0x%0h ",pkt_str,this.io_commits_info_3_debug_otherPdest_3);
    pkt_str = $sformatf("%sio_commits_info_3_debug_otherPdest_4 = 0x%0h ",pkt_str,this.io_commits_info_3_debug_otherPdest_4);
    pkt_str = $sformatf("%sio_commits_info_3_debug_otherPdest_5 = 0x%0h ",pkt_str,this.io_commits_info_3_debug_otherPdest_5);
    pkt_str = $sformatf("%sio_commits_info_3_debug_otherPdest_6 = 0x%0h ",pkt_str,this.io_commits_info_3_debug_otherPdest_6);
    pkt_str = $sformatf("%sio_commits_info_3_debug_fuType = 0x%0h ",pkt_str,this.io_commits_info_3_debug_fuType);
    pkt_str = $sformatf("%sio_commits_info_3_dirtyFs = 0x%0h ",pkt_str,this.io_commits_info_3_dirtyFs);
    pkt_str = $sformatf("%sio_commits_info_3_dirtyVs = 0x%0h ",pkt_str,this.io_commits_info_3_dirtyVs);
    pkt_str = $sformatf("%sio_commits_info_4_walk_v = 0x%0h ",pkt_str,this.io_commits_info_4_walk_v);
    pkt_str = $sformatf("%sio_commits_info_4_commit_v = 0x%0h ",pkt_str,this.io_commits_info_4_commit_v);
    pkt_str = $sformatf("%sio_commits_info_4_commit_w = 0x%0h ",pkt_str,this.io_commits_info_4_commit_w);
    pkt_str = $sformatf("%sio_commits_info_4_realDestSize = 0x%0h ",pkt_str,this.io_commits_info_4_realDestSize);
    pkt_str = $sformatf("%sio_commits_info_4_interrupt_safe = 0x%0h ",pkt_str,this.io_commits_info_4_interrupt_safe);
    pkt_str = $sformatf("%sio_commits_info_4_wflags = 0x%0h ",pkt_str,this.io_commits_info_4_wflags);
    pkt_str = $sformatf("%sio_commits_info_4_fflags = 0x%0h ",pkt_str,this.io_commits_info_4_fflags);
    pkt_str = $sformatf("%sio_commits_info_4_vxsat = 0x%0h ",pkt_str,this.io_commits_info_4_vxsat);
    pkt_str = $sformatf("%sio_commits_info_4_isRVC = 0x%0h ",pkt_str,this.io_commits_info_4_isRVC);
    pkt_str = $sformatf("%sio_commits_info_4_isVset = 0x%0h ",pkt_str,this.io_commits_info_4_isVset);
    pkt_str = $sformatf("%sio_commits_info_4_isHls = 0x%0h ",pkt_str,this.io_commits_info_4_isHls);
    pkt_str = $sformatf("%sio_commits_info_4_isVls = 0x%0h ",pkt_str,this.io_commits_info_4_isVls);
    pkt_str = $sformatf("%sio_commits_info_4_vls = 0x%0h ",pkt_str,this.io_commits_info_4_vls);
    pkt_str = $sformatf("%sio_commits_info_4_mmio = 0x%0h ",pkt_str,this.io_commits_info_4_mmio);
    pkt_str = $sformatf("%sio_commits_info_4_commitType = 0x%0h ",pkt_str,this.io_commits_info_4_commitType);
    pkt_str = $sformatf("%sio_commits_info_4_ftqIdx_flag = 0x%0h ",pkt_str,this.io_commits_info_4_ftqIdx_flag);
    pkt_str = $sformatf("%sio_commits_info_4_ftqIdx_value = 0x%0h ",pkt_str,this.io_commits_info_4_ftqIdx_value);
    pkt_str = $sformatf("%sio_commits_info_4_ftqOffset = 0x%0h ",pkt_str,this.io_commits_info_4_ftqOffset);
    pkt_str = $sformatf("%sio_commits_info_4_instrSize = 0x%0h ",pkt_str,this.io_commits_info_4_instrSize);
    pkt_str = $sformatf("%sio_commits_info_4_fpWen = 0x%0h ",pkt_str,this.io_commits_info_4_fpWen);
    pkt_str = $sformatf("%sio_commits_info_4_rfWen = 0x%0h ",pkt_str,this.io_commits_info_4_rfWen);
    pkt_str = $sformatf("%sio_commits_info_4_needFlush = 0x%0h ",pkt_str,this.io_commits_info_4_needFlush);
    pkt_str = $sformatf("%sio_commits_info_4_traceBlockInPipe_itype = 0x%0h ",pkt_str,this.io_commits_info_4_traceBlockInPipe_itype);
    pkt_str = $sformatf("%sio_commits_info_4_traceBlockInPipe_iretire = 0x%0h ",pkt_str,this.io_commits_info_4_traceBlockInPipe_iretire);
    pkt_str = $sformatf("%sio_commits_info_4_traceBlockInPipe_ilastsize = 0x%0h ",pkt_str,this.io_commits_info_4_traceBlockInPipe_ilastsize);
    pkt_str = $sformatf("%sio_commits_info_4_debug_pc = 0x%0h ",pkt_str,this.io_commits_info_4_debug_pc);
    pkt_str = $sformatf("%sio_commits_info_4_debug_instr = 0x%0h ",pkt_str,this.io_commits_info_4_debug_instr);
    pkt_str = $sformatf("%sio_commits_info_4_debug_ldest = 0x%0h ",pkt_str,this.io_commits_info_4_debug_ldest);
    pkt_str = $sformatf("%sio_commits_info_4_debug_pdest = 0x%0h ",pkt_str,this.io_commits_info_4_debug_pdest);
    pkt_str = $sformatf("%sio_commits_info_4_debug_otherPdest_0 = 0x%0h ",pkt_str,this.io_commits_info_4_debug_otherPdest_0);
    pkt_str = $sformatf("%sio_commits_info_4_debug_otherPdest_1 = 0x%0h ",pkt_str,this.io_commits_info_4_debug_otherPdest_1);
    pkt_str = $sformatf("%sio_commits_info_4_debug_otherPdest_2 = 0x%0h ",pkt_str,this.io_commits_info_4_debug_otherPdest_2);
    pkt_str = $sformatf("%sio_commits_info_4_debug_otherPdest_3 = 0x%0h ",pkt_str,this.io_commits_info_4_debug_otherPdest_3);
    pkt_str = $sformatf("%sio_commits_info_4_debug_otherPdest_4 = 0x%0h ",pkt_str,this.io_commits_info_4_debug_otherPdest_4);
    pkt_str = $sformatf("%sio_commits_info_4_debug_otherPdest_5 = 0x%0h ",pkt_str,this.io_commits_info_4_debug_otherPdest_5);
    pkt_str = $sformatf("%sio_commits_info_4_debug_otherPdest_6 = 0x%0h ",pkt_str,this.io_commits_info_4_debug_otherPdest_6);
    pkt_str = $sformatf("%sio_commits_info_4_debug_fuType = 0x%0h ",pkt_str,this.io_commits_info_4_debug_fuType);
    pkt_str = $sformatf("%sio_commits_info_4_dirtyFs = 0x%0h ",pkt_str,this.io_commits_info_4_dirtyFs);
    pkt_str = $sformatf("%sio_commits_info_4_dirtyVs = 0x%0h ",pkt_str,this.io_commits_info_4_dirtyVs);
    pkt_str = $sformatf("%sio_commits_info_5_walk_v = 0x%0h ",pkt_str,this.io_commits_info_5_walk_v);
    pkt_str = $sformatf("%sio_commits_info_5_commit_v = 0x%0h ",pkt_str,this.io_commits_info_5_commit_v);
    pkt_str = $sformatf("%sio_commits_info_5_commit_w = 0x%0h ",pkt_str,this.io_commits_info_5_commit_w);
    pkt_str = $sformatf("%sio_commits_info_5_realDestSize = 0x%0h ",pkt_str,this.io_commits_info_5_realDestSize);
    pkt_str = $sformatf("%sio_commits_info_5_interrupt_safe = 0x%0h ",pkt_str,this.io_commits_info_5_interrupt_safe);
    pkt_str = $sformatf("%sio_commits_info_5_wflags = 0x%0h ",pkt_str,this.io_commits_info_5_wflags);
    pkt_str = $sformatf("%sio_commits_info_5_fflags = 0x%0h ",pkt_str,this.io_commits_info_5_fflags);
    pkt_str = $sformatf("%sio_commits_info_5_vxsat = 0x%0h ",pkt_str,this.io_commits_info_5_vxsat);
    pkt_str = $sformatf("%sio_commits_info_5_isRVC = 0x%0h ",pkt_str,this.io_commits_info_5_isRVC);
    pkt_str = $sformatf("%sio_commits_info_5_isVset = 0x%0h ",pkt_str,this.io_commits_info_5_isVset);
    pkt_str = $sformatf("%sio_commits_info_5_isHls = 0x%0h ",pkt_str,this.io_commits_info_5_isHls);
    pkt_str = $sformatf("%sio_commits_info_5_isVls = 0x%0h ",pkt_str,this.io_commits_info_5_isVls);
    pkt_str = $sformatf("%sio_commits_info_5_vls = 0x%0h ",pkt_str,this.io_commits_info_5_vls);
    pkt_str = $sformatf("%sio_commits_info_5_mmio = 0x%0h ",pkt_str,this.io_commits_info_5_mmio);
    pkt_str = $sformatf("%sio_commits_info_5_commitType = 0x%0h ",pkt_str,this.io_commits_info_5_commitType);
    pkt_str = $sformatf("%sio_commits_info_5_ftqIdx_flag = 0x%0h ",pkt_str,this.io_commits_info_5_ftqIdx_flag);
    pkt_str = $sformatf("%sio_commits_info_5_ftqIdx_value = 0x%0h ",pkt_str,this.io_commits_info_5_ftqIdx_value);
    pkt_str = $sformatf("%sio_commits_info_5_ftqOffset = 0x%0h ",pkt_str,this.io_commits_info_5_ftqOffset);
    pkt_str = $sformatf("%sio_commits_info_5_instrSize = 0x%0h ",pkt_str,this.io_commits_info_5_instrSize);
    pkt_str = $sformatf("%sio_commits_info_5_fpWen = 0x%0h ",pkt_str,this.io_commits_info_5_fpWen);
    pkt_str = $sformatf("%sio_commits_info_5_rfWen = 0x%0h ",pkt_str,this.io_commits_info_5_rfWen);
    pkt_str = $sformatf("%sio_commits_info_5_needFlush = 0x%0h ",pkt_str,this.io_commits_info_5_needFlush);
    pkt_str = $sformatf("%sio_commits_info_5_traceBlockInPipe_itype = 0x%0h ",pkt_str,this.io_commits_info_5_traceBlockInPipe_itype);
    pkt_str = $sformatf("%sio_commits_info_5_traceBlockInPipe_iretire = 0x%0h ",pkt_str,this.io_commits_info_5_traceBlockInPipe_iretire);
    pkt_str = $sformatf("%sio_commits_info_5_traceBlockInPipe_ilastsize = 0x%0h ",pkt_str,this.io_commits_info_5_traceBlockInPipe_ilastsize);
    pkt_str = $sformatf("%sio_commits_info_5_debug_pc = 0x%0h ",pkt_str,this.io_commits_info_5_debug_pc);
    pkt_str = $sformatf("%sio_commits_info_5_debug_instr = 0x%0h ",pkt_str,this.io_commits_info_5_debug_instr);
    pkt_str = $sformatf("%sio_commits_info_5_debug_ldest = 0x%0h ",pkt_str,this.io_commits_info_5_debug_ldest);
    pkt_str = $sformatf("%sio_commits_info_5_debug_pdest = 0x%0h ",pkt_str,this.io_commits_info_5_debug_pdest);
    pkt_str = $sformatf("%sio_commits_info_5_debug_otherPdest_0 = 0x%0h ",pkt_str,this.io_commits_info_5_debug_otherPdest_0);
    pkt_str = $sformatf("%sio_commits_info_5_debug_otherPdest_1 = 0x%0h ",pkt_str,this.io_commits_info_5_debug_otherPdest_1);
    pkt_str = $sformatf("%sio_commits_info_5_debug_otherPdest_2 = 0x%0h ",pkt_str,this.io_commits_info_5_debug_otherPdest_2);
    pkt_str = $sformatf("%sio_commits_info_5_debug_otherPdest_3 = 0x%0h ",pkt_str,this.io_commits_info_5_debug_otherPdest_3);
    pkt_str = $sformatf("%sio_commits_info_5_debug_otherPdest_4 = 0x%0h ",pkt_str,this.io_commits_info_5_debug_otherPdest_4);
    pkt_str = $sformatf("%sio_commits_info_5_debug_otherPdest_5 = 0x%0h ",pkt_str,this.io_commits_info_5_debug_otherPdest_5);
    pkt_str = $sformatf("%sio_commits_info_5_debug_otherPdest_6 = 0x%0h ",pkt_str,this.io_commits_info_5_debug_otherPdest_6);
    pkt_str = $sformatf("%sio_commits_info_5_debug_fuType = 0x%0h ",pkt_str,this.io_commits_info_5_debug_fuType);
    pkt_str = $sformatf("%sio_commits_info_5_dirtyFs = 0x%0h ",pkt_str,this.io_commits_info_5_dirtyFs);
    pkt_str = $sformatf("%sio_commits_info_5_dirtyVs = 0x%0h ",pkt_str,this.io_commits_info_5_dirtyVs);
    pkt_str = $sformatf("%sio_commits_info_6_walk_v = 0x%0h ",pkt_str,this.io_commits_info_6_walk_v);
    pkt_str = $sformatf("%sio_commits_info_6_commit_v = 0x%0h ",pkt_str,this.io_commits_info_6_commit_v);
    pkt_str = $sformatf("%sio_commits_info_6_commit_w = 0x%0h ",pkt_str,this.io_commits_info_6_commit_w);
    pkt_str = $sformatf("%sio_commits_info_6_realDestSize = 0x%0h ",pkt_str,this.io_commits_info_6_realDestSize);
    pkt_str = $sformatf("%sio_commits_info_6_interrupt_safe = 0x%0h ",pkt_str,this.io_commits_info_6_interrupt_safe);
    pkt_str = $sformatf("%sio_commits_info_6_wflags = 0x%0h ",pkt_str,this.io_commits_info_6_wflags);
    pkt_str = $sformatf("%sio_commits_info_6_fflags = 0x%0h ",pkt_str,this.io_commits_info_6_fflags);
    pkt_str = $sformatf("%sio_commits_info_6_vxsat = 0x%0h ",pkt_str,this.io_commits_info_6_vxsat);
    pkt_str = $sformatf("%sio_commits_info_6_isRVC = 0x%0h ",pkt_str,this.io_commits_info_6_isRVC);
    pkt_str = $sformatf("%sio_commits_info_6_isVset = 0x%0h ",pkt_str,this.io_commits_info_6_isVset);
    pkt_str = $sformatf("%sio_commits_info_6_isHls = 0x%0h ",pkt_str,this.io_commits_info_6_isHls);
    pkt_str = $sformatf("%sio_commits_info_6_isVls = 0x%0h ",pkt_str,this.io_commits_info_6_isVls);
    pkt_str = $sformatf("%sio_commits_info_6_vls = 0x%0h ",pkt_str,this.io_commits_info_6_vls);
    pkt_str = $sformatf("%sio_commits_info_6_mmio = 0x%0h ",pkt_str,this.io_commits_info_6_mmio);
    pkt_str = $sformatf("%sio_commits_info_6_commitType = 0x%0h ",pkt_str,this.io_commits_info_6_commitType);
    pkt_str = $sformatf("%sio_commits_info_6_ftqIdx_flag = 0x%0h ",pkt_str,this.io_commits_info_6_ftqIdx_flag);
    pkt_str = $sformatf("%sio_commits_info_6_ftqIdx_value = 0x%0h ",pkt_str,this.io_commits_info_6_ftqIdx_value);
    pkt_str = $sformatf("%sio_commits_info_6_ftqOffset = 0x%0h ",pkt_str,this.io_commits_info_6_ftqOffset);
    pkt_str = $sformatf("%sio_commits_info_6_instrSize = 0x%0h ",pkt_str,this.io_commits_info_6_instrSize);
    pkt_str = $sformatf("%sio_commits_info_6_fpWen = 0x%0h ",pkt_str,this.io_commits_info_6_fpWen);
    pkt_str = $sformatf("%sio_commits_info_6_rfWen = 0x%0h ",pkt_str,this.io_commits_info_6_rfWen);
    pkt_str = $sformatf("%sio_commits_info_6_needFlush = 0x%0h ",pkt_str,this.io_commits_info_6_needFlush);
    pkt_str = $sformatf("%sio_commits_info_6_traceBlockInPipe_itype = 0x%0h ",pkt_str,this.io_commits_info_6_traceBlockInPipe_itype);
    pkt_str = $sformatf("%sio_commits_info_6_traceBlockInPipe_iretire = 0x%0h ",pkt_str,this.io_commits_info_6_traceBlockInPipe_iretire);
    pkt_str = $sformatf("%sio_commits_info_6_traceBlockInPipe_ilastsize = 0x%0h ",pkt_str,this.io_commits_info_6_traceBlockInPipe_ilastsize);
    pkt_str = $sformatf("%sio_commits_info_6_debug_pc = 0x%0h ",pkt_str,this.io_commits_info_6_debug_pc);
    pkt_str = $sformatf("%sio_commits_info_6_debug_instr = 0x%0h ",pkt_str,this.io_commits_info_6_debug_instr);
    pkt_str = $sformatf("%sio_commits_info_6_debug_ldest = 0x%0h ",pkt_str,this.io_commits_info_6_debug_ldest);
    pkt_str = $sformatf("%sio_commits_info_6_debug_pdest = 0x%0h ",pkt_str,this.io_commits_info_6_debug_pdest);
    pkt_str = $sformatf("%sio_commits_info_6_debug_otherPdest_0 = 0x%0h ",pkt_str,this.io_commits_info_6_debug_otherPdest_0);
    pkt_str = $sformatf("%sio_commits_info_6_debug_otherPdest_1 = 0x%0h ",pkt_str,this.io_commits_info_6_debug_otherPdest_1);
    pkt_str = $sformatf("%sio_commits_info_6_debug_otherPdest_2 = 0x%0h ",pkt_str,this.io_commits_info_6_debug_otherPdest_2);
    pkt_str = $sformatf("%sio_commits_info_6_debug_otherPdest_3 = 0x%0h ",pkt_str,this.io_commits_info_6_debug_otherPdest_3);
    pkt_str = $sformatf("%sio_commits_info_6_debug_otherPdest_4 = 0x%0h ",pkt_str,this.io_commits_info_6_debug_otherPdest_4);
    pkt_str = $sformatf("%sio_commits_info_6_debug_otherPdest_5 = 0x%0h ",pkt_str,this.io_commits_info_6_debug_otherPdest_5);
    pkt_str = $sformatf("%sio_commits_info_6_debug_otherPdest_6 = 0x%0h ",pkt_str,this.io_commits_info_6_debug_otherPdest_6);
    pkt_str = $sformatf("%sio_commits_info_6_debug_fuType = 0x%0h ",pkt_str,this.io_commits_info_6_debug_fuType);
    pkt_str = $sformatf("%sio_commits_info_6_dirtyFs = 0x%0h ",pkt_str,this.io_commits_info_6_dirtyFs);
    pkt_str = $sformatf("%sio_commits_info_6_dirtyVs = 0x%0h ",pkt_str,this.io_commits_info_6_dirtyVs);
    pkt_str = $sformatf("%sio_commits_info_7_walk_v = 0x%0h ",pkt_str,this.io_commits_info_7_walk_v);
    pkt_str = $sformatf("%sio_commits_info_7_commit_v = 0x%0h ",pkt_str,this.io_commits_info_7_commit_v);
    pkt_str = $sformatf("%sio_commits_info_7_commit_w = 0x%0h ",pkt_str,this.io_commits_info_7_commit_w);
    pkt_str = $sformatf("%sio_commits_info_7_realDestSize = 0x%0h ",pkt_str,this.io_commits_info_7_realDestSize);
    pkt_str = $sformatf("%sio_commits_info_7_interrupt_safe = 0x%0h ",pkt_str,this.io_commits_info_7_interrupt_safe);
    pkt_str = $sformatf("%sio_commits_info_7_wflags = 0x%0h ",pkt_str,this.io_commits_info_7_wflags);
    pkt_str = $sformatf("%sio_commits_info_7_fflags = 0x%0h ",pkt_str,this.io_commits_info_7_fflags);
    pkt_str = $sformatf("%sio_commits_info_7_vxsat = 0x%0h ",pkt_str,this.io_commits_info_7_vxsat);
    pkt_str = $sformatf("%sio_commits_info_7_isRVC = 0x%0h ",pkt_str,this.io_commits_info_7_isRVC);
    pkt_str = $sformatf("%sio_commits_info_7_isVset = 0x%0h ",pkt_str,this.io_commits_info_7_isVset);
    pkt_str = $sformatf("%sio_commits_info_7_isHls = 0x%0h ",pkt_str,this.io_commits_info_7_isHls);
    pkt_str = $sformatf("%sio_commits_info_7_isVls = 0x%0h ",pkt_str,this.io_commits_info_7_isVls);
    pkt_str = $sformatf("%sio_commits_info_7_vls = 0x%0h ",pkt_str,this.io_commits_info_7_vls);
    pkt_str = $sformatf("%sio_commits_info_7_mmio = 0x%0h ",pkt_str,this.io_commits_info_7_mmio);
    pkt_str = $sformatf("%sio_commits_info_7_commitType = 0x%0h ",pkt_str,this.io_commits_info_7_commitType);
    pkt_str = $sformatf("%sio_commits_info_7_ftqIdx_flag = 0x%0h ",pkt_str,this.io_commits_info_7_ftqIdx_flag);
    pkt_str = $sformatf("%sio_commits_info_7_ftqIdx_value = 0x%0h ",pkt_str,this.io_commits_info_7_ftqIdx_value);
    pkt_str = $sformatf("%sio_commits_info_7_ftqOffset = 0x%0h ",pkt_str,this.io_commits_info_7_ftqOffset);
    pkt_str = $sformatf("%sio_commits_info_7_instrSize = 0x%0h ",pkt_str,this.io_commits_info_7_instrSize);
    pkt_str = $sformatf("%sio_commits_info_7_fpWen = 0x%0h ",pkt_str,this.io_commits_info_7_fpWen);
    pkt_str = $sformatf("%sio_commits_info_7_rfWen = 0x%0h ",pkt_str,this.io_commits_info_7_rfWen);
    pkt_str = $sformatf("%sio_commits_info_7_needFlush = 0x%0h ",pkt_str,this.io_commits_info_7_needFlush);
    pkt_str = $sformatf("%sio_commits_info_7_traceBlockInPipe_itype = 0x%0h ",pkt_str,this.io_commits_info_7_traceBlockInPipe_itype);
    pkt_str = $sformatf("%sio_commits_info_7_traceBlockInPipe_iretire = 0x%0h ",pkt_str,this.io_commits_info_7_traceBlockInPipe_iretire);
    pkt_str = $sformatf("%sio_commits_info_7_traceBlockInPipe_ilastsize = 0x%0h ",pkt_str,this.io_commits_info_7_traceBlockInPipe_ilastsize);
    pkt_str = $sformatf("%sio_commits_info_7_debug_pc = 0x%0h ",pkt_str,this.io_commits_info_7_debug_pc);
    pkt_str = $sformatf("%sio_commits_info_7_debug_instr = 0x%0h ",pkt_str,this.io_commits_info_7_debug_instr);
    pkt_str = $sformatf("%sio_commits_info_7_debug_ldest = 0x%0h ",pkt_str,this.io_commits_info_7_debug_ldest);
    pkt_str = $sformatf("%sio_commits_info_7_debug_pdest = 0x%0h ",pkt_str,this.io_commits_info_7_debug_pdest);
    pkt_str = $sformatf("%sio_commits_info_7_debug_otherPdest_0 = 0x%0h ",pkt_str,this.io_commits_info_7_debug_otherPdest_0);
    pkt_str = $sformatf("%sio_commits_info_7_debug_otherPdest_1 = 0x%0h ",pkt_str,this.io_commits_info_7_debug_otherPdest_1);
    pkt_str = $sformatf("%sio_commits_info_7_debug_otherPdest_2 = 0x%0h ",pkt_str,this.io_commits_info_7_debug_otherPdest_2);
    pkt_str = $sformatf("%sio_commits_info_7_debug_otherPdest_3 = 0x%0h ",pkt_str,this.io_commits_info_7_debug_otherPdest_3);
    pkt_str = $sformatf("%sio_commits_info_7_debug_otherPdest_4 = 0x%0h ",pkt_str,this.io_commits_info_7_debug_otherPdest_4);
    pkt_str = $sformatf("%sio_commits_info_7_debug_otherPdest_5 = 0x%0h ",pkt_str,this.io_commits_info_7_debug_otherPdest_5);
    pkt_str = $sformatf("%sio_commits_info_7_debug_otherPdest_6 = 0x%0h ",pkt_str,this.io_commits_info_7_debug_otherPdest_6);
    pkt_str = $sformatf("%sio_commits_info_7_debug_fuType = 0x%0h ",pkt_str,this.io_commits_info_7_debug_fuType);
    pkt_str = $sformatf("%sio_commits_info_7_dirtyFs = 0x%0h ",pkt_str,this.io_commits_info_7_dirtyFs);
    pkt_str = $sformatf("%sio_commits_info_7_dirtyVs = 0x%0h ",pkt_str,this.io_commits_info_7_dirtyVs);
    pkt_str = $sformatf("%sio_commits_robIdx_0_flag = 0x%0h ",pkt_str,this.io_commits_robIdx_0_flag);
    pkt_str = $sformatf("%sio_commits_robIdx_0_value = 0x%0h ",pkt_str,this.io_commits_robIdx_0_value);
    pkt_str = $sformatf("%sio_commits_robIdx_1_flag = 0x%0h ",pkt_str,this.io_commits_robIdx_1_flag);
    pkt_str = $sformatf("%sio_commits_robIdx_1_value = 0x%0h ",pkt_str,this.io_commits_robIdx_1_value);
    pkt_str = $sformatf("%sio_commits_robIdx_2_flag = 0x%0h ",pkt_str,this.io_commits_robIdx_2_flag);
    pkt_str = $sformatf("%sio_commits_robIdx_2_value = 0x%0h ",pkt_str,this.io_commits_robIdx_2_value);
    pkt_str = $sformatf("%sio_commits_robIdx_3_flag = 0x%0h ",pkt_str,this.io_commits_robIdx_3_flag);
    pkt_str = $sformatf("%sio_commits_robIdx_3_value = 0x%0h ",pkt_str,this.io_commits_robIdx_3_value);
    pkt_str = $sformatf("%sio_commits_robIdx_4_flag = 0x%0h ",pkt_str,this.io_commits_robIdx_4_flag);
    pkt_str = $sformatf("%sio_commits_robIdx_4_value = 0x%0h ",pkt_str,this.io_commits_robIdx_4_value);
    pkt_str = $sformatf("%sio_commits_robIdx_5_flag = 0x%0h ",pkt_str,this.io_commits_robIdx_5_flag);
    pkt_str = $sformatf("%sio_commits_robIdx_5_value = 0x%0h ",pkt_str,this.io_commits_robIdx_5_value);
    pkt_str = $sformatf("%sio_commits_robIdx_6_flag = 0x%0h ",pkt_str,this.io_commits_robIdx_6_flag);
    pkt_str = $sformatf("%sio_commits_robIdx_6_value = 0x%0h ",pkt_str,this.io_commits_robIdx_6_value);
    pkt_str = $sformatf("%sio_commits_robIdx_7_flag = 0x%0h ",pkt_str,this.io_commits_robIdx_7_flag);
    pkt_str = $sformatf("%sio_commits_robIdx_7_value = 0x%0h ",pkt_str,this.io_commits_robIdx_7_value);
    pkt_str = $sformatf("%sio_trace_blockCommit = 0x%0h ",pkt_str,this.io_trace_blockCommit);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_0_valid = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_0_valid);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_0_bits_ftqOffset = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_0_bits_ftqOffset);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_1_valid = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_1_valid);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_1_bits_ftqOffset = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_1_bits_ftqOffset);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_2_valid = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_2_valid);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_2_bits_ftqOffset = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_2_bits_ftqOffset);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_3_valid = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_3_valid);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_3_bits_ftqOffset = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_3_bits_ftqOffset);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_4_valid = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_4_valid);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_4_bits_ftqOffset = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_4_bits_ftqOffset);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_5_valid = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_5_valid);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_5_bits_ftqOffset = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_5_bits_ftqOffset);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_6_valid = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_6_valid);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_6_bits_ftqOffset = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_6_bits_ftqOffset);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_7_valid = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_7_valid);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_7_bits_ftqOffset = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_7_bits_ftqOffset);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire);
    pkt_str = $sformatf("%sio_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize = 0x%0h ",pkt_str,this.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize);
    pkt_str = $sformatf("%sio_rabCommits_isCommit = 0x%0h ",pkt_str,this.io_rabCommits_isCommit);
    pkt_str = $sformatf("%sio_rabCommits_commitValid_0 = 0x%0h ",pkt_str,this.io_rabCommits_commitValid_0);
    pkt_str = $sformatf("%sio_rabCommits_commitValid_1 = 0x%0h ",pkt_str,this.io_rabCommits_commitValid_1);
    pkt_str = $sformatf("%sio_rabCommits_commitValid_2 = 0x%0h ",pkt_str,this.io_rabCommits_commitValid_2);
    pkt_str = $sformatf("%sio_rabCommits_commitValid_3 = 0x%0h ",pkt_str,this.io_rabCommits_commitValid_3);
    pkt_str = $sformatf("%sio_rabCommits_commitValid_4 = 0x%0h ",pkt_str,this.io_rabCommits_commitValid_4);
    pkt_str = $sformatf("%sio_rabCommits_commitValid_5 = 0x%0h ",pkt_str,this.io_rabCommits_commitValid_5);
    pkt_str = $sformatf("%sio_rabCommits_isWalk = 0x%0h ",pkt_str,this.io_rabCommits_isWalk);
    pkt_str = $sformatf("%sio_rabCommits_walkValid_0 = 0x%0h ",pkt_str,this.io_rabCommits_walkValid_0);
    pkt_str = $sformatf("%sio_rabCommits_walkValid_1 = 0x%0h ",pkt_str,this.io_rabCommits_walkValid_1);
    pkt_str = $sformatf("%sio_rabCommits_walkValid_2 = 0x%0h ",pkt_str,this.io_rabCommits_walkValid_2);
    pkt_str = $sformatf("%sio_rabCommits_walkValid_3 = 0x%0h ",pkt_str,this.io_rabCommits_walkValid_3);
    pkt_str = $sformatf("%sio_rabCommits_walkValid_4 = 0x%0h ",pkt_str,this.io_rabCommits_walkValid_4);
    pkt_str = $sformatf("%sio_rabCommits_walkValid_5 = 0x%0h ",pkt_str,this.io_rabCommits_walkValid_5);
    pkt_str = $sformatf("%sio_rabCommits_info_0_ldest = 0x%0h ",pkt_str,this.io_rabCommits_info_0_ldest);
    pkt_str = $sformatf("%sio_rabCommits_info_0_pdest = 0x%0h ",pkt_str,this.io_rabCommits_info_0_pdest);
    pkt_str = $sformatf("%sio_rabCommits_info_0_rfWen = 0x%0h ",pkt_str,this.io_rabCommits_info_0_rfWen);
    pkt_str = $sformatf("%sio_rabCommits_info_0_fpWen = 0x%0h ",pkt_str,this.io_rabCommits_info_0_fpWen);
    pkt_str = $sformatf("%sio_rabCommits_info_0_vecWen = 0x%0h ",pkt_str,this.io_rabCommits_info_0_vecWen);
    pkt_str = $sformatf("%sio_rabCommits_info_0_v0Wen = 0x%0h ",pkt_str,this.io_rabCommits_info_0_v0Wen);
    pkt_str = $sformatf("%sio_rabCommits_info_0_vlWen = 0x%0h ",pkt_str,this.io_rabCommits_info_0_vlWen);
    pkt_str = $sformatf("%sio_rabCommits_info_0_isMove = 0x%0h ",pkt_str,this.io_rabCommits_info_0_isMove);
    pkt_str = $sformatf("%sio_rabCommits_info_1_ldest = 0x%0h ",pkt_str,this.io_rabCommits_info_1_ldest);
    pkt_str = $sformatf("%sio_rabCommits_info_1_pdest = 0x%0h ",pkt_str,this.io_rabCommits_info_1_pdest);
    pkt_str = $sformatf("%sio_rabCommits_info_1_rfWen = 0x%0h ",pkt_str,this.io_rabCommits_info_1_rfWen);
    pkt_str = $sformatf("%sio_rabCommits_info_1_fpWen = 0x%0h ",pkt_str,this.io_rabCommits_info_1_fpWen);
    pkt_str = $sformatf("%sio_rabCommits_info_1_vecWen = 0x%0h ",pkt_str,this.io_rabCommits_info_1_vecWen);
    pkt_str = $sformatf("%sio_rabCommits_info_1_v0Wen = 0x%0h ",pkt_str,this.io_rabCommits_info_1_v0Wen);
    pkt_str = $sformatf("%sio_rabCommits_info_1_vlWen = 0x%0h ",pkt_str,this.io_rabCommits_info_1_vlWen);
    pkt_str = $sformatf("%sio_rabCommits_info_1_isMove = 0x%0h ",pkt_str,this.io_rabCommits_info_1_isMove);
    pkt_str = $sformatf("%sio_rabCommits_info_2_ldest = 0x%0h ",pkt_str,this.io_rabCommits_info_2_ldest);
    pkt_str = $sformatf("%sio_rabCommits_info_2_pdest = 0x%0h ",pkt_str,this.io_rabCommits_info_2_pdest);
    pkt_str = $sformatf("%sio_rabCommits_info_2_rfWen = 0x%0h ",pkt_str,this.io_rabCommits_info_2_rfWen);
    pkt_str = $sformatf("%sio_rabCommits_info_2_fpWen = 0x%0h ",pkt_str,this.io_rabCommits_info_2_fpWen);
    pkt_str = $sformatf("%sio_rabCommits_info_2_vecWen = 0x%0h ",pkt_str,this.io_rabCommits_info_2_vecWen);
    pkt_str = $sformatf("%sio_rabCommits_info_2_v0Wen = 0x%0h ",pkt_str,this.io_rabCommits_info_2_v0Wen);
    pkt_str = $sformatf("%sio_rabCommits_info_2_vlWen = 0x%0h ",pkt_str,this.io_rabCommits_info_2_vlWen);
    pkt_str = $sformatf("%sio_rabCommits_info_2_isMove = 0x%0h ",pkt_str,this.io_rabCommits_info_2_isMove);
    pkt_str = $sformatf("%sio_rabCommits_info_3_ldest = 0x%0h ",pkt_str,this.io_rabCommits_info_3_ldest);
    pkt_str = $sformatf("%sio_rabCommits_info_3_pdest = 0x%0h ",pkt_str,this.io_rabCommits_info_3_pdest);
    pkt_str = $sformatf("%sio_rabCommits_info_3_rfWen = 0x%0h ",pkt_str,this.io_rabCommits_info_3_rfWen);
    pkt_str = $sformatf("%sio_rabCommits_info_3_fpWen = 0x%0h ",pkt_str,this.io_rabCommits_info_3_fpWen);
    pkt_str = $sformatf("%sio_rabCommits_info_3_vecWen = 0x%0h ",pkt_str,this.io_rabCommits_info_3_vecWen);
    pkt_str = $sformatf("%sio_rabCommits_info_3_v0Wen = 0x%0h ",pkt_str,this.io_rabCommits_info_3_v0Wen);
    pkt_str = $sformatf("%sio_rabCommits_info_3_vlWen = 0x%0h ",pkt_str,this.io_rabCommits_info_3_vlWen);
    pkt_str = $sformatf("%sio_rabCommits_info_3_isMove = 0x%0h ",pkt_str,this.io_rabCommits_info_3_isMove);
    pkt_str = $sformatf("%sio_rabCommits_info_4_ldest = 0x%0h ",pkt_str,this.io_rabCommits_info_4_ldest);
    pkt_str = $sformatf("%sio_rabCommits_info_4_pdest = 0x%0h ",pkt_str,this.io_rabCommits_info_4_pdest);
    pkt_str = $sformatf("%sio_rabCommits_info_4_rfWen = 0x%0h ",pkt_str,this.io_rabCommits_info_4_rfWen);
    pkt_str = $sformatf("%sio_rabCommits_info_4_fpWen = 0x%0h ",pkt_str,this.io_rabCommits_info_4_fpWen);
    pkt_str = $sformatf("%sio_rabCommits_info_4_vecWen = 0x%0h ",pkt_str,this.io_rabCommits_info_4_vecWen);
    pkt_str = $sformatf("%sio_rabCommits_info_4_v0Wen = 0x%0h ",pkt_str,this.io_rabCommits_info_4_v0Wen);
    pkt_str = $sformatf("%sio_rabCommits_info_4_vlWen = 0x%0h ",pkt_str,this.io_rabCommits_info_4_vlWen);
    pkt_str = $sformatf("%sio_rabCommits_info_4_isMove = 0x%0h ",pkt_str,this.io_rabCommits_info_4_isMove);
    pkt_str = $sformatf("%sio_rabCommits_info_5_ldest = 0x%0h ",pkt_str,this.io_rabCommits_info_5_ldest);
    pkt_str = $sformatf("%sio_rabCommits_info_5_pdest = 0x%0h ",pkt_str,this.io_rabCommits_info_5_pdest);
    pkt_str = $sformatf("%sio_rabCommits_info_5_rfWen = 0x%0h ",pkt_str,this.io_rabCommits_info_5_rfWen);
    pkt_str = $sformatf("%sio_rabCommits_info_5_fpWen = 0x%0h ",pkt_str,this.io_rabCommits_info_5_fpWen);
    pkt_str = $sformatf("%sio_rabCommits_info_5_vecWen = 0x%0h ",pkt_str,this.io_rabCommits_info_5_vecWen);
    pkt_str = $sformatf("%sio_rabCommits_info_5_v0Wen = 0x%0h ",pkt_str,this.io_rabCommits_info_5_v0Wen);
    pkt_str = $sformatf("%sio_rabCommits_info_5_vlWen = 0x%0h ",pkt_str,this.io_rabCommits_info_5_vlWen);
    pkt_str = $sformatf("%sio_rabCommits_info_5_isMove = 0x%0h ",pkt_str,this.io_rabCommits_info_5_isMove);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_0 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_0);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_1 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_1);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_2 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_2);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_3 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_3);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_4 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_4);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_5 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_5);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_6 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_6);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_7 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_7);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_8 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_8);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_9 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_9);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_10 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_10);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_11 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_11);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_12 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_12);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_13 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_13);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_14 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_14);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_15 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_15);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_16 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_16);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_17 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_17);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_18 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_18);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_19 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_19);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_20 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_20);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_21 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_21);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_22 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_22);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_23 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_23);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_24 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_24);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_25 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_25);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_26 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_26);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_27 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_27);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_28 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_28);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_29 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_29);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_30 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_30);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_31 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_31);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_32 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_32);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_33 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_33);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_34 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_34);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_35 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_35);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_36 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_36);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_37 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_37);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_38 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_38);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_39 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_39);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_40 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_40);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_41 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_41);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_42 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_42);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_43 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_43);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_44 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_44);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_45 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_45);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_46 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_46);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_47 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_47);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_48 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_48);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_49 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_49);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_50 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_50);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_51 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_51);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_52 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_52);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_53 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_53);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_54 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_54);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_55 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_55);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_56 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_56);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_57 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_57);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_58 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_58);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_59 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_59);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_60 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_60);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_61 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_61);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_62 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_62);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_63 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_63);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_64 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_64);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_65 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_65);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_66 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_66);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_67 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_67);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_68 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_68);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_69 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_69);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_70 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_70);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_71 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_71);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_72 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_72);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_73 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_73);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_74 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_74);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_75 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_75);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_76 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_76);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_77 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_77);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_78 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_78);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_79 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_79);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_80 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_80);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_81 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_81);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_82 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_82);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_83 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_83);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_84 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_84);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_85 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_85);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_86 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_86);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_87 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_87);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_88 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_88);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_89 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_89);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_90 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_90);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_91 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_91);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_92 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_92);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_93 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_93);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_94 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_94);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_95 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_95);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_96 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_96);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_97 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_97);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_98 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_98);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_99 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_99);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_100 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_100);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_101 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_101);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_102 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_102);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_103 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_103);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_104 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_104);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_105 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_105);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_106 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_106);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_107 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_107);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_108 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_108);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_109 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_109);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_110 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_110);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_111 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_111);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_112 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_112);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_113 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_113);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_114 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_114);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_115 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_115);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_116 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_116);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_117 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_117);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_118 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_118);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_119 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_119);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_120 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_120);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_121 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_121);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_122 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_122);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_123 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_123);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_124 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_124);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_125 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_125);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_126 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_126);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_127 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_127);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_128 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_128);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_129 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_129);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_130 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_130);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_131 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_131);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_132 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_132);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_133 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_133);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_134 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_134);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_135 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_135);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_136 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_136);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_137 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_137);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_138 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_138);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_139 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_139);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_140 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_140);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_141 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_141);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_142 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_142);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_143 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_143);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_144 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_144);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_145 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_145);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_146 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_146);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_147 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_147);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_148 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_148);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_149 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_149);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_150 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_150);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_151 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_151);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_152 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_152);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_153 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_153);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_154 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_154);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_155 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_155);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_156 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_156);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_157 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_157);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_158 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_158);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_159 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_159);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_160 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_160);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_161 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_161);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_162 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_162);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_163 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_163);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_164 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_164);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_165 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_165);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_166 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_166);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_167 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_167);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_168 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_168);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_169 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_169);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_170 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_170);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_171 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_171);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_172 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_172);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_173 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_173);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_174 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_174);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_175 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_175);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_176 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_176);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_177 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_177);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_178 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_178);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_179 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_179);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_180 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_180);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_181 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_181);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_182 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_182);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_183 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_183);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_184 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_184);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_185 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_185);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_186 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_186);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_187 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_187);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_188 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_188);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_189 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_189);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_190 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_190);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_191 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_191);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_192 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_192);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_193 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_193);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_194 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_194);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_195 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_195);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_196 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_196);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_197 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_197);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_198 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_198);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_199 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_199);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_200 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_200);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_201 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_201);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_202 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_202);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_203 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_203);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_204 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_204);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_205 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_205);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_206 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_206);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_207 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_207);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_208 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_208);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_209 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_209);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_210 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_210);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_211 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_211);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_212 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_212);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_213 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_213);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_214 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_214);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_215 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_215);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_216 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_216);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_217 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_217);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_218 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_218);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_219 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_219);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_220 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_220);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_221 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_221);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_222 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_222);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_223 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_223);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_224 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_224);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_225 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_225);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_226 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_226);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_227 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_227);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_228 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_228);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_229 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_229);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_230 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_230);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_231 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_231);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_232 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_232);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_233 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_233);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_234 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_234);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_235 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_235);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_236 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_236);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_237 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_237);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_238 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_238);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_239 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_239);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_240 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_240);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_241 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_241);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_242 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_242);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_243 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_243);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_244 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_244);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_245 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_245);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_246 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_246);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_247 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_247);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_248 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_248);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_249 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_249);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_250 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_250);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_251 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_251);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_252 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_252);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_253 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_253);
    pkt_str = $sformatf("%sio_diffCommits_commitValid_254 = 0x%0h ",pkt_str,this.io_diffCommits_commitValid_254);
    pkt_str = $sformatf("%sio_diffCommits_info_0_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_0_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_0_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_0_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_0_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_0_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_0_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_0_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_0_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_0_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_0_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_0_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_0_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_0_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_1_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_1_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_1_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_1_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_1_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_1_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_1_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_1_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_1_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_1_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_1_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_1_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_1_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_1_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_2_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_2_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_2_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_2_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_2_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_2_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_2_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_2_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_2_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_2_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_2_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_2_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_2_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_2_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_3_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_3_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_3_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_3_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_3_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_3_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_3_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_3_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_3_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_3_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_3_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_3_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_3_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_3_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_4_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_4_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_4_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_4_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_4_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_4_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_4_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_4_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_4_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_4_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_4_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_4_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_4_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_4_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_5_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_5_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_5_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_5_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_5_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_5_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_5_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_5_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_5_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_5_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_5_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_5_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_5_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_5_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_6_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_6_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_6_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_6_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_6_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_6_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_6_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_6_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_6_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_6_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_6_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_6_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_6_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_6_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_7_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_7_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_7_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_7_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_7_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_7_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_7_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_7_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_7_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_7_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_7_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_7_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_7_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_7_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_8_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_8_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_8_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_8_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_8_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_8_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_8_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_8_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_8_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_8_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_8_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_8_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_8_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_8_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_9_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_9_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_9_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_9_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_9_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_9_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_9_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_9_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_9_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_9_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_9_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_9_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_9_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_9_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_10_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_10_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_10_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_10_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_10_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_10_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_10_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_10_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_10_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_10_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_10_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_10_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_10_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_10_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_11_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_11_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_11_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_11_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_11_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_11_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_11_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_11_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_11_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_11_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_11_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_11_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_11_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_11_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_12_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_12_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_12_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_12_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_12_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_12_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_12_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_12_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_12_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_12_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_12_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_12_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_12_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_12_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_13_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_13_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_13_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_13_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_13_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_13_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_13_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_13_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_13_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_13_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_13_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_13_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_13_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_13_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_14_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_14_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_14_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_14_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_14_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_14_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_14_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_14_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_14_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_14_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_14_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_14_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_14_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_14_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_15_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_15_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_15_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_15_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_15_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_15_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_15_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_15_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_15_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_15_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_15_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_15_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_15_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_15_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_16_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_16_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_16_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_16_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_16_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_16_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_16_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_16_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_16_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_16_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_16_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_16_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_16_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_16_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_17_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_17_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_17_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_17_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_17_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_17_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_17_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_17_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_17_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_17_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_17_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_17_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_17_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_17_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_18_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_18_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_18_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_18_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_18_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_18_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_18_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_18_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_18_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_18_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_18_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_18_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_18_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_18_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_19_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_19_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_19_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_19_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_19_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_19_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_19_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_19_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_19_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_19_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_19_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_19_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_19_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_19_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_20_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_20_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_20_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_20_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_20_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_20_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_20_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_20_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_20_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_20_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_20_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_20_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_20_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_20_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_21_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_21_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_21_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_21_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_21_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_21_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_21_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_21_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_21_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_21_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_21_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_21_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_21_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_21_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_22_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_22_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_22_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_22_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_22_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_22_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_22_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_22_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_22_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_22_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_22_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_22_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_22_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_22_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_23_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_23_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_23_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_23_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_23_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_23_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_23_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_23_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_23_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_23_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_23_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_23_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_23_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_23_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_24_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_24_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_24_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_24_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_24_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_24_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_24_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_24_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_24_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_24_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_24_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_24_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_24_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_24_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_25_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_25_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_25_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_25_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_25_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_25_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_25_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_25_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_25_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_25_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_25_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_25_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_25_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_25_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_26_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_26_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_26_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_26_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_26_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_26_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_26_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_26_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_26_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_26_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_26_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_26_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_26_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_26_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_27_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_27_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_27_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_27_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_27_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_27_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_27_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_27_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_27_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_27_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_27_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_27_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_27_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_27_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_28_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_28_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_28_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_28_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_28_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_28_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_28_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_28_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_28_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_28_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_28_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_28_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_28_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_28_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_29_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_29_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_29_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_29_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_29_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_29_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_29_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_29_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_29_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_29_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_29_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_29_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_29_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_29_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_30_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_30_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_30_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_30_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_30_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_30_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_30_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_30_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_30_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_30_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_30_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_30_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_30_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_30_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_31_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_31_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_31_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_31_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_31_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_31_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_31_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_31_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_31_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_31_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_31_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_31_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_31_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_31_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_32_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_32_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_32_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_32_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_32_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_32_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_32_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_32_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_32_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_32_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_32_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_32_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_32_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_32_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_33_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_33_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_33_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_33_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_33_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_33_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_33_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_33_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_33_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_33_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_33_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_33_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_33_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_33_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_34_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_34_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_34_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_34_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_34_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_34_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_34_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_34_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_34_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_34_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_34_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_34_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_34_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_34_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_35_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_35_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_35_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_35_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_35_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_35_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_35_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_35_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_35_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_35_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_35_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_35_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_35_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_35_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_36_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_36_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_36_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_36_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_36_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_36_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_36_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_36_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_36_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_36_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_36_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_36_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_36_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_36_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_37_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_37_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_37_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_37_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_37_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_37_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_37_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_37_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_37_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_37_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_37_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_37_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_37_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_37_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_38_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_38_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_38_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_38_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_38_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_38_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_38_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_38_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_38_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_38_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_38_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_38_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_38_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_38_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_39_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_39_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_39_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_39_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_39_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_39_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_39_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_39_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_39_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_39_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_39_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_39_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_39_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_39_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_40_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_40_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_40_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_40_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_40_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_40_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_40_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_40_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_40_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_40_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_40_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_40_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_40_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_40_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_41_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_41_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_41_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_41_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_41_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_41_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_41_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_41_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_41_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_41_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_41_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_41_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_41_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_41_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_42_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_42_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_42_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_42_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_42_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_42_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_42_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_42_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_42_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_42_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_42_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_42_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_42_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_42_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_43_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_43_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_43_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_43_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_43_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_43_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_43_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_43_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_43_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_43_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_43_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_43_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_43_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_43_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_44_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_44_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_44_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_44_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_44_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_44_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_44_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_44_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_44_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_44_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_44_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_44_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_44_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_44_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_45_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_45_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_45_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_45_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_45_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_45_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_45_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_45_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_45_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_45_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_45_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_45_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_45_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_45_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_46_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_46_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_46_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_46_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_46_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_46_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_46_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_46_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_46_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_46_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_46_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_46_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_46_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_46_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_47_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_47_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_47_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_47_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_47_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_47_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_47_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_47_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_47_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_47_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_47_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_47_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_47_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_47_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_48_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_48_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_48_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_48_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_48_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_48_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_48_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_48_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_48_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_48_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_48_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_48_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_48_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_48_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_49_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_49_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_49_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_49_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_49_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_49_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_49_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_49_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_49_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_49_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_49_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_49_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_49_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_49_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_50_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_50_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_50_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_50_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_50_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_50_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_50_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_50_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_50_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_50_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_50_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_50_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_50_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_50_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_51_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_51_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_51_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_51_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_51_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_51_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_51_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_51_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_51_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_51_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_51_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_51_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_51_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_51_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_52_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_52_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_52_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_52_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_52_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_52_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_52_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_52_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_52_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_52_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_52_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_52_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_52_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_52_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_53_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_53_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_53_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_53_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_53_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_53_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_53_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_53_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_53_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_53_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_53_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_53_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_53_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_53_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_54_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_54_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_54_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_54_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_54_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_54_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_54_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_54_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_54_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_54_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_54_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_54_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_54_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_54_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_55_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_55_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_55_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_55_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_55_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_55_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_55_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_55_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_55_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_55_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_55_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_55_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_55_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_55_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_56_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_56_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_56_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_56_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_56_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_56_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_56_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_56_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_56_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_56_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_56_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_56_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_56_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_56_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_57_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_57_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_57_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_57_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_57_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_57_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_57_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_57_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_57_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_57_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_57_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_57_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_57_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_57_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_58_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_58_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_58_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_58_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_58_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_58_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_58_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_58_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_58_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_58_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_58_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_58_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_58_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_58_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_59_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_59_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_59_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_59_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_59_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_59_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_59_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_59_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_59_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_59_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_59_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_59_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_59_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_59_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_60_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_60_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_60_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_60_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_60_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_60_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_60_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_60_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_60_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_60_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_60_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_60_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_60_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_60_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_61_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_61_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_61_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_61_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_61_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_61_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_61_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_61_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_61_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_61_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_61_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_61_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_61_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_61_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_62_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_62_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_62_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_62_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_62_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_62_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_62_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_62_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_62_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_62_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_62_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_62_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_62_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_62_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_63_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_63_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_63_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_63_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_63_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_63_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_63_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_63_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_63_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_63_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_63_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_63_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_63_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_63_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_64_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_64_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_64_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_64_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_64_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_64_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_64_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_64_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_64_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_64_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_64_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_64_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_64_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_64_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_65_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_65_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_65_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_65_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_65_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_65_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_65_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_65_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_65_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_65_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_65_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_65_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_65_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_65_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_66_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_66_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_66_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_66_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_66_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_66_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_66_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_66_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_66_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_66_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_66_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_66_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_66_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_66_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_67_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_67_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_67_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_67_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_67_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_67_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_67_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_67_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_67_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_67_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_67_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_67_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_67_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_67_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_68_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_68_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_68_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_68_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_68_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_68_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_68_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_68_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_68_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_68_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_68_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_68_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_68_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_68_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_69_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_69_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_69_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_69_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_69_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_69_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_69_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_69_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_69_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_69_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_69_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_69_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_69_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_69_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_70_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_70_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_70_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_70_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_70_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_70_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_70_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_70_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_70_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_70_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_70_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_70_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_70_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_70_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_71_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_71_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_71_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_71_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_71_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_71_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_71_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_71_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_71_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_71_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_71_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_71_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_71_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_71_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_72_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_72_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_72_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_72_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_72_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_72_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_72_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_72_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_72_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_72_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_72_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_72_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_72_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_72_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_73_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_73_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_73_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_73_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_73_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_73_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_73_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_73_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_73_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_73_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_73_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_73_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_73_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_73_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_74_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_74_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_74_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_74_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_74_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_74_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_74_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_74_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_74_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_74_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_74_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_74_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_74_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_74_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_75_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_75_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_75_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_75_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_75_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_75_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_75_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_75_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_75_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_75_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_75_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_75_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_75_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_75_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_76_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_76_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_76_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_76_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_76_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_76_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_76_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_76_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_76_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_76_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_76_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_76_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_76_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_76_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_77_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_77_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_77_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_77_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_77_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_77_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_77_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_77_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_77_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_77_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_77_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_77_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_77_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_77_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_78_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_78_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_78_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_78_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_78_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_78_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_78_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_78_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_78_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_78_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_78_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_78_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_78_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_78_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_79_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_79_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_79_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_79_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_79_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_79_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_79_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_79_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_79_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_79_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_79_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_79_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_79_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_79_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_80_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_80_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_80_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_80_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_80_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_80_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_80_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_80_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_80_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_80_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_80_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_80_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_80_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_80_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_81_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_81_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_81_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_81_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_81_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_81_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_81_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_81_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_81_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_81_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_81_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_81_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_81_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_81_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_82_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_82_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_82_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_82_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_82_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_82_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_82_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_82_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_82_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_82_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_82_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_82_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_82_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_82_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_83_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_83_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_83_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_83_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_83_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_83_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_83_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_83_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_83_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_83_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_83_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_83_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_83_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_83_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_84_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_84_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_84_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_84_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_84_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_84_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_84_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_84_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_84_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_84_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_84_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_84_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_84_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_84_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_85_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_85_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_85_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_85_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_85_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_85_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_85_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_85_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_85_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_85_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_85_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_85_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_85_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_85_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_86_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_86_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_86_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_86_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_86_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_86_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_86_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_86_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_86_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_86_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_86_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_86_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_86_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_86_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_87_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_87_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_87_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_87_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_87_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_87_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_87_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_87_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_87_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_87_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_87_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_87_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_87_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_87_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_88_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_88_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_88_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_88_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_88_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_88_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_88_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_88_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_88_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_88_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_88_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_88_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_88_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_88_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_89_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_89_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_89_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_89_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_89_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_89_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_89_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_89_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_89_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_89_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_89_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_89_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_89_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_89_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_90_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_90_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_90_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_90_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_90_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_90_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_90_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_90_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_90_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_90_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_90_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_90_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_90_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_90_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_91_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_91_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_91_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_91_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_91_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_91_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_91_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_91_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_91_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_91_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_91_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_91_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_91_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_91_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_92_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_92_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_92_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_92_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_92_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_92_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_92_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_92_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_92_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_92_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_92_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_92_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_92_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_92_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_93_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_93_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_93_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_93_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_93_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_93_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_93_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_93_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_93_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_93_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_93_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_93_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_93_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_93_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_94_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_94_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_94_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_94_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_94_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_94_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_94_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_94_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_94_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_94_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_94_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_94_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_94_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_94_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_95_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_95_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_95_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_95_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_95_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_95_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_95_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_95_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_95_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_95_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_95_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_95_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_95_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_95_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_96_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_96_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_96_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_96_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_96_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_96_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_96_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_96_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_96_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_96_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_96_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_96_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_96_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_96_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_97_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_97_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_97_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_97_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_97_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_97_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_97_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_97_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_97_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_97_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_97_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_97_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_97_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_97_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_98_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_98_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_98_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_98_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_98_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_98_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_98_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_98_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_98_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_98_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_98_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_98_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_98_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_98_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_99_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_99_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_99_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_99_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_99_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_99_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_99_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_99_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_99_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_99_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_99_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_99_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_99_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_99_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_100_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_100_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_100_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_100_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_100_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_100_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_100_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_100_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_100_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_100_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_100_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_100_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_100_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_100_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_101_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_101_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_101_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_101_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_101_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_101_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_101_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_101_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_101_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_101_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_101_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_101_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_101_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_101_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_102_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_102_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_102_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_102_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_102_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_102_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_102_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_102_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_102_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_102_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_102_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_102_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_102_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_102_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_103_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_103_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_103_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_103_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_103_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_103_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_103_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_103_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_103_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_103_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_103_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_103_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_103_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_103_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_104_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_104_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_104_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_104_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_104_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_104_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_104_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_104_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_104_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_104_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_104_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_104_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_104_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_104_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_105_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_105_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_105_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_105_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_105_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_105_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_105_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_105_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_105_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_105_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_105_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_105_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_105_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_105_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_106_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_106_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_106_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_106_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_106_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_106_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_106_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_106_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_106_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_106_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_106_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_106_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_106_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_106_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_107_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_107_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_107_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_107_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_107_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_107_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_107_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_107_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_107_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_107_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_107_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_107_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_107_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_107_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_108_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_108_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_108_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_108_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_108_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_108_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_108_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_108_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_108_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_108_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_108_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_108_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_108_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_108_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_109_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_109_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_109_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_109_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_109_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_109_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_109_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_109_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_109_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_109_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_109_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_109_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_109_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_109_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_110_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_110_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_110_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_110_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_110_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_110_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_110_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_110_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_110_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_110_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_110_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_110_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_110_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_110_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_111_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_111_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_111_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_111_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_111_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_111_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_111_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_111_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_111_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_111_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_111_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_111_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_111_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_111_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_112_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_112_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_112_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_112_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_112_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_112_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_112_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_112_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_112_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_112_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_112_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_112_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_112_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_112_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_113_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_113_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_113_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_113_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_113_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_113_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_113_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_113_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_113_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_113_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_113_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_113_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_113_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_113_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_114_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_114_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_114_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_114_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_114_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_114_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_114_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_114_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_114_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_114_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_114_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_114_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_114_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_114_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_115_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_115_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_115_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_115_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_115_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_115_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_115_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_115_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_115_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_115_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_115_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_115_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_115_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_115_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_116_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_116_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_116_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_116_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_116_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_116_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_116_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_116_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_116_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_116_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_116_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_116_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_116_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_116_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_117_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_117_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_117_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_117_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_117_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_117_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_117_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_117_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_117_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_117_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_117_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_117_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_117_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_117_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_118_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_118_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_118_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_118_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_118_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_118_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_118_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_118_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_118_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_118_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_118_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_118_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_118_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_118_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_119_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_119_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_119_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_119_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_119_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_119_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_119_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_119_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_119_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_119_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_119_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_119_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_119_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_119_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_120_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_120_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_120_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_120_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_120_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_120_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_120_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_120_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_120_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_120_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_120_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_120_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_120_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_120_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_121_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_121_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_121_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_121_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_121_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_121_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_121_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_121_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_121_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_121_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_121_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_121_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_121_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_121_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_122_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_122_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_122_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_122_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_122_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_122_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_122_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_122_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_122_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_122_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_122_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_122_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_122_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_122_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_123_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_123_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_123_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_123_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_123_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_123_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_123_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_123_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_123_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_123_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_123_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_123_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_123_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_123_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_124_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_124_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_124_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_124_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_124_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_124_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_124_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_124_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_124_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_124_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_124_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_124_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_124_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_124_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_125_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_125_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_125_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_125_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_125_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_125_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_125_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_125_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_125_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_125_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_125_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_125_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_125_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_125_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_126_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_126_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_126_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_126_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_126_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_126_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_126_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_126_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_126_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_126_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_126_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_126_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_126_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_126_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_127_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_127_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_127_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_127_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_127_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_127_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_127_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_127_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_127_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_127_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_127_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_127_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_127_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_127_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_128_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_128_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_128_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_128_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_128_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_128_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_128_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_128_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_128_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_128_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_128_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_128_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_128_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_128_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_129_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_129_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_129_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_129_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_129_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_129_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_129_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_129_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_129_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_129_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_129_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_129_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_129_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_129_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_130_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_130_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_130_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_130_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_130_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_130_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_130_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_130_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_130_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_130_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_130_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_130_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_130_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_130_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_131_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_131_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_131_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_131_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_131_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_131_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_131_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_131_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_131_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_131_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_131_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_131_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_131_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_131_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_132_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_132_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_132_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_132_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_132_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_132_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_132_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_132_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_132_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_132_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_132_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_132_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_132_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_132_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_133_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_133_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_133_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_133_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_133_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_133_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_133_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_133_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_133_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_133_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_133_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_133_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_133_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_133_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_134_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_134_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_134_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_134_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_134_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_134_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_134_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_134_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_134_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_134_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_134_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_134_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_134_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_134_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_135_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_135_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_135_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_135_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_135_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_135_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_135_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_135_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_135_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_135_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_135_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_135_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_135_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_135_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_136_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_136_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_136_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_136_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_136_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_136_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_136_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_136_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_136_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_136_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_136_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_136_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_136_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_136_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_137_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_137_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_137_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_137_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_137_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_137_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_137_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_137_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_137_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_137_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_137_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_137_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_137_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_137_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_138_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_138_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_138_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_138_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_138_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_138_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_138_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_138_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_138_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_138_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_138_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_138_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_138_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_138_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_139_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_139_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_139_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_139_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_139_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_139_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_139_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_139_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_139_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_139_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_139_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_139_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_139_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_139_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_140_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_140_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_140_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_140_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_140_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_140_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_140_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_140_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_140_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_140_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_140_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_140_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_140_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_140_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_141_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_141_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_141_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_141_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_141_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_141_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_141_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_141_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_141_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_141_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_141_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_141_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_141_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_141_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_142_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_142_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_142_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_142_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_142_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_142_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_142_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_142_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_142_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_142_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_142_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_142_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_142_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_142_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_143_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_143_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_143_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_143_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_143_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_143_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_143_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_143_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_143_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_143_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_143_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_143_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_143_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_143_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_144_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_144_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_144_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_144_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_144_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_144_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_144_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_144_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_144_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_144_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_144_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_144_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_144_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_144_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_145_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_145_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_145_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_145_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_145_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_145_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_145_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_145_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_145_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_145_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_145_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_145_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_145_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_145_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_146_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_146_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_146_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_146_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_146_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_146_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_146_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_146_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_146_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_146_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_146_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_146_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_146_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_146_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_147_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_147_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_147_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_147_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_147_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_147_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_147_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_147_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_147_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_147_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_147_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_147_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_147_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_147_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_148_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_148_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_148_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_148_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_148_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_148_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_148_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_148_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_148_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_148_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_148_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_148_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_148_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_148_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_149_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_149_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_149_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_149_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_149_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_149_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_149_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_149_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_149_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_149_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_149_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_149_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_149_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_149_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_150_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_150_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_150_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_150_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_150_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_150_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_150_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_150_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_150_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_150_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_150_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_150_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_150_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_150_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_151_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_151_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_151_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_151_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_151_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_151_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_151_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_151_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_151_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_151_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_151_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_151_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_151_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_151_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_152_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_152_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_152_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_152_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_152_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_152_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_152_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_152_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_152_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_152_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_152_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_152_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_152_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_152_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_153_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_153_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_153_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_153_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_153_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_153_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_153_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_153_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_153_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_153_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_153_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_153_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_153_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_153_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_154_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_154_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_154_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_154_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_154_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_154_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_154_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_154_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_154_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_154_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_154_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_154_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_154_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_154_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_155_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_155_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_155_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_155_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_155_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_155_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_155_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_155_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_155_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_155_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_155_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_155_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_155_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_155_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_156_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_156_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_156_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_156_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_156_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_156_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_156_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_156_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_156_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_156_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_156_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_156_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_156_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_156_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_157_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_157_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_157_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_157_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_157_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_157_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_157_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_157_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_157_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_157_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_157_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_157_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_157_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_157_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_158_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_158_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_158_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_158_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_158_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_158_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_158_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_158_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_158_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_158_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_158_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_158_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_158_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_158_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_159_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_159_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_159_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_159_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_159_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_159_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_159_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_159_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_159_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_159_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_159_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_159_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_159_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_159_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_160_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_160_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_160_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_160_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_160_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_160_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_160_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_160_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_160_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_160_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_160_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_160_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_160_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_160_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_161_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_161_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_161_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_161_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_161_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_161_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_161_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_161_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_161_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_161_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_161_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_161_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_161_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_161_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_162_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_162_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_162_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_162_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_162_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_162_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_162_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_162_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_162_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_162_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_162_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_162_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_162_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_162_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_163_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_163_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_163_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_163_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_163_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_163_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_163_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_163_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_163_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_163_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_163_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_163_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_163_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_163_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_164_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_164_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_164_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_164_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_164_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_164_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_164_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_164_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_164_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_164_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_164_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_164_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_164_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_164_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_165_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_165_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_165_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_165_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_165_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_165_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_165_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_165_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_165_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_165_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_165_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_165_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_165_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_165_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_166_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_166_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_166_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_166_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_166_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_166_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_166_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_166_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_166_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_166_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_166_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_166_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_166_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_166_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_167_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_167_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_167_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_167_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_167_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_167_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_167_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_167_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_167_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_167_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_167_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_167_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_167_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_167_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_168_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_168_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_168_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_168_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_168_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_168_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_168_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_168_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_168_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_168_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_168_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_168_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_168_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_168_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_169_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_169_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_169_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_169_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_169_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_169_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_169_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_169_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_169_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_169_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_169_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_169_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_169_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_169_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_170_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_170_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_170_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_170_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_170_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_170_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_170_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_170_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_170_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_170_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_170_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_170_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_170_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_170_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_171_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_171_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_171_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_171_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_171_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_171_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_171_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_171_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_171_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_171_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_171_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_171_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_171_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_171_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_172_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_172_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_172_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_172_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_172_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_172_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_172_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_172_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_172_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_172_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_172_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_172_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_172_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_172_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_173_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_173_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_173_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_173_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_173_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_173_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_173_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_173_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_173_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_173_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_173_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_173_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_173_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_173_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_174_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_174_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_174_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_174_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_174_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_174_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_174_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_174_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_174_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_174_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_174_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_174_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_174_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_174_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_175_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_175_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_175_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_175_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_175_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_175_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_175_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_175_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_175_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_175_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_175_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_175_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_175_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_175_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_176_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_176_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_176_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_176_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_176_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_176_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_176_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_176_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_176_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_176_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_176_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_176_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_176_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_176_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_177_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_177_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_177_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_177_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_177_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_177_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_177_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_177_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_177_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_177_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_177_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_177_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_177_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_177_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_178_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_178_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_178_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_178_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_178_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_178_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_178_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_178_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_178_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_178_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_178_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_178_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_178_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_178_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_179_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_179_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_179_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_179_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_179_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_179_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_179_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_179_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_179_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_179_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_179_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_179_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_179_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_179_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_180_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_180_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_180_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_180_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_180_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_180_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_180_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_180_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_180_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_180_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_180_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_180_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_180_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_180_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_181_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_181_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_181_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_181_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_181_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_181_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_181_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_181_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_181_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_181_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_181_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_181_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_181_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_181_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_182_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_182_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_182_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_182_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_182_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_182_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_182_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_182_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_182_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_182_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_182_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_182_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_182_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_182_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_183_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_183_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_183_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_183_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_183_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_183_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_183_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_183_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_183_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_183_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_183_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_183_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_183_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_183_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_184_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_184_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_184_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_184_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_184_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_184_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_184_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_184_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_184_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_184_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_184_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_184_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_184_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_184_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_185_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_185_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_185_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_185_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_185_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_185_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_185_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_185_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_185_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_185_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_185_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_185_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_185_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_185_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_186_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_186_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_186_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_186_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_186_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_186_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_186_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_186_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_186_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_186_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_186_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_186_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_186_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_186_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_187_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_187_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_187_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_187_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_187_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_187_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_187_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_187_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_187_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_187_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_187_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_187_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_187_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_187_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_188_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_188_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_188_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_188_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_188_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_188_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_188_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_188_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_188_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_188_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_188_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_188_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_188_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_188_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_189_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_189_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_189_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_189_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_189_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_189_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_189_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_189_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_189_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_189_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_189_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_189_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_189_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_189_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_190_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_190_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_190_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_190_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_190_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_190_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_190_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_190_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_190_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_190_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_190_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_190_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_190_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_190_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_191_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_191_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_191_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_191_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_191_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_191_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_191_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_191_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_191_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_191_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_191_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_191_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_191_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_191_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_192_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_192_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_192_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_192_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_192_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_192_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_192_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_192_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_192_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_192_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_192_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_192_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_192_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_192_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_193_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_193_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_193_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_193_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_193_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_193_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_193_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_193_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_193_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_193_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_193_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_193_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_193_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_193_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_194_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_194_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_194_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_194_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_194_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_194_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_194_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_194_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_194_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_194_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_194_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_194_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_194_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_194_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_195_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_195_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_195_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_195_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_195_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_195_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_195_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_195_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_195_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_195_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_195_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_195_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_195_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_195_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_196_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_196_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_196_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_196_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_196_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_196_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_196_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_196_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_196_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_196_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_196_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_196_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_196_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_196_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_197_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_197_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_197_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_197_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_197_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_197_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_197_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_197_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_197_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_197_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_197_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_197_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_197_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_197_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_198_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_198_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_198_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_198_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_198_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_198_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_198_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_198_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_198_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_198_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_198_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_198_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_198_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_198_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_199_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_199_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_199_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_199_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_199_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_199_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_199_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_199_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_199_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_199_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_199_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_199_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_199_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_199_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_200_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_200_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_200_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_200_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_200_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_200_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_200_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_200_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_200_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_200_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_200_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_200_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_200_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_200_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_201_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_201_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_201_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_201_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_201_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_201_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_201_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_201_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_201_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_201_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_201_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_201_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_201_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_201_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_202_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_202_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_202_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_202_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_202_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_202_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_202_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_202_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_202_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_202_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_202_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_202_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_202_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_202_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_203_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_203_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_203_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_203_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_203_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_203_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_203_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_203_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_203_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_203_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_203_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_203_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_203_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_203_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_204_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_204_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_204_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_204_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_204_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_204_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_204_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_204_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_204_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_204_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_204_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_204_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_204_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_204_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_205_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_205_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_205_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_205_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_205_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_205_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_205_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_205_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_205_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_205_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_205_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_205_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_205_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_205_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_206_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_206_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_206_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_206_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_206_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_206_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_206_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_206_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_206_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_206_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_206_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_206_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_206_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_206_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_207_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_207_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_207_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_207_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_207_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_207_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_207_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_207_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_207_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_207_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_207_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_207_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_207_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_207_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_208_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_208_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_208_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_208_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_208_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_208_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_208_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_208_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_208_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_208_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_208_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_208_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_208_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_208_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_209_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_209_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_209_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_209_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_209_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_209_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_209_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_209_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_209_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_209_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_209_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_209_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_209_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_209_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_210_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_210_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_210_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_210_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_210_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_210_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_210_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_210_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_210_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_210_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_210_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_210_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_210_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_210_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_211_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_211_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_211_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_211_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_211_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_211_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_211_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_211_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_211_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_211_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_211_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_211_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_211_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_211_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_212_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_212_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_212_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_212_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_212_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_212_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_212_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_212_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_212_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_212_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_212_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_212_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_212_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_212_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_213_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_213_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_213_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_213_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_213_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_213_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_213_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_213_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_213_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_213_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_213_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_213_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_213_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_213_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_214_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_214_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_214_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_214_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_214_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_214_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_214_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_214_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_214_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_214_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_214_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_214_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_214_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_214_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_215_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_215_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_215_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_215_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_215_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_215_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_215_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_215_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_215_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_215_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_215_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_215_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_215_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_215_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_216_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_216_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_216_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_216_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_216_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_216_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_216_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_216_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_216_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_216_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_216_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_216_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_216_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_216_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_217_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_217_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_217_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_217_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_217_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_217_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_217_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_217_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_217_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_217_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_217_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_217_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_217_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_217_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_218_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_218_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_218_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_218_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_218_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_218_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_218_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_218_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_218_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_218_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_218_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_218_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_218_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_218_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_219_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_219_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_219_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_219_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_219_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_219_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_219_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_219_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_219_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_219_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_219_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_219_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_219_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_219_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_220_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_220_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_220_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_220_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_220_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_220_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_220_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_220_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_220_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_220_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_220_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_220_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_220_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_220_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_221_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_221_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_221_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_221_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_221_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_221_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_221_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_221_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_221_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_221_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_221_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_221_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_221_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_221_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_222_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_222_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_222_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_222_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_222_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_222_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_222_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_222_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_222_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_222_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_222_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_222_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_222_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_222_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_223_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_223_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_223_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_223_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_223_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_223_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_223_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_223_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_223_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_223_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_223_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_223_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_223_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_223_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_224_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_224_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_224_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_224_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_224_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_224_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_224_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_224_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_224_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_224_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_224_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_224_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_224_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_224_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_225_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_225_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_225_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_225_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_225_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_225_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_225_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_225_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_225_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_225_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_225_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_225_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_225_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_225_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_226_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_226_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_226_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_226_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_226_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_226_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_226_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_226_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_226_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_226_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_226_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_226_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_226_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_226_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_227_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_227_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_227_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_227_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_227_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_227_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_227_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_227_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_227_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_227_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_227_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_227_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_227_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_227_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_228_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_228_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_228_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_228_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_228_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_228_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_228_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_228_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_228_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_228_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_228_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_228_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_228_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_228_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_229_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_229_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_229_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_229_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_229_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_229_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_229_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_229_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_229_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_229_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_229_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_229_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_229_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_229_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_230_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_230_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_230_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_230_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_230_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_230_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_230_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_230_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_230_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_230_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_230_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_230_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_230_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_230_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_231_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_231_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_231_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_231_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_231_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_231_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_231_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_231_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_231_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_231_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_231_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_231_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_231_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_231_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_232_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_232_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_232_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_232_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_232_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_232_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_232_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_232_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_232_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_232_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_232_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_232_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_232_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_232_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_233_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_233_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_233_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_233_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_233_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_233_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_233_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_233_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_233_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_233_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_233_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_233_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_233_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_233_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_234_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_234_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_234_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_234_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_234_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_234_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_234_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_234_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_234_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_234_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_234_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_234_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_234_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_234_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_235_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_235_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_235_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_235_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_235_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_235_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_235_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_235_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_235_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_235_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_235_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_235_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_235_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_235_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_236_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_236_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_236_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_236_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_236_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_236_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_236_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_236_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_236_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_236_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_236_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_236_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_236_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_236_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_237_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_237_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_237_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_237_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_237_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_237_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_237_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_237_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_237_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_237_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_237_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_237_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_237_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_237_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_238_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_238_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_238_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_238_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_238_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_238_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_238_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_238_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_238_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_238_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_238_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_238_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_238_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_238_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_239_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_239_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_239_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_239_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_239_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_239_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_239_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_239_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_239_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_239_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_239_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_239_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_239_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_239_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_240_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_240_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_240_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_240_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_240_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_240_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_240_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_240_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_240_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_240_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_240_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_240_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_240_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_240_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_241_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_241_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_241_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_241_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_241_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_241_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_241_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_241_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_241_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_241_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_241_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_241_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_241_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_241_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_242_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_242_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_242_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_242_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_242_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_242_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_242_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_242_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_242_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_242_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_242_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_242_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_242_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_242_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_243_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_243_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_243_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_243_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_243_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_243_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_243_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_243_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_243_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_243_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_243_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_243_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_243_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_243_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_244_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_244_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_244_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_244_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_244_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_244_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_244_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_244_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_244_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_244_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_244_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_244_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_244_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_244_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_245_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_245_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_245_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_245_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_245_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_245_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_245_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_245_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_245_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_245_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_245_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_245_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_245_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_245_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_246_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_246_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_246_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_246_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_246_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_246_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_246_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_246_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_246_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_246_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_246_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_246_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_246_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_246_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_247_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_247_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_247_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_247_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_247_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_247_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_247_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_247_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_247_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_247_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_247_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_247_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_247_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_247_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_248_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_248_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_248_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_248_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_248_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_248_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_248_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_248_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_248_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_248_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_248_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_248_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_248_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_248_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_249_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_249_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_249_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_249_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_249_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_249_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_249_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_249_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_249_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_249_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_249_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_249_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_249_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_249_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_250_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_250_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_250_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_250_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_250_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_250_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_250_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_250_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_250_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_250_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_250_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_250_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_250_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_250_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_251_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_251_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_251_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_251_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_251_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_251_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_251_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_251_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_251_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_251_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_251_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_251_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_251_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_251_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_252_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_252_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_252_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_252_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_252_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_252_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_252_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_252_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_252_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_252_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_252_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_252_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_252_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_252_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_253_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_253_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_253_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_253_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_253_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_253_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_253_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_253_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_253_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_253_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_253_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_253_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_253_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_253_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_254_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_254_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_254_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_254_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_254_rfWen = 0x%0h ",pkt_str,this.io_diffCommits_info_254_rfWen);
    pkt_str = $sformatf("%sio_diffCommits_info_254_fpWen = 0x%0h ",pkt_str,this.io_diffCommits_info_254_fpWen);
    pkt_str = $sformatf("%sio_diffCommits_info_254_vecWen = 0x%0h ",pkt_str,this.io_diffCommits_info_254_vecWen);
    pkt_str = $sformatf("%sio_diffCommits_info_254_v0Wen = 0x%0h ",pkt_str,this.io_diffCommits_info_254_v0Wen);
    pkt_str = $sformatf("%sio_diffCommits_info_254_vlWen = 0x%0h ",pkt_str,this.io_diffCommits_info_254_vlWen);
    pkt_str = $sformatf("%sio_diffCommits_info_255_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_255_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_255_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_255_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_256_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_256_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_256_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_256_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_257_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_257_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_257_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_257_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_258_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_258_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_258_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_258_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_259_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_259_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_259_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_259_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_260_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_260_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_260_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_260_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_261_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_261_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_261_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_261_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_262_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_262_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_262_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_262_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_263_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_263_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_263_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_263_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_264_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_264_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_264_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_264_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_265_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_265_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_265_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_265_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_266_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_266_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_266_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_266_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_267_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_267_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_267_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_267_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_268_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_268_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_268_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_268_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_269_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_269_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_269_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_269_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_270_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_270_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_270_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_270_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_271_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_271_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_271_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_271_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_272_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_272_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_272_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_272_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_273_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_273_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_273_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_273_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_274_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_274_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_274_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_274_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_275_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_275_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_275_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_275_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_276_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_276_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_276_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_276_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_277_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_277_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_277_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_277_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_278_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_278_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_278_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_278_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_279_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_279_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_279_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_279_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_280_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_280_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_280_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_280_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_281_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_281_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_281_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_281_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_282_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_282_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_282_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_282_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_283_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_283_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_283_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_283_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_284_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_284_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_284_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_284_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_285_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_285_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_285_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_285_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_286_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_286_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_286_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_286_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_287_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_287_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_287_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_287_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_288_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_288_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_288_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_288_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_289_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_289_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_289_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_289_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_290_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_290_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_290_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_290_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_291_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_291_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_291_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_291_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_292_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_292_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_292_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_292_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_293_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_293_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_293_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_293_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_294_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_294_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_294_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_294_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_295_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_295_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_295_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_295_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_296_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_296_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_296_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_296_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_297_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_297_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_297_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_297_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_298_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_298_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_298_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_298_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_299_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_299_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_299_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_299_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_300_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_300_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_300_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_300_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_301_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_301_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_301_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_301_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_302_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_302_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_302_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_302_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_303_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_303_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_303_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_303_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_304_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_304_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_304_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_304_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_305_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_305_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_305_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_305_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_306_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_306_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_306_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_306_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_307_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_307_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_307_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_307_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_308_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_308_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_308_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_308_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_309_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_309_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_309_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_309_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_310_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_310_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_310_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_310_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_311_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_311_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_311_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_311_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_312_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_312_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_312_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_312_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_313_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_313_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_313_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_313_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_314_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_314_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_314_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_314_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_315_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_315_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_315_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_315_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_316_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_316_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_316_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_316_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_317_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_317_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_317_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_317_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_318_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_318_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_318_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_318_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_319_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_319_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_319_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_319_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_320_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_320_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_320_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_320_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_321_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_321_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_321_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_321_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_322_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_322_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_322_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_322_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_323_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_323_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_323_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_323_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_324_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_324_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_324_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_324_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_325_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_325_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_325_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_325_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_326_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_326_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_326_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_326_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_327_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_327_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_327_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_327_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_328_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_328_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_328_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_328_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_329_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_329_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_329_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_329_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_330_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_330_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_330_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_330_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_331_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_331_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_331_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_331_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_332_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_332_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_332_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_332_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_333_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_333_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_333_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_333_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_334_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_334_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_334_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_334_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_335_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_335_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_335_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_335_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_336_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_336_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_336_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_336_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_337_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_337_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_337_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_337_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_338_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_338_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_338_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_338_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_339_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_339_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_339_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_339_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_340_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_340_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_340_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_340_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_341_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_341_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_341_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_341_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_342_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_342_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_342_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_342_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_343_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_343_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_343_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_343_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_344_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_344_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_344_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_344_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_345_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_345_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_345_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_345_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_346_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_346_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_346_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_346_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_347_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_347_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_347_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_347_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_348_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_348_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_348_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_348_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_349_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_349_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_349_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_349_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_350_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_350_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_350_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_350_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_351_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_351_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_351_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_351_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_352_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_352_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_352_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_352_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_353_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_353_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_353_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_353_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_354_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_354_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_354_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_354_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_355_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_355_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_355_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_355_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_356_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_356_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_356_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_356_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_357_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_357_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_357_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_357_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_358_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_358_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_358_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_358_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_359_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_359_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_359_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_359_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_360_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_360_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_360_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_360_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_361_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_361_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_361_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_361_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_362_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_362_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_362_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_362_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_363_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_363_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_363_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_363_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_364_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_364_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_364_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_364_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_365_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_365_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_365_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_365_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_366_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_366_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_366_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_366_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_367_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_367_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_367_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_367_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_368_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_368_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_368_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_368_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_369_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_369_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_369_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_369_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_370_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_370_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_370_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_370_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_371_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_371_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_371_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_371_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_372_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_372_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_372_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_372_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_373_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_373_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_373_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_373_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_374_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_374_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_374_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_374_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_375_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_375_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_375_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_375_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_376_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_376_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_376_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_376_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_377_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_377_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_377_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_377_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_378_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_378_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_378_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_378_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_379_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_379_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_379_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_379_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_380_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_380_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_380_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_380_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_381_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_381_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_381_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_381_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_382_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_382_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_382_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_382_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_383_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_383_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_383_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_383_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_384_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_384_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_384_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_384_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_385_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_385_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_385_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_385_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_386_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_386_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_386_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_386_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_387_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_387_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_387_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_387_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_388_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_388_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_388_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_388_pdest);
    pkt_str = $sformatf("%sio_diffCommits_info_389_ldest = 0x%0h ",pkt_str,this.io_diffCommits_info_389_ldest);
    pkt_str = $sformatf("%sio_diffCommits_info_389_pdest = 0x%0h ",pkt_str,this.io_diffCommits_info_389_pdest);
    pkt_str = $sformatf("%sio_lsq_scommit = 0x%0h ",pkt_str,this.io_lsq_scommit);
    pkt_str = $sformatf("%sio_lsq_pendingMMIOld = 0x%0h ",pkt_str,this.io_lsq_pendingMMIOld);
    pkt_str = $sformatf("%sio_lsq_pendingst = 0x%0h ",pkt_str,this.io_lsq_pendingst);
    pkt_str = $sformatf("%sio_lsq_pendingPtr_flag = 0x%0h ",pkt_str,this.io_lsq_pendingPtr_flag);
    pkt_str = $sformatf("%sio_lsq_pendingPtr_value = 0x%0h ",pkt_str,this.io_lsq_pendingPtr_value);
    pkt_str = $sformatf("%sio_robDeqPtr_flag = 0x%0h ",pkt_str,this.io_robDeqPtr_flag);
    pkt_str = $sformatf("%sio_robDeqPtr_value = 0x%0h ",pkt_str,this.io_robDeqPtr_value);
    pkt_str = $sformatf("%sio_csr_fflags_valid = 0x%0h ",pkt_str,this.io_csr_fflags_valid);
    pkt_str = $sformatf("%sio_csr_fflags_bits = 0x%0h ",pkt_str,this.io_csr_fflags_bits);
    pkt_str = $sformatf("%sio_csr_vxsat_valid = 0x%0h ",pkt_str,this.io_csr_vxsat_valid);
    pkt_str = $sformatf("%sio_csr_vxsat_bits = 0x%0h ",pkt_str,this.io_csr_vxsat_bits);
    pkt_str = $sformatf("%sio_csr_vstart_valid = 0x%0h ",pkt_str,this.io_csr_vstart_valid);
    pkt_str = $sformatf("%sio_csr_vstart_bits = 0x%0h ",pkt_str,this.io_csr_vstart_bits);
    pkt_str = $sformatf("%sio_csr_dirty_fs = 0x%0h ",pkt_str,this.io_csr_dirty_fs);
    pkt_str = $sformatf("%sio_csr_dirty_vs = 0x%0h ",pkt_str,this.io_csr_dirty_vs);
    pkt_str = $sformatf("%sio_csr_perfinfo_retiredInstr = 0x%0h ",pkt_str,this.io_csr_perfinfo_retiredInstr);
    pkt_str = $sformatf("%sio_cpu_halt = 0x%0h ",pkt_str,this.io_cpu_halt);
    pkt_str = $sformatf("%sio_wfi_wfiReq = 0x%0h ",pkt_str,this.io_wfi_wfiReq);
    pkt_str = $sformatf("%sio_toDecode_isResumeVType = 0x%0h ",pkt_str,this.io_toDecode_isResumeVType);
    pkt_str = $sformatf("%sio_toDecode_walkToArchVType = 0x%0h ",pkt_str,this.io_toDecode_walkToArchVType);
    pkt_str = $sformatf("%sio_toDecode_walkVType_valid = 0x%0h ",pkt_str,this.io_toDecode_walkVType_valid);
    pkt_str = $sformatf("%sio_toDecode_walkVType_bits_illegal = 0x%0h ",pkt_str,this.io_toDecode_walkVType_bits_illegal);
    pkt_str = $sformatf("%sio_toDecode_walkVType_bits_vma = 0x%0h ",pkt_str,this.io_toDecode_walkVType_bits_vma);
    pkt_str = $sformatf("%sio_toDecode_walkVType_bits_vta = 0x%0h ",pkt_str,this.io_toDecode_walkVType_bits_vta);
    pkt_str = $sformatf("%sio_toDecode_walkVType_bits_vsew = 0x%0h ",pkt_str,this.io_toDecode_walkVType_bits_vsew);
    pkt_str = $sformatf("%sio_toDecode_walkVType_bits_vlmul = 0x%0h ",pkt_str,this.io_toDecode_walkVType_bits_vlmul);
    pkt_str = $sformatf("%sio_toDecode_commitVType_vtype_valid = 0x%0h ",pkt_str,this.io_toDecode_commitVType_vtype_valid);
    pkt_str = $sformatf("%sio_toDecode_commitVType_vtype_bits_illegal = 0x%0h ",pkt_str,this.io_toDecode_commitVType_vtype_bits_illegal);
    pkt_str = $sformatf("%sio_toDecode_commitVType_vtype_bits_vma = 0x%0h ",pkt_str,this.io_toDecode_commitVType_vtype_bits_vma);
    pkt_str = $sformatf("%sio_toDecode_commitVType_vtype_bits_vta = 0x%0h ",pkt_str,this.io_toDecode_commitVType_vtype_bits_vta);
    pkt_str = $sformatf("%sio_toDecode_commitVType_vtype_bits_vsew = 0x%0h ",pkt_str,this.io_toDecode_commitVType_vtype_bits_vsew);
    pkt_str = $sformatf("%sio_toDecode_commitVType_vtype_bits_vlmul = 0x%0h ",pkt_str,this.io_toDecode_commitVType_vtype_bits_vlmul);
    pkt_str = $sformatf("%sio_toDecode_commitVType_hasVsetvl = 0x%0h ",pkt_str,this.io_toDecode_commitVType_hasVsetvl);
    pkt_str = $sformatf("%sio_readGPAMemAddr_valid = 0x%0h ",pkt_str,this.io_readGPAMemAddr_valid);
    pkt_str = $sformatf("%sio_readGPAMemAddr_bits_ftqPtr_value = 0x%0h ",pkt_str,this.io_readGPAMemAddr_bits_ftqPtr_value);
    pkt_str = $sformatf("%sio_readGPAMemAddr_bits_ftqOffset = 0x%0h ",pkt_str,this.io_readGPAMemAddr_bits_ftqOffset);
    pkt_str = $sformatf("%sio_toVecExcpMod_logicPhyRegMap_0_valid = 0x%0h ",pkt_str,this.io_toVecExcpMod_logicPhyRegMap_0_valid);
    pkt_str = $sformatf("%sio_toVecExcpMod_logicPhyRegMap_0_bits_lreg = 0x%0h ",pkt_str,this.io_toVecExcpMod_logicPhyRegMap_0_bits_lreg);
    pkt_str = $sformatf("%sio_toVecExcpMod_logicPhyRegMap_0_bits_preg = 0x%0h ",pkt_str,this.io_toVecExcpMod_logicPhyRegMap_0_bits_preg);
    pkt_str = $sformatf("%sio_toVecExcpMod_logicPhyRegMap_1_valid = 0x%0h ",pkt_str,this.io_toVecExcpMod_logicPhyRegMap_1_valid);
    pkt_str = $sformatf("%sio_toVecExcpMod_logicPhyRegMap_1_bits_lreg = 0x%0h ",pkt_str,this.io_toVecExcpMod_logicPhyRegMap_1_bits_lreg);
    pkt_str = $sformatf("%sio_toVecExcpMod_logicPhyRegMap_1_bits_preg = 0x%0h ",pkt_str,this.io_toVecExcpMod_logicPhyRegMap_1_bits_preg);
    pkt_str = $sformatf("%sio_toVecExcpMod_logicPhyRegMap_2_valid = 0x%0h ",pkt_str,this.io_toVecExcpMod_logicPhyRegMap_2_valid);
    pkt_str = $sformatf("%sio_toVecExcpMod_logicPhyRegMap_2_bits_lreg = 0x%0h ",pkt_str,this.io_toVecExcpMod_logicPhyRegMap_2_bits_lreg);
    pkt_str = $sformatf("%sio_toVecExcpMod_logicPhyRegMap_2_bits_preg = 0x%0h ",pkt_str,this.io_toVecExcpMod_logicPhyRegMap_2_bits_preg);
    pkt_str = $sformatf("%sio_toVecExcpMod_logicPhyRegMap_3_valid = 0x%0h ",pkt_str,this.io_toVecExcpMod_logicPhyRegMap_3_valid);
    pkt_str = $sformatf("%sio_toVecExcpMod_logicPhyRegMap_3_bits_lreg = 0x%0h ",pkt_str,this.io_toVecExcpMod_logicPhyRegMap_3_bits_lreg);
    pkt_str = $sformatf("%sio_toVecExcpMod_logicPhyRegMap_3_bits_preg = 0x%0h ",pkt_str,this.io_toVecExcpMod_logicPhyRegMap_3_bits_preg);
    pkt_str = $sformatf("%sio_toVecExcpMod_logicPhyRegMap_4_valid = 0x%0h ",pkt_str,this.io_toVecExcpMod_logicPhyRegMap_4_valid);
    pkt_str = $sformatf("%sio_toVecExcpMod_logicPhyRegMap_4_bits_lreg = 0x%0h ",pkt_str,this.io_toVecExcpMod_logicPhyRegMap_4_bits_lreg);
    pkt_str = $sformatf("%sio_toVecExcpMod_logicPhyRegMap_4_bits_preg = 0x%0h ",pkt_str,this.io_toVecExcpMod_logicPhyRegMap_4_bits_preg);
    pkt_str = $sformatf("%sio_toVecExcpMod_logicPhyRegMap_5_valid = 0x%0h ",pkt_str,this.io_toVecExcpMod_logicPhyRegMap_5_valid);
    pkt_str = $sformatf("%sio_toVecExcpMod_logicPhyRegMap_5_bits_lreg = 0x%0h ",pkt_str,this.io_toVecExcpMod_logicPhyRegMap_5_bits_lreg);
    pkt_str = $sformatf("%sio_toVecExcpMod_logicPhyRegMap_5_bits_preg = 0x%0h ",pkt_str,this.io_toVecExcpMod_logicPhyRegMap_5_bits_preg);
    pkt_str = $sformatf("%sio_toVecExcpMod_excpInfo_valid = 0x%0h ",pkt_str,this.io_toVecExcpMod_excpInfo_valid);
    pkt_str = $sformatf("%sio_toVecExcpMod_excpInfo_bits_vstart = 0x%0h ",pkt_str,this.io_toVecExcpMod_excpInfo_bits_vstart);
    pkt_str = $sformatf("%sio_toVecExcpMod_excpInfo_bits_vsew = 0x%0h ",pkt_str,this.io_toVecExcpMod_excpInfo_bits_vsew);
    pkt_str = $sformatf("%sio_toVecExcpMod_excpInfo_bits_veew = 0x%0h ",pkt_str,this.io_toVecExcpMod_excpInfo_bits_veew);
    pkt_str = $sformatf("%sio_toVecExcpMod_excpInfo_bits_vlmul = 0x%0h ",pkt_str,this.io_toVecExcpMod_excpInfo_bits_vlmul);
    pkt_str = $sformatf("%sio_toVecExcpMod_excpInfo_bits_nf = 0x%0h ",pkt_str,this.io_toVecExcpMod_excpInfo_bits_nf);
    pkt_str = $sformatf("%sio_toVecExcpMod_excpInfo_bits_isStride = 0x%0h ",pkt_str,this.io_toVecExcpMod_excpInfo_bits_isStride);
    pkt_str = $sformatf("%sio_toVecExcpMod_excpInfo_bits_isIndexed = 0x%0h ",pkt_str,this.io_toVecExcpMod_excpInfo_bits_isIndexed);
    pkt_str = $sformatf("%sio_toVecExcpMod_excpInfo_bits_isWhole = 0x%0h ",pkt_str,this.io_toVecExcpMod_excpInfo_bits_isWhole);
    pkt_str = $sformatf("%sio_toVecExcpMod_excpInfo_bits_isVlm = 0x%0h ",pkt_str,this.io_toVecExcpMod_excpInfo_bits_isVlm);
    pkt_str = $sformatf("%sio_storeDebugInfo_1_pc = 0x%0h ",pkt_str,this.io_storeDebugInfo_1_pc);
    pkt_str = $sformatf("%sio_perf_0_value = 0x%0h ",pkt_str,this.io_perf_0_value);
    pkt_str = $sformatf("%sio_perf_1_value = 0x%0h ",pkt_str,this.io_perf_1_value);
    pkt_str = $sformatf("%sio_perf_2_value = 0x%0h ",pkt_str,this.io_perf_2_value);
    pkt_str = $sformatf("%sio_perf_3_value = 0x%0h ",pkt_str,this.io_perf_3_value);
    pkt_str = $sformatf("%sio_perf_4_value = 0x%0h ",pkt_str,this.io_perf_4_value);
    pkt_str = $sformatf("%sio_perf_5_value = 0x%0h ",pkt_str,this.io_perf_5_value);
    pkt_str = $sformatf("%sio_perf_6_value = 0x%0h ",pkt_str,this.io_perf_6_value);
    pkt_str = $sformatf("%sio_perf_7_value = 0x%0h ",pkt_str,this.io_perf_7_value);
    pkt_str = $sformatf("%sio_perf_8_value = 0x%0h ",pkt_str,this.io_perf_8_value);
    pkt_str = $sformatf("%sio_perf_9_value = 0x%0h ",pkt_str,this.io_perf_9_value);
    pkt_str = $sformatf("%sio_perf_10_value = 0x%0h ",pkt_str,this.io_perf_10_value);
    pkt_str = $sformatf("%sio_perf_11_value = 0x%0h ",pkt_str,this.io_perf_11_value);
    pkt_str = $sformatf("%sio_perf_12_value = 0x%0h ",pkt_str,this.io_perf_12_value);
    pkt_str = $sformatf("%sio_perf_13_value = 0x%0h ",pkt_str,this.io_perf_13_value);
    pkt_str = $sformatf("%sio_perf_14_value = 0x%0h ",pkt_str,this.io_perf_14_value);
    pkt_str = $sformatf("%sio_perf_15_value = 0x%0h ",pkt_str,this.io_perf_15_value);
    pkt_str = $sformatf("%sio_perf_16_value = 0x%0h ",pkt_str,this.io_perf_16_value);
    pkt_str = $sformatf("%sio_perf_17_value = 0x%0h ",pkt_str,this.io_perf_17_value);
    pkt_str = $sformatf("%sio_error_0 = 0x%0h ",pkt_str,this.io_error_0);

    return pkt_str;
endfunction:psdisplay

function bit Rob_output_agent_xaction::compare(uvm_object rhs, uvm_comparer comparer=null);
    bit super_result;
    Rob_output_agent_xaction  rhs_;
    if(!$cast(rhs_, rhs)) begin
        `uvm_fatal(get_type_name(),$sformatf("rhs is not a Rob_output_agent_xaction or its extend"))
    end
    super_result = super.compare(rhs_,comparer);
    if(super_result==0) begin
        super_result = 1;
        //foreach(this.pload_q[i]) begin
        //    if(this.pload_q[i]!=rhs_.pload_q[i]) begin
        //        super_result = 0;
        //        `uvm_info(get_type_name(),$sformatf("compare fail for this.pload[%0d]=0x%2h while the rhs_.pload[%0d]=0x%2h",i,this.pload_q[i],i,rhs_.pload_q[i]),UVM_NONE)
        //    end
        //end

        if(this.io_enq_canAccept!=rhs_.io_enq_canAccept) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_enq_canAccept=0x%0h while the rhs_.io_enq_canAccept=0x%0h",this.io_enq_canAccept,rhs_.io_enq_canAccept),UVM_NONE)
        end

        if(this.io_enq_canAcceptForDispatch!=rhs_.io_enq_canAcceptForDispatch) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_enq_canAcceptForDispatch=0x%0h while the rhs_.io_enq_canAcceptForDispatch=0x%0h",this.io_enq_canAcceptForDispatch,rhs_.io_enq_canAcceptForDispatch),UVM_NONE)
        end

        if(this.io_enq_isEmpty!=rhs_.io_enq_isEmpty) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_enq_isEmpty=0x%0h while the rhs_.io_enq_isEmpty=0x%0h",this.io_enq_isEmpty,rhs_.io_enq_isEmpty),UVM_NONE)
        end

        if(this.io_flushOut_valid!=rhs_.io_flushOut_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_flushOut_valid=0x%0h while the rhs_.io_flushOut_valid=0x%0h",this.io_flushOut_valid,rhs_.io_flushOut_valid),UVM_NONE)
        end

        if(this.io_flushOut_bits_isRVC!=rhs_.io_flushOut_bits_isRVC) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_flushOut_bits_isRVC=0x%0h while the rhs_.io_flushOut_bits_isRVC=0x%0h",this.io_flushOut_bits_isRVC,rhs_.io_flushOut_bits_isRVC),UVM_NONE)
        end

        if(this.io_flushOut_bits_robIdx_flag!=rhs_.io_flushOut_bits_robIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_flushOut_bits_robIdx_flag=0x%0h while the rhs_.io_flushOut_bits_robIdx_flag=0x%0h",this.io_flushOut_bits_robIdx_flag,rhs_.io_flushOut_bits_robIdx_flag),UVM_NONE)
        end

        if(this.io_flushOut_bits_robIdx_value!=rhs_.io_flushOut_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_flushOut_bits_robIdx_value=0x%0h while the rhs_.io_flushOut_bits_robIdx_value=0x%0h",this.io_flushOut_bits_robIdx_value,rhs_.io_flushOut_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_flushOut_bits_ftqIdx_flag!=rhs_.io_flushOut_bits_ftqIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_flushOut_bits_ftqIdx_flag=0x%0h while the rhs_.io_flushOut_bits_ftqIdx_flag=0x%0h",this.io_flushOut_bits_ftqIdx_flag,rhs_.io_flushOut_bits_ftqIdx_flag),UVM_NONE)
        end

        if(this.io_flushOut_bits_ftqIdx_value!=rhs_.io_flushOut_bits_ftqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_flushOut_bits_ftqIdx_value=0x%0h while the rhs_.io_flushOut_bits_ftqIdx_value=0x%0h",this.io_flushOut_bits_ftqIdx_value,rhs_.io_flushOut_bits_ftqIdx_value),UVM_NONE)
        end

        if(this.io_flushOut_bits_ftqOffset!=rhs_.io_flushOut_bits_ftqOffset) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_flushOut_bits_ftqOffset=0x%0h while the rhs_.io_flushOut_bits_ftqOffset=0x%0h",this.io_flushOut_bits_ftqOffset,rhs_.io_flushOut_bits_ftqOffset),UVM_NONE)
        end

        if(this.io_flushOut_bits_level!=rhs_.io_flushOut_bits_level) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_flushOut_bits_level=0x%0h while the rhs_.io_flushOut_bits_level=0x%0h",this.io_flushOut_bits_level,rhs_.io_flushOut_bits_level),UVM_NONE)
        end

        if(this.io_exception_valid!=rhs_.io_exception_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_valid=0x%0h while the rhs_.io_exception_valid=0x%0h",this.io_exception_valid,rhs_.io_exception_valid),UVM_NONE)
        end

        if(this.io_exception_bits_instr!=rhs_.io_exception_bits_instr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_instr=0x%0h while the rhs_.io_exception_bits_instr=0x%0h",this.io_exception_bits_instr,rhs_.io_exception_bits_instr),UVM_NONE)
        end

        if(this.io_exception_bits_commitType!=rhs_.io_exception_bits_commitType) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_commitType=0x%0h while the rhs_.io_exception_bits_commitType=0x%0h",this.io_exception_bits_commitType,rhs_.io_exception_bits_commitType),UVM_NONE)
        end

        if(this.io_exception_bits_exceptionVec_0!=rhs_.io_exception_bits_exceptionVec_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_exceptionVec_0=0x%0h while the rhs_.io_exception_bits_exceptionVec_0=0x%0h",this.io_exception_bits_exceptionVec_0,rhs_.io_exception_bits_exceptionVec_0),UVM_NONE)
        end

        if(this.io_exception_bits_exceptionVec_1!=rhs_.io_exception_bits_exceptionVec_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_exceptionVec_1=0x%0h while the rhs_.io_exception_bits_exceptionVec_1=0x%0h",this.io_exception_bits_exceptionVec_1,rhs_.io_exception_bits_exceptionVec_1),UVM_NONE)
        end

        if(this.io_exception_bits_exceptionVec_2!=rhs_.io_exception_bits_exceptionVec_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_exceptionVec_2=0x%0h while the rhs_.io_exception_bits_exceptionVec_2=0x%0h",this.io_exception_bits_exceptionVec_2,rhs_.io_exception_bits_exceptionVec_2),UVM_NONE)
        end

        if(this.io_exception_bits_exceptionVec_3!=rhs_.io_exception_bits_exceptionVec_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_exceptionVec_3=0x%0h while the rhs_.io_exception_bits_exceptionVec_3=0x%0h",this.io_exception_bits_exceptionVec_3,rhs_.io_exception_bits_exceptionVec_3),UVM_NONE)
        end

        if(this.io_exception_bits_exceptionVec_4!=rhs_.io_exception_bits_exceptionVec_4) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_exceptionVec_4=0x%0h while the rhs_.io_exception_bits_exceptionVec_4=0x%0h",this.io_exception_bits_exceptionVec_4,rhs_.io_exception_bits_exceptionVec_4),UVM_NONE)
        end

        if(this.io_exception_bits_exceptionVec_5!=rhs_.io_exception_bits_exceptionVec_5) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_exceptionVec_5=0x%0h while the rhs_.io_exception_bits_exceptionVec_5=0x%0h",this.io_exception_bits_exceptionVec_5,rhs_.io_exception_bits_exceptionVec_5),UVM_NONE)
        end

        if(this.io_exception_bits_exceptionVec_6!=rhs_.io_exception_bits_exceptionVec_6) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_exceptionVec_6=0x%0h while the rhs_.io_exception_bits_exceptionVec_6=0x%0h",this.io_exception_bits_exceptionVec_6,rhs_.io_exception_bits_exceptionVec_6),UVM_NONE)
        end

        if(this.io_exception_bits_exceptionVec_7!=rhs_.io_exception_bits_exceptionVec_7) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_exceptionVec_7=0x%0h while the rhs_.io_exception_bits_exceptionVec_7=0x%0h",this.io_exception_bits_exceptionVec_7,rhs_.io_exception_bits_exceptionVec_7),UVM_NONE)
        end

        if(this.io_exception_bits_exceptionVec_8!=rhs_.io_exception_bits_exceptionVec_8) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_exceptionVec_8=0x%0h while the rhs_.io_exception_bits_exceptionVec_8=0x%0h",this.io_exception_bits_exceptionVec_8,rhs_.io_exception_bits_exceptionVec_8),UVM_NONE)
        end

        if(this.io_exception_bits_exceptionVec_9!=rhs_.io_exception_bits_exceptionVec_9) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_exceptionVec_9=0x%0h while the rhs_.io_exception_bits_exceptionVec_9=0x%0h",this.io_exception_bits_exceptionVec_9,rhs_.io_exception_bits_exceptionVec_9),UVM_NONE)
        end

        if(this.io_exception_bits_exceptionVec_10!=rhs_.io_exception_bits_exceptionVec_10) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_exceptionVec_10=0x%0h while the rhs_.io_exception_bits_exceptionVec_10=0x%0h",this.io_exception_bits_exceptionVec_10,rhs_.io_exception_bits_exceptionVec_10),UVM_NONE)
        end

        if(this.io_exception_bits_exceptionVec_11!=rhs_.io_exception_bits_exceptionVec_11) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_exceptionVec_11=0x%0h while the rhs_.io_exception_bits_exceptionVec_11=0x%0h",this.io_exception_bits_exceptionVec_11,rhs_.io_exception_bits_exceptionVec_11),UVM_NONE)
        end

        if(this.io_exception_bits_exceptionVec_12!=rhs_.io_exception_bits_exceptionVec_12) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_exceptionVec_12=0x%0h while the rhs_.io_exception_bits_exceptionVec_12=0x%0h",this.io_exception_bits_exceptionVec_12,rhs_.io_exception_bits_exceptionVec_12),UVM_NONE)
        end

        if(this.io_exception_bits_exceptionVec_13!=rhs_.io_exception_bits_exceptionVec_13) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_exceptionVec_13=0x%0h while the rhs_.io_exception_bits_exceptionVec_13=0x%0h",this.io_exception_bits_exceptionVec_13,rhs_.io_exception_bits_exceptionVec_13),UVM_NONE)
        end

        if(this.io_exception_bits_exceptionVec_14!=rhs_.io_exception_bits_exceptionVec_14) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_exceptionVec_14=0x%0h while the rhs_.io_exception_bits_exceptionVec_14=0x%0h",this.io_exception_bits_exceptionVec_14,rhs_.io_exception_bits_exceptionVec_14),UVM_NONE)
        end

        if(this.io_exception_bits_exceptionVec_15!=rhs_.io_exception_bits_exceptionVec_15) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_exceptionVec_15=0x%0h while the rhs_.io_exception_bits_exceptionVec_15=0x%0h",this.io_exception_bits_exceptionVec_15,rhs_.io_exception_bits_exceptionVec_15),UVM_NONE)
        end

        if(this.io_exception_bits_exceptionVec_16!=rhs_.io_exception_bits_exceptionVec_16) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_exceptionVec_16=0x%0h while the rhs_.io_exception_bits_exceptionVec_16=0x%0h",this.io_exception_bits_exceptionVec_16,rhs_.io_exception_bits_exceptionVec_16),UVM_NONE)
        end

        if(this.io_exception_bits_exceptionVec_17!=rhs_.io_exception_bits_exceptionVec_17) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_exceptionVec_17=0x%0h while the rhs_.io_exception_bits_exceptionVec_17=0x%0h",this.io_exception_bits_exceptionVec_17,rhs_.io_exception_bits_exceptionVec_17),UVM_NONE)
        end

        if(this.io_exception_bits_exceptionVec_18!=rhs_.io_exception_bits_exceptionVec_18) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_exceptionVec_18=0x%0h while the rhs_.io_exception_bits_exceptionVec_18=0x%0h",this.io_exception_bits_exceptionVec_18,rhs_.io_exception_bits_exceptionVec_18),UVM_NONE)
        end

        if(this.io_exception_bits_exceptionVec_19!=rhs_.io_exception_bits_exceptionVec_19) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_exceptionVec_19=0x%0h while the rhs_.io_exception_bits_exceptionVec_19=0x%0h",this.io_exception_bits_exceptionVec_19,rhs_.io_exception_bits_exceptionVec_19),UVM_NONE)
        end

        if(this.io_exception_bits_exceptionVec_20!=rhs_.io_exception_bits_exceptionVec_20) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_exceptionVec_20=0x%0h while the rhs_.io_exception_bits_exceptionVec_20=0x%0h",this.io_exception_bits_exceptionVec_20,rhs_.io_exception_bits_exceptionVec_20),UVM_NONE)
        end

        if(this.io_exception_bits_exceptionVec_21!=rhs_.io_exception_bits_exceptionVec_21) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_exceptionVec_21=0x%0h while the rhs_.io_exception_bits_exceptionVec_21=0x%0h",this.io_exception_bits_exceptionVec_21,rhs_.io_exception_bits_exceptionVec_21),UVM_NONE)
        end

        if(this.io_exception_bits_exceptionVec_22!=rhs_.io_exception_bits_exceptionVec_22) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_exceptionVec_22=0x%0h while the rhs_.io_exception_bits_exceptionVec_22=0x%0h",this.io_exception_bits_exceptionVec_22,rhs_.io_exception_bits_exceptionVec_22),UVM_NONE)
        end

        if(this.io_exception_bits_exceptionVec_23!=rhs_.io_exception_bits_exceptionVec_23) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_exceptionVec_23=0x%0h while the rhs_.io_exception_bits_exceptionVec_23=0x%0h",this.io_exception_bits_exceptionVec_23,rhs_.io_exception_bits_exceptionVec_23),UVM_NONE)
        end

        if(this.io_exception_bits_isPcBkpt!=rhs_.io_exception_bits_isPcBkpt) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_isPcBkpt=0x%0h while the rhs_.io_exception_bits_isPcBkpt=0x%0h",this.io_exception_bits_isPcBkpt,rhs_.io_exception_bits_isPcBkpt),UVM_NONE)
        end

        if(this.io_exception_bits_isFetchMalAddr!=rhs_.io_exception_bits_isFetchMalAddr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_isFetchMalAddr=0x%0h while the rhs_.io_exception_bits_isFetchMalAddr=0x%0h",this.io_exception_bits_isFetchMalAddr,rhs_.io_exception_bits_isFetchMalAddr),UVM_NONE)
        end

        if(this.io_exception_bits_gpaddr!=rhs_.io_exception_bits_gpaddr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_gpaddr=0x%0h while the rhs_.io_exception_bits_gpaddr=0x%0h",this.io_exception_bits_gpaddr,rhs_.io_exception_bits_gpaddr),UVM_NONE)
        end

        if(this.io_exception_bits_singleStep!=rhs_.io_exception_bits_singleStep) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_singleStep=0x%0h while the rhs_.io_exception_bits_singleStep=0x%0h",this.io_exception_bits_singleStep,rhs_.io_exception_bits_singleStep),UVM_NONE)
        end

        if(this.io_exception_bits_crossPageIPFFix!=rhs_.io_exception_bits_crossPageIPFFix) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_crossPageIPFFix=0x%0h while the rhs_.io_exception_bits_crossPageIPFFix=0x%0h",this.io_exception_bits_crossPageIPFFix,rhs_.io_exception_bits_crossPageIPFFix),UVM_NONE)
        end

        if(this.io_exception_bits_isInterrupt!=rhs_.io_exception_bits_isInterrupt) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_isInterrupt=0x%0h while the rhs_.io_exception_bits_isInterrupt=0x%0h",this.io_exception_bits_isInterrupt,rhs_.io_exception_bits_isInterrupt),UVM_NONE)
        end

        if(this.io_exception_bits_isHls!=rhs_.io_exception_bits_isHls) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_isHls=0x%0h while the rhs_.io_exception_bits_isHls=0x%0h",this.io_exception_bits_isHls,rhs_.io_exception_bits_isHls),UVM_NONE)
        end

        if(this.io_exception_bits_trigger!=rhs_.io_exception_bits_trigger) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_trigger=0x%0h while the rhs_.io_exception_bits_trigger=0x%0h",this.io_exception_bits_trigger,rhs_.io_exception_bits_trigger),UVM_NONE)
        end

        if(this.io_exception_bits_isForVSnonLeafPTE!=rhs_.io_exception_bits_isForVSnonLeafPTE) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exception_bits_isForVSnonLeafPTE=0x%0h while the rhs_.io_exception_bits_isForVSnonLeafPTE=0x%0h",this.io_exception_bits_isForVSnonLeafPTE,rhs_.io_exception_bits_isForVSnonLeafPTE),UVM_NONE)
        end

        if(this.io_commits_isCommit!=rhs_.io_commits_isCommit) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_isCommit=0x%0h while the rhs_.io_commits_isCommit=0x%0h",this.io_commits_isCommit,rhs_.io_commits_isCommit),UVM_NONE)
        end

        if(this.io_commits_commitValid_0!=rhs_.io_commits_commitValid_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_commitValid_0=0x%0h while the rhs_.io_commits_commitValid_0=0x%0h",this.io_commits_commitValid_0,rhs_.io_commits_commitValid_0),UVM_NONE)
        end

        if(this.io_commits_commitValid_1!=rhs_.io_commits_commitValid_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_commitValid_1=0x%0h while the rhs_.io_commits_commitValid_1=0x%0h",this.io_commits_commitValid_1,rhs_.io_commits_commitValid_1),UVM_NONE)
        end

        if(this.io_commits_commitValid_2!=rhs_.io_commits_commitValid_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_commitValid_2=0x%0h while the rhs_.io_commits_commitValid_2=0x%0h",this.io_commits_commitValid_2,rhs_.io_commits_commitValid_2),UVM_NONE)
        end

        if(this.io_commits_commitValid_3!=rhs_.io_commits_commitValid_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_commitValid_3=0x%0h while the rhs_.io_commits_commitValid_3=0x%0h",this.io_commits_commitValid_3,rhs_.io_commits_commitValid_3),UVM_NONE)
        end

        if(this.io_commits_commitValid_4!=rhs_.io_commits_commitValid_4) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_commitValid_4=0x%0h while the rhs_.io_commits_commitValid_4=0x%0h",this.io_commits_commitValid_4,rhs_.io_commits_commitValid_4),UVM_NONE)
        end

        if(this.io_commits_commitValid_5!=rhs_.io_commits_commitValid_5) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_commitValid_5=0x%0h while the rhs_.io_commits_commitValid_5=0x%0h",this.io_commits_commitValid_5,rhs_.io_commits_commitValid_5),UVM_NONE)
        end

        if(this.io_commits_commitValid_6!=rhs_.io_commits_commitValid_6) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_commitValid_6=0x%0h while the rhs_.io_commits_commitValid_6=0x%0h",this.io_commits_commitValid_6,rhs_.io_commits_commitValid_6),UVM_NONE)
        end

        if(this.io_commits_commitValid_7!=rhs_.io_commits_commitValid_7) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_commitValid_7=0x%0h while the rhs_.io_commits_commitValid_7=0x%0h",this.io_commits_commitValid_7,rhs_.io_commits_commitValid_7),UVM_NONE)
        end

        if(this.io_commits_isWalk!=rhs_.io_commits_isWalk) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_isWalk=0x%0h while the rhs_.io_commits_isWalk=0x%0h",this.io_commits_isWalk,rhs_.io_commits_isWalk),UVM_NONE)
        end

        if(this.io_commits_walkValid_0!=rhs_.io_commits_walkValid_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_walkValid_0=0x%0h while the rhs_.io_commits_walkValid_0=0x%0h",this.io_commits_walkValid_0,rhs_.io_commits_walkValid_0),UVM_NONE)
        end

        if(this.io_commits_walkValid_1!=rhs_.io_commits_walkValid_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_walkValid_1=0x%0h while the rhs_.io_commits_walkValid_1=0x%0h",this.io_commits_walkValid_1,rhs_.io_commits_walkValid_1),UVM_NONE)
        end

        if(this.io_commits_walkValid_2!=rhs_.io_commits_walkValid_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_walkValid_2=0x%0h while the rhs_.io_commits_walkValid_2=0x%0h",this.io_commits_walkValid_2,rhs_.io_commits_walkValid_2),UVM_NONE)
        end

        if(this.io_commits_walkValid_3!=rhs_.io_commits_walkValid_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_walkValid_3=0x%0h while the rhs_.io_commits_walkValid_3=0x%0h",this.io_commits_walkValid_3,rhs_.io_commits_walkValid_3),UVM_NONE)
        end

        if(this.io_commits_walkValid_4!=rhs_.io_commits_walkValid_4) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_walkValid_4=0x%0h while the rhs_.io_commits_walkValid_4=0x%0h",this.io_commits_walkValid_4,rhs_.io_commits_walkValid_4),UVM_NONE)
        end

        if(this.io_commits_walkValid_5!=rhs_.io_commits_walkValid_5) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_walkValid_5=0x%0h while the rhs_.io_commits_walkValid_5=0x%0h",this.io_commits_walkValid_5,rhs_.io_commits_walkValid_5),UVM_NONE)
        end

        if(this.io_commits_walkValid_6!=rhs_.io_commits_walkValid_6) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_walkValid_6=0x%0h while the rhs_.io_commits_walkValid_6=0x%0h",this.io_commits_walkValid_6,rhs_.io_commits_walkValid_6),UVM_NONE)
        end

        if(this.io_commits_walkValid_7!=rhs_.io_commits_walkValid_7) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_walkValid_7=0x%0h while the rhs_.io_commits_walkValid_7=0x%0h",this.io_commits_walkValid_7,rhs_.io_commits_walkValid_7),UVM_NONE)
        end

        if(this.io_commits_info_0_walk_v!=rhs_.io_commits_info_0_walk_v) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_walk_v=0x%0h while the rhs_.io_commits_info_0_walk_v=0x%0h",this.io_commits_info_0_walk_v,rhs_.io_commits_info_0_walk_v),UVM_NONE)
        end

        if(this.io_commits_info_0_commit_v!=rhs_.io_commits_info_0_commit_v) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_commit_v=0x%0h while the rhs_.io_commits_info_0_commit_v=0x%0h",this.io_commits_info_0_commit_v,rhs_.io_commits_info_0_commit_v),UVM_NONE)
        end

        if(this.io_commits_info_0_commit_w!=rhs_.io_commits_info_0_commit_w) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_commit_w=0x%0h while the rhs_.io_commits_info_0_commit_w=0x%0h",this.io_commits_info_0_commit_w,rhs_.io_commits_info_0_commit_w),UVM_NONE)
        end

        if(this.io_commits_info_0_realDestSize!=rhs_.io_commits_info_0_realDestSize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_realDestSize=0x%0h while the rhs_.io_commits_info_0_realDestSize=0x%0h",this.io_commits_info_0_realDestSize,rhs_.io_commits_info_0_realDestSize),UVM_NONE)
        end

        if(this.io_commits_info_0_interrupt_safe!=rhs_.io_commits_info_0_interrupt_safe) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_interrupt_safe=0x%0h while the rhs_.io_commits_info_0_interrupt_safe=0x%0h",this.io_commits_info_0_interrupt_safe,rhs_.io_commits_info_0_interrupt_safe),UVM_NONE)
        end

        if(this.io_commits_info_0_wflags!=rhs_.io_commits_info_0_wflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_wflags=0x%0h while the rhs_.io_commits_info_0_wflags=0x%0h",this.io_commits_info_0_wflags,rhs_.io_commits_info_0_wflags),UVM_NONE)
        end

        if(this.io_commits_info_0_fflags!=rhs_.io_commits_info_0_fflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_fflags=0x%0h while the rhs_.io_commits_info_0_fflags=0x%0h",this.io_commits_info_0_fflags,rhs_.io_commits_info_0_fflags),UVM_NONE)
        end

        if(this.io_commits_info_0_vxsat!=rhs_.io_commits_info_0_vxsat) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_vxsat=0x%0h while the rhs_.io_commits_info_0_vxsat=0x%0h",this.io_commits_info_0_vxsat,rhs_.io_commits_info_0_vxsat),UVM_NONE)
        end

        if(this.io_commits_info_0_isRVC!=rhs_.io_commits_info_0_isRVC) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_isRVC=0x%0h while the rhs_.io_commits_info_0_isRVC=0x%0h",this.io_commits_info_0_isRVC,rhs_.io_commits_info_0_isRVC),UVM_NONE)
        end

        if(this.io_commits_info_0_isVset!=rhs_.io_commits_info_0_isVset) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_isVset=0x%0h while the rhs_.io_commits_info_0_isVset=0x%0h",this.io_commits_info_0_isVset,rhs_.io_commits_info_0_isVset),UVM_NONE)
        end

        if(this.io_commits_info_0_isHls!=rhs_.io_commits_info_0_isHls) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_isHls=0x%0h while the rhs_.io_commits_info_0_isHls=0x%0h",this.io_commits_info_0_isHls,rhs_.io_commits_info_0_isHls),UVM_NONE)
        end

        if(this.io_commits_info_0_isVls!=rhs_.io_commits_info_0_isVls) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_isVls=0x%0h while the rhs_.io_commits_info_0_isVls=0x%0h",this.io_commits_info_0_isVls,rhs_.io_commits_info_0_isVls),UVM_NONE)
        end

        if(this.io_commits_info_0_vls!=rhs_.io_commits_info_0_vls) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_vls=0x%0h while the rhs_.io_commits_info_0_vls=0x%0h",this.io_commits_info_0_vls,rhs_.io_commits_info_0_vls),UVM_NONE)
        end

        if(this.io_commits_info_0_mmio!=rhs_.io_commits_info_0_mmio) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_mmio=0x%0h while the rhs_.io_commits_info_0_mmio=0x%0h",this.io_commits_info_0_mmio,rhs_.io_commits_info_0_mmio),UVM_NONE)
        end

        if(this.io_commits_info_0_commitType!=rhs_.io_commits_info_0_commitType) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_commitType=0x%0h while the rhs_.io_commits_info_0_commitType=0x%0h",this.io_commits_info_0_commitType,rhs_.io_commits_info_0_commitType),UVM_NONE)
        end

        if(this.io_commits_info_0_ftqIdx_flag!=rhs_.io_commits_info_0_ftqIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_ftqIdx_flag=0x%0h while the rhs_.io_commits_info_0_ftqIdx_flag=0x%0h",this.io_commits_info_0_ftqIdx_flag,rhs_.io_commits_info_0_ftqIdx_flag),UVM_NONE)
        end

        if(this.io_commits_info_0_ftqIdx_value!=rhs_.io_commits_info_0_ftqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_ftqIdx_value=0x%0h while the rhs_.io_commits_info_0_ftqIdx_value=0x%0h",this.io_commits_info_0_ftqIdx_value,rhs_.io_commits_info_0_ftqIdx_value),UVM_NONE)
        end

        if(this.io_commits_info_0_ftqOffset!=rhs_.io_commits_info_0_ftqOffset) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_ftqOffset=0x%0h while the rhs_.io_commits_info_0_ftqOffset=0x%0h",this.io_commits_info_0_ftqOffset,rhs_.io_commits_info_0_ftqOffset),UVM_NONE)
        end

        if(this.io_commits_info_0_instrSize!=rhs_.io_commits_info_0_instrSize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_instrSize=0x%0h while the rhs_.io_commits_info_0_instrSize=0x%0h",this.io_commits_info_0_instrSize,rhs_.io_commits_info_0_instrSize),UVM_NONE)
        end

        if(this.io_commits_info_0_fpWen!=rhs_.io_commits_info_0_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_fpWen=0x%0h while the rhs_.io_commits_info_0_fpWen=0x%0h",this.io_commits_info_0_fpWen,rhs_.io_commits_info_0_fpWen),UVM_NONE)
        end

        if(this.io_commits_info_0_rfWen!=rhs_.io_commits_info_0_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_rfWen=0x%0h while the rhs_.io_commits_info_0_rfWen=0x%0h",this.io_commits_info_0_rfWen,rhs_.io_commits_info_0_rfWen),UVM_NONE)
        end

        if(this.io_commits_info_0_needFlush!=rhs_.io_commits_info_0_needFlush) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_needFlush=0x%0h while the rhs_.io_commits_info_0_needFlush=0x%0h",this.io_commits_info_0_needFlush,rhs_.io_commits_info_0_needFlush),UVM_NONE)
        end

        if(this.io_commits_info_0_traceBlockInPipe_itype!=rhs_.io_commits_info_0_traceBlockInPipe_itype) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_traceBlockInPipe_itype=0x%0h while the rhs_.io_commits_info_0_traceBlockInPipe_itype=0x%0h",this.io_commits_info_0_traceBlockInPipe_itype,rhs_.io_commits_info_0_traceBlockInPipe_itype),UVM_NONE)
        end

        if(this.io_commits_info_0_traceBlockInPipe_iretire!=rhs_.io_commits_info_0_traceBlockInPipe_iretire) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_traceBlockInPipe_iretire=0x%0h while the rhs_.io_commits_info_0_traceBlockInPipe_iretire=0x%0h",this.io_commits_info_0_traceBlockInPipe_iretire,rhs_.io_commits_info_0_traceBlockInPipe_iretire),UVM_NONE)
        end

        if(this.io_commits_info_0_traceBlockInPipe_ilastsize!=rhs_.io_commits_info_0_traceBlockInPipe_ilastsize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_traceBlockInPipe_ilastsize=0x%0h while the rhs_.io_commits_info_0_traceBlockInPipe_ilastsize=0x%0h",this.io_commits_info_0_traceBlockInPipe_ilastsize,rhs_.io_commits_info_0_traceBlockInPipe_ilastsize),UVM_NONE)
        end

        if(this.io_commits_info_0_debug_pc!=rhs_.io_commits_info_0_debug_pc) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_debug_pc=0x%0h while the rhs_.io_commits_info_0_debug_pc=0x%0h",this.io_commits_info_0_debug_pc,rhs_.io_commits_info_0_debug_pc),UVM_NONE)
        end

        if(this.io_commits_info_0_debug_instr!=rhs_.io_commits_info_0_debug_instr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_debug_instr=0x%0h while the rhs_.io_commits_info_0_debug_instr=0x%0h",this.io_commits_info_0_debug_instr,rhs_.io_commits_info_0_debug_instr),UVM_NONE)
        end

        if(this.io_commits_info_0_debug_ldest!=rhs_.io_commits_info_0_debug_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_debug_ldest=0x%0h while the rhs_.io_commits_info_0_debug_ldest=0x%0h",this.io_commits_info_0_debug_ldest,rhs_.io_commits_info_0_debug_ldest),UVM_NONE)
        end

        if(this.io_commits_info_0_debug_pdest!=rhs_.io_commits_info_0_debug_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_debug_pdest=0x%0h while the rhs_.io_commits_info_0_debug_pdest=0x%0h",this.io_commits_info_0_debug_pdest,rhs_.io_commits_info_0_debug_pdest),UVM_NONE)
        end

        if(this.io_commits_info_0_debug_otherPdest_0!=rhs_.io_commits_info_0_debug_otherPdest_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_debug_otherPdest_0=0x%0h while the rhs_.io_commits_info_0_debug_otherPdest_0=0x%0h",this.io_commits_info_0_debug_otherPdest_0,rhs_.io_commits_info_0_debug_otherPdest_0),UVM_NONE)
        end

        if(this.io_commits_info_0_debug_otherPdest_1!=rhs_.io_commits_info_0_debug_otherPdest_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_debug_otherPdest_1=0x%0h while the rhs_.io_commits_info_0_debug_otherPdest_1=0x%0h",this.io_commits_info_0_debug_otherPdest_1,rhs_.io_commits_info_0_debug_otherPdest_1),UVM_NONE)
        end

        if(this.io_commits_info_0_debug_otherPdest_2!=rhs_.io_commits_info_0_debug_otherPdest_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_debug_otherPdest_2=0x%0h while the rhs_.io_commits_info_0_debug_otherPdest_2=0x%0h",this.io_commits_info_0_debug_otherPdest_2,rhs_.io_commits_info_0_debug_otherPdest_2),UVM_NONE)
        end

        if(this.io_commits_info_0_debug_otherPdest_3!=rhs_.io_commits_info_0_debug_otherPdest_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_debug_otherPdest_3=0x%0h while the rhs_.io_commits_info_0_debug_otherPdest_3=0x%0h",this.io_commits_info_0_debug_otherPdest_3,rhs_.io_commits_info_0_debug_otherPdest_3),UVM_NONE)
        end

        if(this.io_commits_info_0_debug_otherPdest_4!=rhs_.io_commits_info_0_debug_otherPdest_4) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_debug_otherPdest_4=0x%0h while the rhs_.io_commits_info_0_debug_otherPdest_4=0x%0h",this.io_commits_info_0_debug_otherPdest_4,rhs_.io_commits_info_0_debug_otherPdest_4),UVM_NONE)
        end

        if(this.io_commits_info_0_debug_otherPdest_5!=rhs_.io_commits_info_0_debug_otherPdest_5) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_debug_otherPdest_5=0x%0h while the rhs_.io_commits_info_0_debug_otherPdest_5=0x%0h",this.io_commits_info_0_debug_otherPdest_5,rhs_.io_commits_info_0_debug_otherPdest_5),UVM_NONE)
        end

        if(this.io_commits_info_0_debug_otherPdest_6!=rhs_.io_commits_info_0_debug_otherPdest_6) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_debug_otherPdest_6=0x%0h while the rhs_.io_commits_info_0_debug_otherPdest_6=0x%0h",this.io_commits_info_0_debug_otherPdest_6,rhs_.io_commits_info_0_debug_otherPdest_6),UVM_NONE)
        end

        if(this.io_commits_info_0_debug_fuType!=rhs_.io_commits_info_0_debug_fuType) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_debug_fuType=0x%0h while the rhs_.io_commits_info_0_debug_fuType=0x%0h",this.io_commits_info_0_debug_fuType,rhs_.io_commits_info_0_debug_fuType),UVM_NONE)
        end

        if(this.io_commits_info_0_dirtyFs!=rhs_.io_commits_info_0_dirtyFs) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_dirtyFs=0x%0h while the rhs_.io_commits_info_0_dirtyFs=0x%0h",this.io_commits_info_0_dirtyFs,rhs_.io_commits_info_0_dirtyFs),UVM_NONE)
        end

        if(this.io_commits_info_0_dirtyVs!=rhs_.io_commits_info_0_dirtyVs) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_0_dirtyVs=0x%0h while the rhs_.io_commits_info_0_dirtyVs=0x%0h",this.io_commits_info_0_dirtyVs,rhs_.io_commits_info_0_dirtyVs),UVM_NONE)
        end

        if(this.io_commits_info_1_walk_v!=rhs_.io_commits_info_1_walk_v) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_walk_v=0x%0h while the rhs_.io_commits_info_1_walk_v=0x%0h",this.io_commits_info_1_walk_v,rhs_.io_commits_info_1_walk_v),UVM_NONE)
        end

        if(this.io_commits_info_1_commit_v!=rhs_.io_commits_info_1_commit_v) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_commit_v=0x%0h while the rhs_.io_commits_info_1_commit_v=0x%0h",this.io_commits_info_1_commit_v,rhs_.io_commits_info_1_commit_v),UVM_NONE)
        end

        if(this.io_commits_info_1_commit_w!=rhs_.io_commits_info_1_commit_w) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_commit_w=0x%0h while the rhs_.io_commits_info_1_commit_w=0x%0h",this.io_commits_info_1_commit_w,rhs_.io_commits_info_1_commit_w),UVM_NONE)
        end

        if(this.io_commits_info_1_realDestSize!=rhs_.io_commits_info_1_realDestSize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_realDestSize=0x%0h while the rhs_.io_commits_info_1_realDestSize=0x%0h",this.io_commits_info_1_realDestSize,rhs_.io_commits_info_1_realDestSize),UVM_NONE)
        end

        if(this.io_commits_info_1_interrupt_safe!=rhs_.io_commits_info_1_interrupt_safe) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_interrupt_safe=0x%0h while the rhs_.io_commits_info_1_interrupt_safe=0x%0h",this.io_commits_info_1_interrupt_safe,rhs_.io_commits_info_1_interrupt_safe),UVM_NONE)
        end

        if(this.io_commits_info_1_wflags!=rhs_.io_commits_info_1_wflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_wflags=0x%0h while the rhs_.io_commits_info_1_wflags=0x%0h",this.io_commits_info_1_wflags,rhs_.io_commits_info_1_wflags),UVM_NONE)
        end

        if(this.io_commits_info_1_fflags!=rhs_.io_commits_info_1_fflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_fflags=0x%0h while the rhs_.io_commits_info_1_fflags=0x%0h",this.io_commits_info_1_fflags,rhs_.io_commits_info_1_fflags),UVM_NONE)
        end

        if(this.io_commits_info_1_vxsat!=rhs_.io_commits_info_1_vxsat) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_vxsat=0x%0h while the rhs_.io_commits_info_1_vxsat=0x%0h",this.io_commits_info_1_vxsat,rhs_.io_commits_info_1_vxsat),UVM_NONE)
        end

        if(this.io_commits_info_1_isRVC!=rhs_.io_commits_info_1_isRVC) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_isRVC=0x%0h while the rhs_.io_commits_info_1_isRVC=0x%0h",this.io_commits_info_1_isRVC,rhs_.io_commits_info_1_isRVC),UVM_NONE)
        end

        if(this.io_commits_info_1_isVset!=rhs_.io_commits_info_1_isVset) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_isVset=0x%0h while the rhs_.io_commits_info_1_isVset=0x%0h",this.io_commits_info_1_isVset,rhs_.io_commits_info_1_isVset),UVM_NONE)
        end

        if(this.io_commits_info_1_isHls!=rhs_.io_commits_info_1_isHls) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_isHls=0x%0h while the rhs_.io_commits_info_1_isHls=0x%0h",this.io_commits_info_1_isHls,rhs_.io_commits_info_1_isHls),UVM_NONE)
        end

        if(this.io_commits_info_1_isVls!=rhs_.io_commits_info_1_isVls) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_isVls=0x%0h while the rhs_.io_commits_info_1_isVls=0x%0h",this.io_commits_info_1_isVls,rhs_.io_commits_info_1_isVls),UVM_NONE)
        end

        if(this.io_commits_info_1_vls!=rhs_.io_commits_info_1_vls) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_vls=0x%0h while the rhs_.io_commits_info_1_vls=0x%0h",this.io_commits_info_1_vls,rhs_.io_commits_info_1_vls),UVM_NONE)
        end

        if(this.io_commits_info_1_mmio!=rhs_.io_commits_info_1_mmio) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_mmio=0x%0h while the rhs_.io_commits_info_1_mmio=0x%0h",this.io_commits_info_1_mmio,rhs_.io_commits_info_1_mmio),UVM_NONE)
        end

        if(this.io_commits_info_1_commitType!=rhs_.io_commits_info_1_commitType) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_commitType=0x%0h while the rhs_.io_commits_info_1_commitType=0x%0h",this.io_commits_info_1_commitType,rhs_.io_commits_info_1_commitType),UVM_NONE)
        end

        if(this.io_commits_info_1_ftqIdx_flag!=rhs_.io_commits_info_1_ftqIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_ftqIdx_flag=0x%0h while the rhs_.io_commits_info_1_ftqIdx_flag=0x%0h",this.io_commits_info_1_ftqIdx_flag,rhs_.io_commits_info_1_ftqIdx_flag),UVM_NONE)
        end

        if(this.io_commits_info_1_ftqIdx_value!=rhs_.io_commits_info_1_ftqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_ftqIdx_value=0x%0h while the rhs_.io_commits_info_1_ftqIdx_value=0x%0h",this.io_commits_info_1_ftqIdx_value,rhs_.io_commits_info_1_ftqIdx_value),UVM_NONE)
        end

        if(this.io_commits_info_1_ftqOffset!=rhs_.io_commits_info_1_ftqOffset) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_ftqOffset=0x%0h while the rhs_.io_commits_info_1_ftqOffset=0x%0h",this.io_commits_info_1_ftqOffset,rhs_.io_commits_info_1_ftqOffset),UVM_NONE)
        end

        if(this.io_commits_info_1_instrSize!=rhs_.io_commits_info_1_instrSize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_instrSize=0x%0h while the rhs_.io_commits_info_1_instrSize=0x%0h",this.io_commits_info_1_instrSize,rhs_.io_commits_info_1_instrSize),UVM_NONE)
        end

        if(this.io_commits_info_1_fpWen!=rhs_.io_commits_info_1_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_fpWen=0x%0h while the rhs_.io_commits_info_1_fpWen=0x%0h",this.io_commits_info_1_fpWen,rhs_.io_commits_info_1_fpWen),UVM_NONE)
        end

        if(this.io_commits_info_1_rfWen!=rhs_.io_commits_info_1_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_rfWen=0x%0h while the rhs_.io_commits_info_1_rfWen=0x%0h",this.io_commits_info_1_rfWen,rhs_.io_commits_info_1_rfWen),UVM_NONE)
        end

        if(this.io_commits_info_1_needFlush!=rhs_.io_commits_info_1_needFlush) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_needFlush=0x%0h while the rhs_.io_commits_info_1_needFlush=0x%0h",this.io_commits_info_1_needFlush,rhs_.io_commits_info_1_needFlush),UVM_NONE)
        end

        if(this.io_commits_info_1_traceBlockInPipe_itype!=rhs_.io_commits_info_1_traceBlockInPipe_itype) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_traceBlockInPipe_itype=0x%0h while the rhs_.io_commits_info_1_traceBlockInPipe_itype=0x%0h",this.io_commits_info_1_traceBlockInPipe_itype,rhs_.io_commits_info_1_traceBlockInPipe_itype),UVM_NONE)
        end

        if(this.io_commits_info_1_traceBlockInPipe_iretire!=rhs_.io_commits_info_1_traceBlockInPipe_iretire) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_traceBlockInPipe_iretire=0x%0h while the rhs_.io_commits_info_1_traceBlockInPipe_iretire=0x%0h",this.io_commits_info_1_traceBlockInPipe_iretire,rhs_.io_commits_info_1_traceBlockInPipe_iretire),UVM_NONE)
        end

        if(this.io_commits_info_1_traceBlockInPipe_ilastsize!=rhs_.io_commits_info_1_traceBlockInPipe_ilastsize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_traceBlockInPipe_ilastsize=0x%0h while the rhs_.io_commits_info_1_traceBlockInPipe_ilastsize=0x%0h",this.io_commits_info_1_traceBlockInPipe_ilastsize,rhs_.io_commits_info_1_traceBlockInPipe_ilastsize),UVM_NONE)
        end

        if(this.io_commits_info_1_debug_pc!=rhs_.io_commits_info_1_debug_pc) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_debug_pc=0x%0h while the rhs_.io_commits_info_1_debug_pc=0x%0h",this.io_commits_info_1_debug_pc,rhs_.io_commits_info_1_debug_pc),UVM_NONE)
        end

        if(this.io_commits_info_1_debug_instr!=rhs_.io_commits_info_1_debug_instr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_debug_instr=0x%0h while the rhs_.io_commits_info_1_debug_instr=0x%0h",this.io_commits_info_1_debug_instr,rhs_.io_commits_info_1_debug_instr),UVM_NONE)
        end

        if(this.io_commits_info_1_debug_ldest!=rhs_.io_commits_info_1_debug_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_debug_ldest=0x%0h while the rhs_.io_commits_info_1_debug_ldest=0x%0h",this.io_commits_info_1_debug_ldest,rhs_.io_commits_info_1_debug_ldest),UVM_NONE)
        end

        if(this.io_commits_info_1_debug_pdest!=rhs_.io_commits_info_1_debug_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_debug_pdest=0x%0h while the rhs_.io_commits_info_1_debug_pdest=0x%0h",this.io_commits_info_1_debug_pdest,rhs_.io_commits_info_1_debug_pdest),UVM_NONE)
        end

        if(this.io_commits_info_1_debug_otherPdest_0!=rhs_.io_commits_info_1_debug_otherPdest_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_debug_otherPdest_0=0x%0h while the rhs_.io_commits_info_1_debug_otherPdest_0=0x%0h",this.io_commits_info_1_debug_otherPdest_0,rhs_.io_commits_info_1_debug_otherPdest_0),UVM_NONE)
        end

        if(this.io_commits_info_1_debug_otherPdest_1!=rhs_.io_commits_info_1_debug_otherPdest_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_debug_otherPdest_1=0x%0h while the rhs_.io_commits_info_1_debug_otherPdest_1=0x%0h",this.io_commits_info_1_debug_otherPdest_1,rhs_.io_commits_info_1_debug_otherPdest_1),UVM_NONE)
        end

        if(this.io_commits_info_1_debug_otherPdest_2!=rhs_.io_commits_info_1_debug_otherPdest_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_debug_otherPdest_2=0x%0h while the rhs_.io_commits_info_1_debug_otherPdest_2=0x%0h",this.io_commits_info_1_debug_otherPdest_2,rhs_.io_commits_info_1_debug_otherPdest_2),UVM_NONE)
        end

        if(this.io_commits_info_1_debug_otherPdest_3!=rhs_.io_commits_info_1_debug_otherPdest_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_debug_otherPdest_3=0x%0h while the rhs_.io_commits_info_1_debug_otherPdest_3=0x%0h",this.io_commits_info_1_debug_otherPdest_3,rhs_.io_commits_info_1_debug_otherPdest_3),UVM_NONE)
        end

        if(this.io_commits_info_1_debug_otherPdest_4!=rhs_.io_commits_info_1_debug_otherPdest_4) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_debug_otherPdest_4=0x%0h while the rhs_.io_commits_info_1_debug_otherPdest_4=0x%0h",this.io_commits_info_1_debug_otherPdest_4,rhs_.io_commits_info_1_debug_otherPdest_4),UVM_NONE)
        end

        if(this.io_commits_info_1_debug_otherPdest_5!=rhs_.io_commits_info_1_debug_otherPdest_5) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_debug_otherPdest_5=0x%0h while the rhs_.io_commits_info_1_debug_otherPdest_5=0x%0h",this.io_commits_info_1_debug_otherPdest_5,rhs_.io_commits_info_1_debug_otherPdest_5),UVM_NONE)
        end

        if(this.io_commits_info_1_debug_otherPdest_6!=rhs_.io_commits_info_1_debug_otherPdest_6) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_debug_otherPdest_6=0x%0h while the rhs_.io_commits_info_1_debug_otherPdest_6=0x%0h",this.io_commits_info_1_debug_otherPdest_6,rhs_.io_commits_info_1_debug_otherPdest_6),UVM_NONE)
        end

        if(this.io_commits_info_1_debug_fuType!=rhs_.io_commits_info_1_debug_fuType) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_debug_fuType=0x%0h while the rhs_.io_commits_info_1_debug_fuType=0x%0h",this.io_commits_info_1_debug_fuType,rhs_.io_commits_info_1_debug_fuType),UVM_NONE)
        end

        if(this.io_commits_info_1_dirtyFs!=rhs_.io_commits_info_1_dirtyFs) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_dirtyFs=0x%0h while the rhs_.io_commits_info_1_dirtyFs=0x%0h",this.io_commits_info_1_dirtyFs,rhs_.io_commits_info_1_dirtyFs),UVM_NONE)
        end

        if(this.io_commits_info_1_dirtyVs!=rhs_.io_commits_info_1_dirtyVs) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_1_dirtyVs=0x%0h while the rhs_.io_commits_info_1_dirtyVs=0x%0h",this.io_commits_info_1_dirtyVs,rhs_.io_commits_info_1_dirtyVs),UVM_NONE)
        end

        if(this.io_commits_info_2_walk_v!=rhs_.io_commits_info_2_walk_v) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_walk_v=0x%0h while the rhs_.io_commits_info_2_walk_v=0x%0h",this.io_commits_info_2_walk_v,rhs_.io_commits_info_2_walk_v),UVM_NONE)
        end

        if(this.io_commits_info_2_commit_v!=rhs_.io_commits_info_2_commit_v) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_commit_v=0x%0h while the rhs_.io_commits_info_2_commit_v=0x%0h",this.io_commits_info_2_commit_v,rhs_.io_commits_info_2_commit_v),UVM_NONE)
        end

        if(this.io_commits_info_2_commit_w!=rhs_.io_commits_info_2_commit_w) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_commit_w=0x%0h while the rhs_.io_commits_info_2_commit_w=0x%0h",this.io_commits_info_2_commit_w,rhs_.io_commits_info_2_commit_w),UVM_NONE)
        end

        if(this.io_commits_info_2_realDestSize!=rhs_.io_commits_info_2_realDestSize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_realDestSize=0x%0h while the rhs_.io_commits_info_2_realDestSize=0x%0h",this.io_commits_info_2_realDestSize,rhs_.io_commits_info_2_realDestSize),UVM_NONE)
        end

        if(this.io_commits_info_2_interrupt_safe!=rhs_.io_commits_info_2_interrupt_safe) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_interrupt_safe=0x%0h while the rhs_.io_commits_info_2_interrupt_safe=0x%0h",this.io_commits_info_2_interrupt_safe,rhs_.io_commits_info_2_interrupt_safe),UVM_NONE)
        end

        if(this.io_commits_info_2_wflags!=rhs_.io_commits_info_2_wflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_wflags=0x%0h while the rhs_.io_commits_info_2_wflags=0x%0h",this.io_commits_info_2_wflags,rhs_.io_commits_info_2_wflags),UVM_NONE)
        end

        if(this.io_commits_info_2_fflags!=rhs_.io_commits_info_2_fflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_fflags=0x%0h while the rhs_.io_commits_info_2_fflags=0x%0h",this.io_commits_info_2_fflags,rhs_.io_commits_info_2_fflags),UVM_NONE)
        end

        if(this.io_commits_info_2_vxsat!=rhs_.io_commits_info_2_vxsat) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_vxsat=0x%0h while the rhs_.io_commits_info_2_vxsat=0x%0h",this.io_commits_info_2_vxsat,rhs_.io_commits_info_2_vxsat),UVM_NONE)
        end

        if(this.io_commits_info_2_isRVC!=rhs_.io_commits_info_2_isRVC) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_isRVC=0x%0h while the rhs_.io_commits_info_2_isRVC=0x%0h",this.io_commits_info_2_isRVC,rhs_.io_commits_info_2_isRVC),UVM_NONE)
        end

        if(this.io_commits_info_2_isVset!=rhs_.io_commits_info_2_isVset) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_isVset=0x%0h while the rhs_.io_commits_info_2_isVset=0x%0h",this.io_commits_info_2_isVset,rhs_.io_commits_info_2_isVset),UVM_NONE)
        end

        if(this.io_commits_info_2_isHls!=rhs_.io_commits_info_2_isHls) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_isHls=0x%0h while the rhs_.io_commits_info_2_isHls=0x%0h",this.io_commits_info_2_isHls,rhs_.io_commits_info_2_isHls),UVM_NONE)
        end

        if(this.io_commits_info_2_isVls!=rhs_.io_commits_info_2_isVls) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_isVls=0x%0h while the rhs_.io_commits_info_2_isVls=0x%0h",this.io_commits_info_2_isVls,rhs_.io_commits_info_2_isVls),UVM_NONE)
        end

        if(this.io_commits_info_2_vls!=rhs_.io_commits_info_2_vls) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_vls=0x%0h while the rhs_.io_commits_info_2_vls=0x%0h",this.io_commits_info_2_vls,rhs_.io_commits_info_2_vls),UVM_NONE)
        end

        if(this.io_commits_info_2_mmio!=rhs_.io_commits_info_2_mmio) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_mmio=0x%0h while the rhs_.io_commits_info_2_mmio=0x%0h",this.io_commits_info_2_mmio,rhs_.io_commits_info_2_mmio),UVM_NONE)
        end

        if(this.io_commits_info_2_commitType!=rhs_.io_commits_info_2_commitType) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_commitType=0x%0h while the rhs_.io_commits_info_2_commitType=0x%0h",this.io_commits_info_2_commitType,rhs_.io_commits_info_2_commitType),UVM_NONE)
        end

        if(this.io_commits_info_2_ftqIdx_flag!=rhs_.io_commits_info_2_ftqIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_ftqIdx_flag=0x%0h while the rhs_.io_commits_info_2_ftqIdx_flag=0x%0h",this.io_commits_info_2_ftqIdx_flag,rhs_.io_commits_info_2_ftqIdx_flag),UVM_NONE)
        end

        if(this.io_commits_info_2_ftqIdx_value!=rhs_.io_commits_info_2_ftqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_ftqIdx_value=0x%0h while the rhs_.io_commits_info_2_ftqIdx_value=0x%0h",this.io_commits_info_2_ftqIdx_value,rhs_.io_commits_info_2_ftqIdx_value),UVM_NONE)
        end

        if(this.io_commits_info_2_ftqOffset!=rhs_.io_commits_info_2_ftqOffset) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_ftqOffset=0x%0h while the rhs_.io_commits_info_2_ftqOffset=0x%0h",this.io_commits_info_2_ftqOffset,rhs_.io_commits_info_2_ftqOffset),UVM_NONE)
        end

        if(this.io_commits_info_2_instrSize!=rhs_.io_commits_info_2_instrSize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_instrSize=0x%0h while the rhs_.io_commits_info_2_instrSize=0x%0h",this.io_commits_info_2_instrSize,rhs_.io_commits_info_2_instrSize),UVM_NONE)
        end

        if(this.io_commits_info_2_fpWen!=rhs_.io_commits_info_2_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_fpWen=0x%0h while the rhs_.io_commits_info_2_fpWen=0x%0h",this.io_commits_info_2_fpWen,rhs_.io_commits_info_2_fpWen),UVM_NONE)
        end

        if(this.io_commits_info_2_rfWen!=rhs_.io_commits_info_2_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_rfWen=0x%0h while the rhs_.io_commits_info_2_rfWen=0x%0h",this.io_commits_info_2_rfWen,rhs_.io_commits_info_2_rfWen),UVM_NONE)
        end

        if(this.io_commits_info_2_needFlush!=rhs_.io_commits_info_2_needFlush) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_needFlush=0x%0h while the rhs_.io_commits_info_2_needFlush=0x%0h",this.io_commits_info_2_needFlush,rhs_.io_commits_info_2_needFlush),UVM_NONE)
        end

        if(this.io_commits_info_2_traceBlockInPipe_itype!=rhs_.io_commits_info_2_traceBlockInPipe_itype) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_traceBlockInPipe_itype=0x%0h while the rhs_.io_commits_info_2_traceBlockInPipe_itype=0x%0h",this.io_commits_info_2_traceBlockInPipe_itype,rhs_.io_commits_info_2_traceBlockInPipe_itype),UVM_NONE)
        end

        if(this.io_commits_info_2_traceBlockInPipe_iretire!=rhs_.io_commits_info_2_traceBlockInPipe_iretire) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_traceBlockInPipe_iretire=0x%0h while the rhs_.io_commits_info_2_traceBlockInPipe_iretire=0x%0h",this.io_commits_info_2_traceBlockInPipe_iretire,rhs_.io_commits_info_2_traceBlockInPipe_iretire),UVM_NONE)
        end

        if(this.io_commits_info_2_traceBlockInPipe_ilastsize!=rhs_.io_commits_info_2_traceBlockInPipe_ilastsize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_traceBlockInPipe_ilastsize=0x%0h while the rhs_.io_commits_info_2_traceBlockInPipe_ilastsize=0x%0h",this.io_commits_info_2_traceBlockInPipe_ilastsize,rhs_.io_commits_info_2_traceBlockInPipe_ilastsize),UVM_NONE)
        end

        if(this.io_commits_info_2_debug_pc!=rhs_.io_commits_info_2_debug_pc) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_debug_pc=0x%0h while the rhs_.io_commits_info_2_debug_pc=0x%0h",this.io_commits_info_2_debug_pc,rhs_.io_commits_info_2_debug_pc),UVM_NONE)
        end

        if(this.io_commits_info_2_debug_instr!=rhs_.io_commits_info_2_debug_instr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_debug_instr=0x%0h while the rhs_.io_commits_info_2_debug_instr=0x%0h",this.io_commits_info_2_debug_instr,rhs_.io_commits_info_2_debug_instr),UVM_NONE)
        end

        if(this.io_commits_info_2_debug_ldest!=rhs_.io_commits_info_2_debug_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_debug_ldest=0x%0h while the rhs_.io_commits_info_2_debug_ldest=0x%0h",this.io_commits_info_2_debug_ldest,rhs_.io_commits_info_2_debug_ldest),UVM_NONE)
        end

        if(this.io_commits_info_2_debug_pdest!=rhs_.io_commits_info_2_debug_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_debug_pdest=0x%0h while the rhs_.io_commits_info_2_debug_pdest=0x%0h",this.io_commits_info_2_debug_pdest,rhs_.io_commits_info_2_debug_pdest),UVM_NONE)
        end

        if(this.io_commits_info_2_debug_otherPdest_0!=rhs_.io_commits_info_2_debug_otherPdest_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_debug_otherPdest_0=0x%0h while the rhs_.io_commits_info_2_debug_otherPdest_0=0x%0h",this.io_commits_info_2_debug_otherPdest_0,rhs_.io_commits_info_2_debug_otherPdest_0),UVM_NONE)
        end

        if(this.io_commits_info_2_debug_otherPdest_1!=rhs_.io_commits_info_2_debug_otherPdest_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_debug_otherPdest_1=0x%0h while the rhs_.io_commits_info_2_debug_otherPdest_1=0x%0h",this.io_commits_info_2_debug_otherPdest_1,rhs_.io_commits_info_2_debug_otherPdest_1),UVM_NONE)
        end

        if(this.io_commits_info_2_debug_otherPdest_2!=rhs_.io_commits_info_2_debug_otherPdest_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_debug_otherPdest_2=0x%0h while the rhs_.io_commits_info_2_debug_otherPdest_2=0x%0h",this.io_commits_info_2_debug_otherPdest_2,rhs_.io_commits_info_2_debug_otherPdest_2),UVM_NONE)
        end

        if(this.io_commits_info_2_debug_otherPdest_3!=rhs_.io_commits_info_2_debug_otherPdest_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_debug_otherPdest_3=0x%0h while the rhs_.io_commits_info_2_debug_otherPdest_3=0x%0h",this.io_commits_info_2_debug_otherPdest_3,rhs_.io_commits_info_2_debug_otherPdest_3),UVM_NONE)
        end

        if(this.io_commits_info_2_debug_otherPdest_4!=rhs_.io_commits_info_2_debug_otherPdest_4) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_debug_otherPdest_4=0x%0h while the rhs_.io_commits_info_2_debug_otherPdest_4=0x%0h",this.io_commits_info_2_debug_otherPdest_4,rhs_.io_commits_info_2_debug_otherPdest_4),UVM_NONE)
        end

        if(this.io_commits_info_2_debug_otherPdest_5!=rhs_.io_commits_info_2_debug_otherPdest_5) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_debug_otherPdest_5=0x%0h while the rhs_.io_commits_info_2_debug_otherPdest_5=0x%0h",this.io_commits_info_2_debug_otherPdest_5,rhs_.io_commits_info_2_debug_otherPdest_5),UVM_NONE)
        end

        if(this.io_commits_info_2_debug_otherPdest_6!=rhs_.io_commits_info_2_debug_otherPdest_6) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_debug_otherPdest_6=0x%0h while the rhs_.io_commits_info_2_debug_otherPdest_6=0x%0h",this.io_commits_info_2_debug_otherPdest_6,rhs_.io_commits_info_2_debug_otherPdest_6),UVM_NONE)
        end

        if(this.io_commits_info_2_debug_fuType!=rhs_.io_commits_info_2_debug_fuType) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_debug_fuType=0x%0h while the rhs_.io_commits_info_2_debug_fuType=0x%0h",this.io_commits_info_2_debug_fuType,rhs_.io_commits_info_2_debug_fuType),UVM_NONE)
        end

        if(this.io_commits_info_2_dirtyFs!=rhs_.io_commits_info_2_dirtyFs) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_dirtyFs=0x%0h while the rhs_.io_commits_info_2_dirtyFs=0x%0h",this.io_commits_info_2_dirtyFs,rhs_.io_commits_info_2_dirtyFs),UVM_NONE)
        end

        if(this.io_commits_info_2_dirtyVs!=rhs_.io_commits_info_2_dirtyVs) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_2_dirtyVs=0x%0h while the rhs_.io_commits_info_2_dirtyVs=0x%0h",this.io_commits_info_2_dirtyVs,rhs_.io_commits_info_2_dirtyVs),UVM_NONE)
        end

        if(this.io_commits_info_3_walk_v!=rhs_.io_commits_info_3_walk_v) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_walk_v=0x%0h while the rhs_.io_commits_info_3_walk_v=0x%0h",this.io_commits_info_3_walk_v,rhs_.io_commits_info_3_walk_v),UVM_NONE)
        end

        if(this.io_commits_info_3_commit_v!=rhs_.io_commits_info_3_commit_v) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_commit_v=0x%0h while the rhs_.io_commits_info_3_commit_v=0x%0h",this.io_commits_info_3_commit_v,rhs_.io_commits_info_3_commit_v),UVM_NONE)
        end

        if(this.io_commits_info_3_commit_w!=rhs_.io_commits_info_3_commit_w) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_commit_w=0x%0h while the rhs_.io_commits_info_3_commit_w=0x%0h",this.io_commits_info_3_commit_w,rhs_.io_commits_info_3_commit_w),UVM_NONE)
        end

        if(this.io_commits_info_3_realDestSize!=rhs_.io_commits_info_3_realDestSize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_realDestSize=0x%0h while the rhs_.io_commits_info_3_realDestSize=0x%0h",this.io_commits_info_3_realDestSize,rhs_.io_commits_info_3_realDestSize),UVM_NONE)
        end

        if(this.io_commits_info_3_interrupt_safe!=rhs_.io_commits_info_3_interrupt_safe) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_interrupt_safe=0x%0h while the rhs_.io_commits_info_3_interrupt_safe=0x%0h",this.io_commits_info_3_interrupt_safe,rhs_.io_commits_info_3_interrupt_safe),UVM_NONE)
        end

        if(this.io_commits_info_3_wflags!=rhs_.io_commits_info_3_wflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_wflags=0x%0h while the rhs_.io_commits_info_3_wflags=0x%0h",this.io_commits_info_3_wflags,rhs_.io_commits_info_3_wflags),UVM_NONE)
        end

        if(this.io_commits_info_3_fflags!=rhs_.io_commits_info_3_fflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_fflags=0x%0h while the rhs_.io_commits_info_3_fflags=0x%0h",this.io_commits_info_3_fflags,rhs_.io_commits_info_3_fflags),UVM_NONE)
        end

        if(this.io_commits_info_3_vxsat!=rhs_.io_commits_info_3_vxsat) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_vxsat=0x%0h while the rhs_.io_commits_info_3_vxsat=0x%0h",this.io_commits_info_3_vxsat,rhs_.io_commits_info_3_vxsat),UVM_NONE)
        end

        if(this.io_commits_info_3_isRVC!=rhs_.io_commits_info_3_isRVC) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_isRVC=0x%0h while the rhs_.io_commits_info_3_isRVC=0x%0h",this.io_commits_info_3_isRVC,rhs_.io_commits_info_3_isRVC),UVM_NONE)
        end

        if(this.io_commits_info_3_isVset!=rhs_.io_commits_info_3_isVset) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_isVset=0x%0h while the rhs_.io_commits_info_3_isVset=0x%0h",this.io_commits_info_3_isVset,rhs_.io_commits_info_3_isVset),UVM_NONE)
        end

        if(this.io_commits_info_3_isHls!=rhs_.io_commits_info_3_isHls) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_isHls=0x%0h while the rhs_.io_commits_info_3_isHls=0x%0h",this.io_commits_info_3_isHls,rhs_.io_commits_info_3_isHls),UVM_NONE)
        end

        if(this.io_commits_info_3_isVls!=rhs_.io_commits_info_3_isVls) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_isVls=0x%0h while the rhs_.io_commits_info_3_isVls=0x%0h",this.io_commits_info_3_isVls,rhs_.io_commits_info_3_isVls),UVM_NONE)
        end

        if(this.io_commits_info_3_vls!=rhs_.io_commits_info_3_vls) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_vls=0x%0h while the rhs_.io_commits_info_3_vls=0x%0h",this.io_commits_info_3_vls,rhs_.io_commits_info_3_vls),UVM_NONE)
        end

        if(this.io_commits_info_3_mmio!=rhs_.io_commits_info_3_mmio) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_mmio=0x%0h while the rhs_.io_commits_info_3_mmio=0x%0h",this.io_commits_info_3_mmio,rhs_.io_commits_info_3_mmio),UVM_NONE)
        end

        if(this.io_commits_info_3_commitType!=rhs_.io_commits_info_3_commitType) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_commitType=0x%0h while the rhs_.io_commits_info_3_commitType=0x%0h",this.io_commits_info_3_commitType,rhs_.io_commits_info_3_commitType),UVM_NONE)
        end

        if(this.io_commits_info_3_ftqIdx_flag!=rhs_.io_commits_info_3_ftqIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_ftqIdx_flag=0x%0h while the rhs_.io_commits_info_3_ftqIdx_flag=0x%0h",this.io_commits_info_3_ftqIdx_flag,rhs_.io_commits_info_3_ftqIdx_flag),UVM_NONE)
        end

        if(this.io_commits_info_3_ftqIdx_value!=rhs_.io_commits_info_3_ftqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_ftqIdx_value=0x%0h while the rhs_.io_commits_info_3_ftqIdx_value=0x%0h",this.io_commits_info_3_ftqIdx_value,rhs_.io_commits_info_3_ftqIdx_value),UVM_NONE)
        end

        if(this.io_commits_info_3_ftqOffset!=rhs_.io_commits_info_3_ftqOffset) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_ftqOffset=0x%0h while the rhs_.io_commits_info_3_ftqOffset=0x%0h",this.io_commits_info_3_ftqOffset,rhs_.io_commits_info_3_ftqOffset),UVM_NONE)
        end

        if(this.io_commits_info_3_instrSize!=rhs_.io_commits_info_3_instrSize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_instrSize=0x%0h while the rhs_.io_commits_info_3_instrSize=0x%0h",this.io_commits_info_3_instrSize,rhs_.io_commits_info_3_instrSize),UVM_NONE)
        end

        if(this.io_commits_info_3_fpWen!=rhs_.io_commits_info_3_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_fpWen=0x%0h while the rhs_.io_commits_info_3_fpWen=0x%0h",this.io_commits_info_3_fpWen,rhs_.io_commits_info_3_fpWen),UVM_NONE)
        end

        if(this.io_commits_info_3_rfWen!=rhs_.io_commits_info_3_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_rfWen=0x%0h while the rhs_.io_commits_info_3_rfWen=0x%0h",this.io_commits_info_3_rfWen,rhs_.io_commits_info_3_rfWen),UVM_NONE)
        end

        if(this.io_commits_info_3_needFlush!=rhs_.io_commits_info_3_needFlush) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_needFlush=0x%0h while the rhs_.io_commits_info_3_needFlush=0x%0h",this.io_commits_info_3_needFlush,rhs_.io_commits_info_3_needFlush),UVM_NONE)
        end

        if(this.io_commits_info_3_traceBlockInPipe_itype!=rhs_.io_commits_info_3_traceBlockInPipe_itype) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_traceBlockInPipe_itype=0x%0h while the rhs_.io_commits_info_3_traceBlockInPipe_itype=0x%0h",this.io_commits_info_3_traceBlockInPipe_itype,rhs_.io_commits_info_3_traceBlockInPipe_itype),UVM_NONE)
        end

        if(this.io_commits_info_3_traceBlockInPipe_iretire!=rhs_.io_commits_info_3_traceBlockInPipe_iretire) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_traceBlockInPipe_iretire=0x%0h while the rhs_.io_commits_info_3_traceBlockInPipe_iretire=0x%0h",this.io_commits_info_3_traceBlockInPipe_iretire,rhs_.io_commits_info_3_traceBlockInPipe_iretire),UVM_NONE)
        end

        if(this.io_commits_info_3_traceBlockInPipe_ilastsize!=rhs_.io_commits_info_3_traceBlockInPipe_ilastsize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_traceBlockInPipe_ilastsize=0x%0h while the rhs_.io_commits_info_3_traceBlockInPipe_ilastsize=0x%0h",this.io_commits_info_3_traceBlockInPipe_ilastsize,rhs_.io_commits_info_3_traceBlockInPipe_ilastsize),UVM_NONE)
        end

        if(this.io_commits_info_3_debug_pc!=rhs_.io_commits_info_3_debug_pc) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_debug_pc=0x%0h while the rhs_.io_commits_info_3_debug_pc=0x%0h",this.io_commits_info_3_debug_pc,rhs_.io_commits_info_3_debug_pc),UVM_NONE)
        end

        if(this.io_commits_info_3_debug_instr!=rhs_.io_commits_info_3_debug_instr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_debug_instr=0x%0h while the rhs_.io_commits_info_3_debug_instr=0x%0h",this.io_commits_info_3_debug_instr,rhs_.io_commits_info_3_debug_instr),UVM_NONE)
        end

        if(this.io_commits_info_3_debug_ldest!=rhs_.io_commits_info_3_debug_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_debug_ldest=0x%0h while the rhs_.io_commits_info_3_debug_ldest=0x%0h",this.io_commits_info_3_debug_ldest,rhs_.io_commits_info_3_debug_ldest),UVM_NONE)
        end

        if(this.io_commits_info_3_debug_pdest!=rhs_.io_commits_info_3_debug_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_debug_pdest=0x%0h while the rhs_.io_commits_info_3_debug_pdest=0x%0h",this.io_commits_info_3_debug_pdest,rhs_.io_commits_info_3_debug_pdest),UVM_NONE)
        end

        if(this.io_commits_info_3_debug_otherPdest_0!=rhs_.io_commits_info_3_debug_otherPdest_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_debug_otherPdest_0=0x%0h while the rhs_.io_commits_info_3_debug_otherPdest_0=0x%0h",this.io_commits_info_3_debug_otherPdest_0,rhs_.io_commits_info_3_debug_otherPdest_0),UVM_NONE)
        end

        if(this.io_commits_info_3_debug_otherPdest_1!=rhs_.io_commits_info_3_debug_otherPdest_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_debug_otherPdest_1=0x%0h while the rhs_.io_commits_info_3_debug_otherPdest_1=0x%0h",this.io_commits_info_3_debug_otherPdest_1,rhs_.io_commits_info_3_debug_otherPdest_1),UVM_NONE)
        end

        if(this.io_commits_info_3_debug_otherPdest_2!=rhs_.io_commits_info_3_debug_otherPdest_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_debug_otherPdest_2=0x%0h while the rhs_.io_commits_info_3_debug_otherPdest_2=0x%0h",this.io_commits_info_3_debug_otherPdest_2,rhs_.io_commits_info_3_debug_otherPdest_2),UVM_NONE)
        end

        if(this.io_commits_info_3_debug_otherPdest_3!=rhs_.io_commits_info_3_debug_otherPdest_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_debug_otherPdest_3=0x%0h while the rhs_.io_commits_info_3_debug_otherPdest_3=0x%0h",this.io_commits_info_3_debug_otherPdest_3,rhs_.io_commits_info_3_debug_otherPdest_3),UVM_NONE)
        end

        if(this.io_commits_info_3_debug_otherPdest_4!=rhs_.io_commits_info_3_debug_otherPdest_4) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_debug_otherPdest_4=0x%0h while the rhs_.io_commits_info_3_debug_otherPdest_4=0x%0h",this.io_commits_info_3_debug_otherPdest_4,rhs_.io_commits_info_3_debug_otherPdest_4),UVM_NONE)
        end

        if(this.io_commits_info_3_debug_otherPdest_5!=rhs_.io_commits_info_3_debug_otherPdest_5) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_debug_otherPdest_5=0x%0h while the rhs_.io_commits_info_3_debug_otherPdest_5=0x%0h",this.io_commits_info_3_debug_otherPdest_5,rhs_.io_commits_info_3_debug_otherPdest_5),UVM_NONE)
        end

        if(this.io_commits_info_3_debug_otherPdest_6!=rhs_.io_commits_info_3_debug_otherPdest_6) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_debug_otherPdest_6=0x%0h while the rhs_.io_commits_info_3_debug_otherPdest_6=0x%0h",this.io_commits_info_3_debug_otherPdest_6,rhs_.io_commits_info_3_debug_otherPdest_6),UVM_NONE)
        end

        if(this.io_commits_info_3_debug_fuType!=rhs_.io_commits_info_3_debug_fuType) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_debug_fuType=0x%0h while the rhs_.io_commits_info_3_debug_fuType=0x%0h",this.io_commits_info_3_debug_fuType,rhs_.io_commits_info_3_debug_fuType),UVM_NONE)
        end

        if(this.io_commits_info_3_dirtyFs!=rhs_.io_commits_info_3_dirtyFs) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_dirtyFs=0x%0h while the rhs_.io_commits_info_3_dirtyFs=0x%0h",this.io_commits_info_3_dirtyFs,rhs_.io_commits_info_3_dirtyFs),UVM_NONE)
        end

        if(this.io_commits_info_3_dirtyVs!=rhs_.io_commits_info_3_dirtyVs) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_3_dirtyVs=0x%0h while the rhs_.io_commits_info_3_dirtyVs=0x%0h",this.io_commits_info_3_dirtyVs,rhs_.io_commits_info_3_dirtyVs),UVM_NONE)
        end

        if(this.io_commits_info_4_walk_v!=rhs_.io_commits_info_4_walk_v) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_walk_v=0x%0h while the rhs_.io_commits_info_4_walk_v=0x%0h",this.io_commits_info_4_walk_v,rhs_.io_commits_info_4_walk_v),UVM_NONE)
        end

        if(this.io_commits_info_4_commit_v!=rhs_.io_commits_info_4_commit_v) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_commit_v=0x%0h while the rhs_.io_commits_info_4_commit_v=0x%0h",this.io_commits_info_4_commit_v,rhs_.io_commits_info_4_commit_v),UVM_NONE)
        end

        if(this.io_commits_info_4_commit_w!=rhs_.io_commits_info_4_commit_w) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_commit_w=0x%0h while the rhs_.io_commits_info_4_commit_w=0x%0h",this.io_commits_info_4_commit_w,rhs_.io_commits_info_4_commit_w),UVM_NONE)
        end

        if(this.io_commits_info_4_realDestSize!=rhs_.io_commits_info_4_realDestSize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_realDestSize=0x%0h while the rhs_.io_commits_info_4_realDestSize=0x%0h",this.io_commits_info_4_realDestSize,rhs_.io_commits_info_4_realDestSize),UVM_NONE)
        end

        if(this.io_commits_info_4_interrupt_safe!=rhs_.io_commits_info_4_interrupt_safe) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_interrupt_safe=0x%0h while the rhs_.io_commits_info_4_interrupt_safe=0x%0h",this.io_commits_info_4_interrupt_safe,rhs_.io_commits_info_4_interrupt_safe),UVM_NONE)
        end

        if(this.io_commits_info_4_wflags!=rhs_.io_commits_info_4_wflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_wflags=0x%0h while the rhs_.io_commits_info_4_wflags=0x%0h",this.io_commits_info_4_wflags,rhs_.io_commits_info_4_wflags),UVM_NONE)
        end

        if(this.io_commits_info_4_fflags!=rhs_.io_commits_info_4_fflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_fflags=0x%0h while the rhs_.io_commits_info_4_fflags=0x%0h",this.io_commits_info_4_fflags,rhs_.io_commits_info_4_fflags),UVM_NONE)
        end

        if(this.io_commits_info_4_vxsat!=rhs_.io_commits_info_4_vxsat) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_vxsat=0x%0h while the rhs_.io_commits_info_4_vxsat=0x%0h",this.io_commits_info_4_vxsat,rhs_.io_commits_info_4_vxsat),UVM_NONE)
        end

        if(this.io_commits_info_4_isRVC!=rhs_.io_commits_info_4_isRVC) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_isRVC=0x%0h while the rhs_.io_commits_info_4_isRVC=0x%0h",this.io_commits_info_4_isRVC,rhs_.io_commits_info_4_isRVC),UVM_NONE)
        end

        if(this.io_commits_info_4_isVset!=rhs_.io_commits_info_4_isVset) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_isVset=0x%0h while the rhs_.io_commits_info_4_isVset=0x%0h",this.io_commits_info_4_isVset,rhs_.io_commits_info_4_isVset),UVM_NONE)
        end

        if(this.io_commits_info_4_isHls!=rhs_.io_commits_info_4_isHls) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_isHls=0x%0h while the rhs_.io_commits_info_4_isHls=0x%0h",this.io_commits_info_4_isHls,rhs_.io_commits_info_4_isHls),UVM_NONE)
        end

        if(this.io_commits_info_4_isVls!=rhs_.io_commits_info_4_isVls) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_isVls=0x%0h while the rhs_.io_commits_info_4_isVls=0x%0h",this.io_commits_info_4_isVls,rhs_.io_commits_info_4_isVls),UVM_NONE)
        end

        if(this.io_commits_info_4_vls!=rhs_.io_commits_info_4_vls) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_vls=0x%0h while the rhs_.io_commits_info_4_vls=0x%0h",this.io_commits_info_4_vls,rhs_.io_commits_info_4_vls),UVM_NONE)
        end

        if(this.io_commits_info_4_mmio!=rhs_.io_commits_info_4_mmio) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_mmio=0x%0h while the rhs_.io_commits_info_4_mmio=0x%0h",this.io_commits_info_4_mmio,rhs_.io_commits_info_4_mmio),UVM_NONE)
        end

        if(this.io_commits_info_4_commitType!=rhs_.io_commits_info_4_commitType) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_commitType=0x%0h while the rhs_.io_commits_info_4_commitType=0x%0h",this.io_commits_info_4_commitType,rhs_.io_commits_info_4_commitType),UVM_NONE)
        end

        if(this.io_commits_info_4_ftqIdx_flag!=rhs_.io_commits_info_4_ftqIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_ftqIdx_flag=0x%0h while the rhs_.io_commits_info_4_ftqIdx_flag=0x%0h",this.io_commits_info_4_ftqIdx_flag,rhs_.io_commits_info_4_ftqIdx_flag),UVM_NONE)
        end

        if(this.io_commits_info_4_ftqIdx_value!=rhs_.io_commits_info_4_ftqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_ftqIdx_value=0x%0h while the rhs_.io_commits_info_4_ftqIdx_value=0x%0h",this.io_commits_info_4_ftqIdx_value,rhs_.io_commits_info_4_ftqIdx_value),UVM_NONE)
        end

        if(this.io_commits_info_4_ftqOffset!=rhs_.io_commits_info_4_ftqOffset) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_ftqOffset=0x%0h while the rhs_.io_commits_info_4_ftqOffset=0x%0h",this.io_commits_info_4_ftqOffset,rhs_.io_commits_info_4_ftqOffset),UVM_NONE)
        end

        if(this.io_commits_info_4_instrSize!=rhs_.io_commits_info_4_instrSize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_instrSize=0x%0h while the rhs_.io_commits_info_4_instrSize=0x%0h",this.io_commits_info_4_instrSize,rhs_.io_commits_info_4_instrSize),UVM_NONE)
        end

        if(this.io_commits_info_4_fpWen!=rhs_.io_commits_info_4_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_fpWen=0x%0h while the rhs_.io_commits_info_4_fpWen=0x%0h",this.io_commits_info_4_fpWen,rhs_.io_commits_info_4_fpWen),UVM_NONE)
        end

        if(this.io_commits_info_4_rfWen!=rhs_.io_commits_info_4_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_rfWen=0x%0h while the rhs_.io_commits_info_4_rfWen=0x%0h",this.io_commits_info_4_rfWen,rhs_.io_commits_info_4_rfWen),UVM_NONE)
        end

        if(this.io_commits_info_4_needFlush!=rhs_.io_commits_info_4_needFlush) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_needFlush=0x%0h while the rhs_.io_commits_info_4_needFlush=0x%0h",this.io_commits_info_4_needFlush,rhs_.io_commits_info_4_needFlush),UVM_NONE)
        end

        if(this.io_commits_info_4_traceBlockInPipe_itype!=rhs_.io_commits_info_4_traceBlockInPipe_itype) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_traceBlockInPipe_itype=0x%0h while the rhs_.io_commits_info_4_traceBlockInPipe_itype=0x%0h",this.io_commits_info_4_traceBlockInPipe_itype,rhs_.io_commits_info_4_traceBlockInPipe_itype),UVM_NONE)
        end

        if(this.io_commits_info_4_traceBlockInPipe_iretire!=rhs_.io_commits_info_4_traceBlockInPipe_iretire) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_traceBlockInPipe_iretire=0x%0h while the rhs_.io_commits_info_4_traceBlockInPipe_iretire=0x%0h",this.io_commits_info_4_traceBlockInPipe_iretire,rhs_.io_commits_info_4_traceBlockInPipe_iretire),UVM_NONE)
        end

        if(this.io_commits_info_4_traceBlockInPipe_ilastsize!=rhs_.io_commits_info_4_traceBlockInPipe_ilastsize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_traceBlockInPipe_ilastsize=0x%0h while the rhs_.io_commits_info_4_traceBlockInPipe_ilastsize=0x%0h",this.io_commits_info_4_traceBlockInPipe_ilastsize,rhs_.io_commits_info_4_traceBlockInPipe_ilastsize),UVM_NONE)
        end

        if(this.io_commits_info_4_debug_pc!=rhs_.io_commits_info_4_debug_pc) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_debug_pc=0x%0h while the rhs_.io_commits_info_4_debug_pc=0x%0h",this.io_commits_info_4_debug_pc,rhs_.io_commits_info_4_debug_pc),UVM_NONE)
        end

        if(this.io_commits_info_4_debug_instr!=rhs_.io_commits_info_4_debug_instr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_debug_instr=0x%0h while the rhs_.io_commits_info_4_debug_instr=0x%0h",this.io_commits_info_4_debug_instr,rhs_.io_commits_info_4_debug_instr),UVM_NONE)
        end

        if(this.io_commits_info_4_debug_ldest!=rhs_.io_commits_info_4_debug_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_debug_ldest=0x%0h while the rhs_.io_commits_info_4_debug_ldest=0x%0h",this.io_commits_info_4_debug_ldest,rhs_.io_commits_info_4_debug_ldest),UVM_NONE)
        end

        if(this.io_commits_info_4_debug_pdest!=rhs_.io_commits_info_4_debug_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_debug_pdest=0x%0h while the rhs_.io_commits_info_4_debug_pdest=0x%0h",this.io_commits_info_4_debug_pdest,rhs_.io_commits_info_4_debug_pdest),UVM_NONE)
        end

        if(this.io_commits_info_4_debug_otherPdest_0!=rhs_.io_commits_info_4_debug_otherPdest_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_debug_otherPdest_0=0x%0h while the rhs_.io_commits_info_4_debug_otherPdest_0=0x%0h",this.io_commits_info_4_debug_otherPdest_0,rhs_.io_commits_info_4_debug_otherPdest_0),UVM_NONE)
        end

        if(this.io_commits_info_4_debug_otherPdest_1!=rhs_.io_commits_info_4_debug_otherPdest_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_debug_otherPdest_1=0x%0h while the rhs_.io_commits_info_4_debug_otherPdest_1=0x%0h",this.io_commits_info_4_debug_otherPdest_1,rhs_.io_commits_info_4_debug_otherPdest_1),UVM_NONE)
        end

        if(this.io_commits_info_4_debug_otherPdest_2!=rhs_.io_commits_info_4_debug_otherPdest_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_debug_otherPdest_2=0x%0h while the rhs_.io_commits_info_4_debug_otherPdest_2=0x%0h",this.io_commits_info_4_debug_otherPdest_2,rhs_.io_commits_info_4_debug_otherPdest_2),UVM_NONE)
        end

        if(this.io_commits_info_4_debug_otherPdest_3!=rhs_.io_commits_info_4_debug_otherPdest_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_debug_otherPdest_3=0x%0h while the rhs_.io_commits_info_4_debug_otherPdest_3=0x%0h",this.io_commits_info_4_debug_otherPdest_3,rhs_.io_commits_info_4_debug_otherPdest_3),UVM_NONE)
        end

        if(this.io_commits_info_4_debug_otherPdest_4!=rhs_.io_commits_info_4_debug_otherPdest_4) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_debug_otherPdest_4=0x%0h while the rhs_.io_commits_info_4_debug_otherPdest_4=0x%0h",this.io_commits_info_4_debug_otherPdest_4,rhs_.io_commits_info_4_debug_otherPdest_4),UVM_NONE)
        end

        if(this.io_commits_info_4_debug_otherPdest_5!=rhs_.io_commits_info_4_debug_otherPdest_5) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_debug_otherPdest_5=0x%0h while the rhs_.io_commits_info_4_debug_otherPdest_5=0x%0h",this.io_commits_info_4_debug_otherPdest_5,rhs_.io_commits_info_4_debug_otherPdest_5),UVM_NONE)
        end

        if(this.io_commits_info_4_debug_otherPdest_6!=rhs_.io_commits_info_4_debug_otherPdest_6) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_debug_otherPdest_6=0x%0h while the rhs_.io_commits_info_4_debug_otherPdest_6=0x%0h",this.io_commits_info_4_debug_otherPdest_6,rhs_.io_commits_info_4_debug_otherPdest_6),UVM_NONE)
        end

        if(this.io_commits_info_4_debug_fuType!=rhs_.io_commits_info_4_debug_fuType) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_debug_fuType=0x%0h while the rhs_.io_commits_info_4_debug_fuType=0x%0h",this.io_commits_info_4_debug_fuType,rhs_.io_commits_info_4_debug_fuType),UVM_NONE)
        end

        if(this.io_commits_info_4_dirtyFs!=rhs_.io_commits_info_4_dirtyFs) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_dirtyFs=0x%0h while the rhs_.io_commits_info_4_dirtyFs=0x%0h",this.io_commits_info_4_dirtyFs,rhs_.io_commits_info_4_dirtyFs),UVM_NONE)
        end

        if(this.io_commits_info_4_dirtyVs!=rhs_.io_commits_info_4_dirtyVs) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_4_dirtyVs=0x%0h while the rhs_.io_commits_info_4_dirtyVs=0x%0h",this.io_commits_info_4_dirtyVs,rhs_.io_commits_info_4_dirtyVs),UVM_NONE)
        end

        if(this.io_commits_info_5_walk_v!=rhs_.io_commits_info_5_walk_v) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_walk_v=0x%0h while the rhs_.io_commits_info_5_walk_v=0x%0h",this.io_commits_info_5_walk_v,rhs_.io_commits_info_5_walk_v),UVM_NONE)
        end

        if(this.io_commits_info_5_commit_v!=rhs_.io_commits_info_5_commit_v) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_commit_v=0x%0h while the rhs_.io_commits_info_5_commit_v=0x%0h",this.io_commits_info_5_commit_v,rhs_.io_commits_info_5_commit_v),UVM_NONE)
        end

        if(this.io_commits_info_5_commit_w!=rhs_.io_commits_info_5_commit_w) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_commit_w=0x%0h while the rhs_.io_commits_info_5_commit_w=0x%0h",this.io_commits_info_5_commit_w,rhs_.io_commits_info_5_commit_w),UVM_NONE)
        end

        if(this.io_commits_info_5_realDestSize!=rhs_.io_commits_info_5_realDestSize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_realDestSize=0x%0h while the rhs_.io_commits_info_5_realDestSize=0x%0h",this.io_commits_info_5_realDestSize,rhs_.io_commits_info_5_realDestSize),UVM_NONE)
        end

        if(this.io_commits_info_5_interrupt_safe!=rhs_.io_commits_info_5_interrupt_safe) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_interrupt_safe=0x%0h while the rhs_.io_commits_info_5_interrupt_safe=0x%0h",this.io_commits_info_5_interrupt_safe,rhs_.io_commits_info_5_interrupt_safe),UVM_NONE)
        end

        if(this.io_commits_info_5_wflags!=rhs_.io_commits_info_5_wflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_wflags=0x%0h while the rhs_.io_commits_info_5_wflags=0x%0h",this.io_commits_info_5_wflags,rhs_.io_commits_info_5_wflags),UVM_NONE)
        end

        if(this.io_commits_info_5_fflags!=rhs_.io_commits_info_5_fflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_fflags=0x%0h while the rhs_.io_commits_info_5_fflags=0x%0h",this.io_commits_info_5_fflags,rhs_.io_commits_info_5_fflags),UVM_NONE)
        end

        if(this.io_commits_info_5_vxsat!=rhs_.io_commits_info_5_vxsat) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_vxsat=0x%0h while the rhs_.io_commits_info_5_vxsat=0x%0h",this.io_commits_info_5_vxsat,rhs_.io_commits_info_5_vxsat),UVM_NONE)
        end

        if(this.io_commits_info_5_isRVC!=rhs_.io_commits_info_5_isRVC) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_isRVC=0x%0h while the rhs_.io_commits_info_5_isRVC=0x%0h",this.io_commits_info_5_isRVC,rhs_.io_commits_info_5_isRVC),UVM_NONE)
        end

        if(this.io_commits_info_5_isVset!=rhs_.io_commits_info_5_isVset) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_isVset=0x%0h while the rhs_.io_commits_info_5_isVset=0x%0h",this.io_commits_info_5_isVset,rhs_.io_commits_info_5_isVset),UVM_NONE)
        end

        if(this.io_commits_info_5_isHls!=rhs_.io_commits_info_5_isHls) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_isHls=0x%0h while the rhs_.io_commits_info_5_isHls=0x%0h",this.io_commits_info_5_isHls,rhs_.io_commits_info_5_isHls),UVM_NONE)
        end

        if(this.io_commits_info_5_isVls!=rhs_.io_commits_info_5_isVls) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_isVls=0x%0h while the rhs_.io_commits_info_5_isVls=0x%0h",this.io_commits_info_5_isVls,rhs_.io_commits_info_5_isVls),UVM_NONE)
        end

        if(this.io_commits_info_5_vls!=rhs_.io_commits_info_5_vls) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_vls=0x%0h while the rhs_.io_commits_info_5_vls=0x%0h",this.io_commits_info_5_vls,rhs_.io_commits_info_5_vls),UVM_NONE)
        end

        if(this.io_commits_info_5_mmio!=rhs_.io_commits_info_5_mmio) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_mmio=0x%0h while the rhs_.io_commits_info_5_mmio=0x%0h",this.io_commits_info_5_mmio,rhs_.io_commits_info_5_mmio),UVM_NONE)
        end

        if(this.io_commits_info_5_commitType!=rhs_.io_commits_info_5_commitType) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_commitType=0x%0h while the rhs_.io_commits_info_5_commitType=0x%0h",this.io_commits_info_5_commitType,rhs_.io_commits_info_5_commitType),UVM_NONE)
        end

        if(this.io_commits_info_5_ftqIdx_flag!=rhs_.io_commits_info_5_ftqIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_ftqIdx_flag=0x%0h while the rhs_.io_commits_info_5_ftqIdx_flag=0x%0h",this.io_commits_info_5_ftqIdx_flag,rhs_.io_commits_info_5_ftqIdx_flag),UVM_NONE)
        end

        if(this.io_commits_info_5_ftqIdx_value!=rhs_.io_commits_info_5_ftqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_ftqIdx_value=0x%0h while the rhs_.io_commits_info_5_ftqIdx_value=0x%0h",this.io_commits_info_5_ftqIdx_value,rhs_.io_commits_info_5_ftqIdx_value),UVM_NONE)
        end

        if(this.io_commits_info_5_ftqOffset!=rhs_.io_commits_info_5_ftqOffset) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_ftqOffset=0x%0h while the rhs_.io_commits_info_5_ftqOffset=0x%0h",this.io_commits_info_5_ftqOffset,rhs_.io_commits_info_5_ftqOffset),UVM_NONE)
        end

        if(this.io_commits_info_5_instrSize!=rhs_.io_commits_info_5_instrSize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_instrSize=0x%0h while the rhs_.io_commits_info_5_instrSize=0x%0h",this.io_commits_info_5_instrSize,rhs_.io_commits_info_5_instrSize),UVM_NONE)
        end

        if(this.io_commits_info_5_fpWen!=rhs_.io_commits_info_5_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_fpWen=0x%0h while the rhs_.io_commits_info_5_fpWen=0x%0h",this.io_commits_info_5_fpWen,rhs_.io_commits_info_5_fpWen),UVM_NONE)
        end

        if(this.io_commits_info_5_rfWen!=rhs_.io_commits_info_5_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_rfWen=0x%0h while the rhs_.io_commits_info_5_rfWen=0x%0h",this.io_commits_info_5_rfWen,rhs_.io_commits_info_5_rfWen),UVM_NONE)
        end

        if(this.io_commits_info_5_needFlush!=rhs_.io_commits_info_5_needFlush) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_needFlush=0x%0h while the rhs_.io_commits_info_5_needFlush=0x%0h",this.io_commits_info_5_needFlush,rhs_.io_commits_info_5_needFlush),UVM_NONE)
        end

        if(this.io_commits_info_5_traceBlockInPipe_itype!=rhs_.io_commits_info_5_traceBlockInPipe_itype) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_traceBlockInPipe_itype=0x%0h while the rhs_.io_commits_info_5_traceBlockInPipe_itype=0x%0h",this.io_commits_info_5_traceBlockInPipe_itype,rhs_.io_commits_info_5_traceBlockInPipe_itype),UVM_NONE)
        end

        if(this.io_commits_info_5_traceBlockInPipe_iretire!=rhs_.io_commits_info_5_traceBlockInPipe_iretire) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_traceBlockInPipe_iretire=0x%0h while the rhs_.io_commits_info_5_traceBlockInPipe_iretire=0x%0h",this.io_commits_info_5_traceBlockInPipe_iretire,rhs_.io_commits_info_5_traceBlockInPipe_iretire),UVM_NONE)
        end

        if(this.io_commits_info_5_traceBlockInPipe_ilastsize!=rhs_.io_commits_info_5_traceBlockInPipe_ilastsize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_traceBlockInPipe_ilastsize=0x%0h while the rhs_.io_commits_info_5_traceBlockInPipe_ilastsize=0x%0h",this.io_commits_info_5_traceBlockInPipe_ilastsize,rhs_.io_commits_info_5_traceBlockInPipe_ilastsize),UVM_NONE)
        end

        if(this.io_commits_info_5_debug_pc!=rhs_.io_commits_info_5_debug_pc) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_debug_pc=0x%0h while the rhs_.io_commits_info_5_debug_pc=0x%0h",this.io_commits_info_5_debug_pc,rhs_.io_commits_info_5_debug_pc),UVM_NONE)
        end

        if(this.io_commits_info_5_debug_instr!=rhs_.io_commits_info_5_debug_instr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_debug_instr=0x%0h while the rhs_.io_commits_info_5_debug_instr=0x%0h",this.io_commits_info_5_debug_instr,rhs_.io_commits_info_5_debug_instr),UVM_NONE)
        end

        if(this.io_commits_info_5_debug_ldest!=rhs_.io_commits_info_5_debug_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_debug_ldest=0x%0h while the rhs_.io_commits_info_5_debug_ldest=0x%0h",this.io_commits_info_5_debug_ldest,rhs_.io_commits_info_5_debug_ldest),UVM_NONE)
        end

        if(this.io_commits_info_5_debug_pdest!=rhs_.io_commits_info_5_debug_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_debug_pdest=0x%0h while the rhs_.io_commits_info_5_debug_pdest=0x%0h",this.io_commits_info_5_debug_pdest,rhs_.io_commits_info_5_debug_pdest),UVM_NONE)
        end

        if(this.io_commits_info_5_debug_otherPdest_0!=rhs_.io_commits_info_5_debug_otherPdest_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_debug_otherPdest_0=0x%0h while the rhs_.io_commits_info_5_debug_otherPdest_0=0x%0h",this.io_commits_info_5_debug_otherPdest_0,rhs_.io_commits_info_5_debug_otherPdest_0),UVM_NONE)
        end

        if(this.io_commits_info_5_debug_otherPdest_1!=rhs_.io_commits_info_5_debug_otherPdest_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_debug_otherPdest_1=0x%0h while the rhs_.io_commits_info_5_debug_otherPdest_1=0x%0h",this.io_commits_info_5_debug_otherPdest_1,rhs_.io_commits_info_5_debug_otherPdest_1),UVM_NONE)
        end

        if(this.io_commits_info_5_debug_otherPdest_2!=rhs_.io_commits_info_5_debug_otherPdest_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_debug_otherPdest_2=0x%0h while the rhs_.io_commits_info_5_debug_otherPdest_2=0x%0h",this.io_commits_info_5_debug_otherPdest_2,rhs_.io_commits_info_5_debug_otherPdest_2),UVM_NONE)
        end

        if(this.io_commits_info_5_debug_otherPdest_3!=rhs_.io_commits_info_5_debug_otherPdest_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_debug_otherPdest_3=0x%0h while the rhs_.io_commits_info_5_debug_otherPdest_3=0x%0h",this.io_commits_info_5_debug_otherPdest_3,rhs_.io_commits_info_5_debug_otherPdest_3),UVM_NONE)
        end

        if(this.io_commits_info_5_debug_otherPdest_4!=rhs_.io_commits_info_5_debug_otherPdest_4) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_debug_otherPdest_4=0x%0h while the rhs_.io_commits_info_5_debug_otherPdest_4=0x%0h",this.io_commits_info_5_debug_otherPdest_4,rhs_.io_commits_info_5_debug_otherPdest_4),UVM_NONE)
        end

        if(this.io_commits_info_5_debug_otherPdest_5!=rhs_.io_commits_info_5_debug_otherPdest_5) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_debug_otherPdest_5=0x%0h while the rhs_.io_commits_info_5_debug_otherPdest_5=0x%0h",this.io_commits_info_5_debug_otherPdest_5,rhs_.io_commits_info_5_debug_otherPdest_5),UVM_NONE)
        end

        if(this.io_commits_info_5_debug_otherPdest_6!=rhs_.io_commits_info_5_debug_otherPdest_6) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_debug_otherPdest_6=0x%0h while the rhs_.io_commits_info_5_debug_otherPdest_6=0x%0h",this.io_commits_info_5_debug_otherPdest_6,rhs_.io_commits_info_5_debug_otherPdest_6),UVM_NONE)
        end

        if(this.io_commits_info_5_debug_fuType!=rhs_.io_commits_info_5_debug_fuType) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_debug_fuType=0x%0h while the rhs_.io_commits_info_5_debug_fuType=0x%0h",this.io_commits_info_5_debug_fuType,rhs_.io_commits_info_5_debug_fuType),UVM_NONE)
        end

        if(this.io_commits_info_5_dirtyFs!=rhs_.io_commits_info_5_dirtyFs) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_dirtyFs=0x%0h while the rhs_.io_commits_info_5_dirtyFs=0x%0h",this.io_commits_info_5_dirtyFs,rhs_.io_commits_info_5_dirtyFs),UVM_NONE)
        end

        if(this.io_commits_info_5_dirtyVs!=rhs_.io_commits_info_5_dirtyVs) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_5_dirtyVs=0x%0h while the rhs_.io_commits_info_5_dirtyVs=0x%0h",this.io_commits_info_5_dirtyVs,rhs_.io_commits_info_5_dirtyVs),UVM_NONE)
        end

        if(this.io_commits_info_6_walk_v!=rhs_.io_commits_info_6_walk_v) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_walk_v=0x%0h while the rhs_.io_commits_info_6_walk_v=0x%0h",this.io_commits_info_6_walk_v,rhs_.io_commits_info_6_walk_v),UVM_NONE)
        end

        if(this.io_commits_info_6_commit_v!=rhs_.io_commits_info_6_commit_v) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_commit_v=0x%0h while the rhs_.io_commits_info_6_commit_v=0x%0h",this.io_commits_info_6_commit_v,rhs_.io_commits_info_6_commit_v),UVM_NONE)
        end

        if(this.io_commits_info_6_commit_w!=rhs_.io_commits_info_6_commit_w) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_commit_w=0x%0h while the rhs_.io_commits_info_6_commit_w=0x%0h",this.io_commits_info_6_commit_w,rhs_.io_commits_info_6_commit_w),UVM_NONE)
        end

        if(this.io_commits_info_6_realDestSize!=rhs_.io_commits_info_6_realDestSize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_realDestSize=0x%0h while the rhs_.io_commits_info_6_realDestSize=0x%0h",this.io_commits_info_6_realDestSize,rhs_.io_commits_info_6_realDestSize),UVM_NONE)
        end

        if(this.io_commits_info_6_interrupt_safe!=rhs_.io_commits_info_6_interrupt_safe) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_interrupt_safe=0x%0h while the rhs_.io_commits_info_6_interrupt_safe=0x%0h",this.io_commits_info_6_interrupt_safe,rhs_.io_commits_info_6_interrupt_safe),UVM_NONE)
        end

        if(this.io_commits_info_6_wflags!=rhs_.io_commits_info_6_wflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_wflags=0x%0h while the rhs_.io_commits_info_6_wflags=0x%0h",this.io_commits_info_6_wflags,rhs_.io_commits_info_6_wflags),UVM_NONE)
        end

        if(this.io_commits_info_6_fflags!=rhs_.io_commits_info_6_fflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_fflags=0x%0h while the rhs_.io_commits_info_6_fflags=0x%0h",this.io_commits_info_6_fflags,rhs_.io_commits_info_6_fflags),UVM_NONE)
        end

        if(this.io_commits_info_6_vxsat!=rhs_.io_commits_info_6_vxsat) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_vxsat=0x%0h while the rhs_.io_commits_info_6_vxsat=0x%0h",this.io_commits_info_6_vxsat,rhs_.io_commits_info_6_vxsat),UVM_NONE)
        end

        if(this.io_commits_info_6_isRVC!=rhs_.io_commits_info_6_isRVC) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_isRVC=0x%0h while the rhs_.io_commits_info_6_isRVC=0x%0h",this.io_commits_info_6_isRVC,rhs_.io_commits_info_6_isRVC),UVM_NONE)
        end

        if(this.io_commits_info_6_isVset!=rhs_.io_commits_info_6_isVset) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_isVset=0x%0h while the rhs_.io_commits_info_6_isVset=0x%0h",this.io_commits_info_6_isVset,rhs_.io_commits_info_6_isVset),UVM_NONE)
        end

        if(this.io_commits_info_6_isHls!=rhs_.io_commits_info_6_isHls) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_isHls=0x%0h while the rhs_.io_commits_info_6_isHls=0x%0h",this.io_commits_info_6_isHls,rhs_.io_commits_info_6_isHls),UVM_NONE)
        end

        if(this.io_commits_info_6_isVls!=rhs_.io_commits_info_6_isVls) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_isVls=0x%0h while the rhs_.io_commits_info_6_isVls=0x%0h",this.io_commits_info_6_isVls,rhs_.io_commits_info_6_isVls),UVM_NONE)
        end

        if(this.io_commits_info_6_vls!=rhs_.io_commits_info_6_vls) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_vls=0x%0h while the rhs_.io_commits_info_6_vls=0x%0h",this.io_commits_info_6_vls,rhs_.io_commits_info_6_vls),UVM_NONE)
        end

        if(this.io_commits_info_6_mmio!=rhs_.io_commits_info_6_mmio) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_mmio=0x%0h while the rhs_.io_commits_info_6_mmio=0x%0h",this.io_commits_info_6_mmio,rhs_.io_commits_info_6_mmio),UVM_NONE)
        end

        if(this.io_commits_info_6_commitType!=rhs_.io_commits_info_6_commitType) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_commitType=0x%0h while the rhs_.io_commits_info_6_commitType=0x%0h",this.io_commits_info_6_commitType,rhs_.io_commits_info_6_commitType),UVM_NONE)
        end

        if(this.io_commits_info_6_ftqIdx_flag!=rhs_.io_commits_info_6_ftqIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_ftqIdx_flag=0x%0h while the rhs_.io_commits_info_6_ftqIdx_flag=0x%0h",this.io_commits_info_6_ftqIdx_flag,rhs_.io_commits_info_6_ftqIdx_flag),UVM_NONE)
        end

        if(this.io_commits_info_6_ftqIdx_value!=rhs_.io_commits_info_6_ftqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_ftqIdx_value=0x%0h while the rhs_.io_commits_info_6_ftqIdx_value=0x%0h",this.io_commits_info_6_ftqIdx_value,rhs_.io_commits_info_6_ftqIdx_value),UVM_NONE)
        end

        if(this.io_commits_info_6_ftqOffset!=rhs_.io_commits_info_6_ftqOffset) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_ftqOffset=0x%0h while the rhs_.io_commits_info_6_ftqOffset=0x%0h",this.io_commits_info_6_ftqOffset,rhs_.io_commits_info_6_ftqOffset),UVM_NONE)
        end

        if(this.io_commits_info_6_instrSize!=rhs_.io_commits_info_6_instrSize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_instrSize=0x%0h while the rhs_.io_commits_info_6_instrSize=0x%0h",this.io_commits_info_6_instrSize,rhs_.io_commits_info_6_instrSize),UVM_NONE)
        end

        if(this.io_commits_info_6_fpWen!=rhs_.io_commits_info_6_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_fpWen=0x%0h while the rhs_.io_commits_info_6_fpWen=0x%0h",this.io_commits_info_6_fpWen,rhs_.io_commits_info_6_fpWen),UVM_NONE)
        end

        if(this.io_commits_info_6_rfWen!=rhs_.io_commits_info_6_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_rfWen=0x%0h while the rhs_.io_commits_info_6_rfWen=0x%0h",this.io_commits_info_6_rfWen,rhs_.io_commits_info_6_rfWen),UVM_NONE)
        end

        if(this.io_commits_info_6_needFlush!=rhs_.io_commits_info_6_needFlush) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_needFlush=0x%0h while the rhs_.io_commits_info_6_needFlush=0x%0h",this.io_commits_info_6_needFlush,rhs_.io_commits_info_6_needFlush),UVM_NONE)
        end

        if(this.io_commits_info_6_traceBlockInPipe_itype!=rhs_.io_commits_info_6_traceBlockInPipe_itype) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_traceBlockInPipe_itype=0x%0h while the rhs_.io_commits_info_6_traceBlockInPipe_itype=0x%0h",this.io_commits_info_6_traceBlockInPipe_itype,rhs_.io_commits_info_6_traceBlockInPipe_itype),UVM_NONE)
        end

        if(this.io_commits_info_6_traceBlockInPipe_iretire!=rhs_.io_commits_info_6_traceBlockInPipe_iretire) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_traceBlockInPipe_iretire=0x%0h while the rhs_.io_commits_info_6_traceBlockInPipe_iretire=0x%0h",this.io_commits_info_6_traceBlockInPipe_iretire,rhs_.io_commits_info_6_traceBlockInPipe_iretire),UVM_NONE)
        end

        if(this.io_commits_info_6_traceBlockInPipe_ilastsize!=rhs_.io_commits_info_6_traceBlockInPipe_ilastsize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_traceBlockInPipe_ilastsize=0x%0h while the rhs_.io_commits_info_6_traceBlockInPipe_ilastsize=0x%0h",this.io_commits_info_6_traceBlockInPipe_ilastsize,rhs_.io_commits_info_6_traceBlockInPipe_ilastsize),UVM_NONE)
        end

        if(this.io_commits_info_6_debug_pc!=rhs_.io_commits_info_6_debug_pc) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_debug_pc=0x%0h while the rhs_.io_commits_info_6_debug_pc=0x%0h",this.io_commits_info_6_debug_pc,rhs_.io_commits_info_6_debug_pc),UVM_NONE)
        end

        if(this.io_commits_info_6_debug_instr!=rhs_.io_commits_info_6_debug_instr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_debug_instr=0x%0h while the rhs_.io_commits_info_6_debug_instr=0x%0h",this.io_commits_info_6_debug_instr,rhs_.io_commits_info_6_debug_instr),UVM_NONE)
        end

        if(this.io_commits_info_6_debug_ldest!=rhs_.io_commits_info_6_debug_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_debug_ldest=0x%0h while the rhs_.io_commits_info_6_debug_ldest=0x%0h",this.io_commits_info_6_debug_ldest,rhs_.io_commits_info_6_debug_ldest),UVM_NONE)
        end

        if(this.io_commits_info_6_debug_pdest!=rhs_.io_commits_info_6_debug_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_debug_pdest=0x%0h while the rhs_.io_commits_info_6_debug_pdest=0x%0h",this.io_commits_info_6_debug_pdest,rhs_.io_commits_info_6_debug_pdest),UVM_NONE)
        end

        if(this.io_commits_info_6_debug_otherPdest_0!=rhs_.io_commits_info_6_debug_otherPdest_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_debug_otherPdest_0=0x%0h while the rhs_.io_commits_info_6_debug_otherPdest_0=0x%0h",this.io_commits_info_6_debug_otherPdest_0,rhs_.io_commits_info_6_debug_otherPdest_0),UVM_NONE)
        end

        if(this.io_commits_info_6_debug_otherPdest_1!=rhs_.io_commits_info_6_debug_otherPdest_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_debug_otherPdest_1=0x%0h while the rhs_.io_commits_info_6_debug_otherPdest_1=0x%0h",this.io_commits_info_6_debug_otherPdest_1,rhs_.io_commits_info_6_debug_otherPdest_1),UVM_NONE)
        end

        if(this.io_commits_info_6_debug_otherPdest_2!=rhs_.io_commits_info_6_debug_otherPdest_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_debug_otherPdest_2=0x%0h while the rhs_.io_commits_info_6_debug_otherPdest_2=0x%0h",this.io_commits_info_6_debug_otherPdest_2,rhs_.io_commits_info_6_debug_otherPdest_2),UVM_NONE)
        end

        if(this.io_commits_info_6_debug_otherPdest_3!=rhs_.io_commits_info_6_debug_otherPdest_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_debug_otherPdest_3=0x%0h while the rhs_.io_commits_info_6_debug_otherPdest_3=0x%0h",this.io_commits_info_6_debug_otherPdest_3,rhs_.io_commits_info_6_debug_otherPdest_3),UVM_NONE)
        end

        if(this.io_commits_info_6_debug_otherPdest_4!=rhs_.io_commits_info_6_debug_otherPdest_4) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_debug_otherPdest_4=0x%0h while the rhs_.io_commits_info_6_debug_otherPdest_4=0x%0h",this.io_commits_info_6_debug_otherPdest_4,rhs_.io_commits_info_6_debug_otherPdest_4),UVM_NONE)
        end

        if(this.io_commits_info_6_debug_otherPdest_5!=rhs_.io_commits_info_6_debug_otherPdest_5) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_debug_otherPdest_5=0x%0h while the rhs_.io_commits_info_6_debug_otherPdest_5=0x%0h",this.io_commits_info_6_debug_otherPdest_5,rhs_.io_commits_info_6_debug_otherPdest_5),UVM_NONE)
        end

        if(this.io_commits_info_6_debug_otherPdest_6!=rhs_.io_commits_info_6_debug_otherPdest_6) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_debug_otherPdest_6=0x%0h while the rhs_.io_commits_info_6_debug_otherPdest_6=0x%0h",this.io_commits_info_6_debug_otherPdest_6,rhs_.io_commits_info_6_debug_otherPdest_6),UVM_NONE)
        end

        if(this.io_commits_info_6_debug_fuType!=rhs_.io_commits_info_6_debug_fuType) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_debug_fuType=0x%0h while the rhs_.io_commits_info_6_debug_fuType=0x%0h",this.io_commits_info_6_debug_fuType,rhs_.io_commits_info_6_debug_fuType),UVM_NONE)
        end

        if(this.io_commits_info_6_dirtyFs!=rhs_.io_commits_info_6_dirtyFs) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_dirtyFs=0x%0h while the rhs_.io_commits_info_6_dirtyFs=0x%0h",this.io_commits_info_6_dirtyFs,rhs_.io_commits_info_6_dirtyFs),UVM_NONE)
        end

        if(this.io_commits_info_6_dirtyVs!=rhs_.io_commits_info_6_dirtyVs) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_6_dirtyVs=0x%0h while the rhs_.io_commits_info_6_dirtyVs=0x%0h",this.io_commits_info_6_dirtyVs,rhs_.io_commits_info_6_dirtyVs),UVM_NONE)
        end

        if(this.io_commits_info_7_walk_v!=rhs_.io_commits_info_7_walk_v) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_walk_v=0x%0h while the rhs_.io_commits_info_7_walk_v=0x%0h",this.io_commits_info_7_walk_v,rhs_.io_commits_info_7_walk_v),UVM_NONE)
        end

        if(this.io_commits_info_7_commit_v!=rhs_.io_commits_info_7_commit_v) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_commit_v=0x%0h while the rhs_.io_commits_info_7_commit_v=0x%0h",this.io_commits_info_7_commit_v,rhs_.io_commits_info_7_commit_v),UVM_NONE)
        end

        if(this.io_commits_info_7_commit_w!=rhs_.io_commits_info_7_commit_w) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_commit_w=0x%0h while the rhs_.io_commits_info_7_commit_w=0x%0h",this.io_commits_info_7_commit_w,rhs_.io_commits_info_7_commit_w),UVM_NONE)
        end

        if(this.io_commits_info_7_realDestSize!=rhs_.io_commits_info_7_realDestSize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_realDestSize=0x%0h while the rhs_.io_commits_info_7_realDestSize=0x%0h",this.io_commits_info_7_realDestSize,rhs_.io_commits_info_7_realDestSize),UVM_NONE)
        end

        if(this.io_commits_info_7_interrupt_safe!=rhs_.io_commits_info_7_interrupt_safe) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_interrupt_safe=0x%0h while the rhs_.io_commits_info_7_interrupt_safe=0x%0h",this.io_commits_info_7_interrupt_safe,rhs_.io_commits_info_7_interrupt_safe),UVM_NONE)
        end

        if(this.io_commits_info_7_wflags!=rhs_.io_commits_info_7_wflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_wflags=0x%0h while the rhs_.io_commits_info_7_wflags=0x%0h",this.io_commits_info_7_wflags,rhs_.io_commits_info_7_wflags),UVM_NONE)
        end

        if(this.io_commits_info_7_fflags!=rhs_.io_commits_info_7_fflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_fflags=0x%0h while the rhs_.io_commits_info_7_fflags=0x%0h",this.io_commits_info_7_fflags,rhs_.io_commits_info_7_fflags),UVM_NONE)
        end

        if(this.io_commits_info_7_vxsat!=rhs_.io_commits_info_7_vxsat) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_vxsat=0x%0h while the rhs_.io_commits_info_7_vxsat=0x%0h",this.io_commits_info_7_vxsat,rhs_.io_commits_info_7_vxsat),UVM_NONE)
        end

        if(this.io_commits_info_7_isRVC!=rhs_.io_commits_info_7_isRVC) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_isRVC=0x%0h while the rhs_.io_commits_info_7_isRVC=0x%0h",this.io_commits_info_7_isRVC,rhs_.io_commits_info_7_isRVC),UVM_NONE)
        end

        if(this.io_commits_info_7_isVset!=rhs_.io_commits_info_7_isVset) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_isVset=0x%0h while the rhs_.io_commits_info_7_isVset=0x%0h",this.io_commits_info_7_isVset,rhs_.io_commits_info_7_isVset),UVM_NONE)
        end

        if(this.io_commits_info_7_isHls!=rhs_.io_commits_info_7_isHls) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_isHls=0x%0h while the rhs_.io_commits_info_7_isHls=0x%0h",this.io_commits_info_7_isHls,rhs_.io_commits_info_7_isHls),UVM_NONE)
        end

        if(this.io_commits_info_7_isVls!=rhs_.io_commits_info_7_isVls) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_isVls=0x%0h while the rhs_.io_commits_info_7_isVls=0x%0h",this.io_commits_info_7_isVls,rhs_.io_commits_info_7_isVls),UVM_NONE)
        end

        if(this.io_commits_info_7_vls!=rhs_.io_commits_info_7_vls) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_vls=0x%0h while the rhs_.io_commits_info_7_vls=0x%0h",this.io_commits_info_7_vls,rhs_.io_commits_info_7_vls),UVM_NONE)
        end

        if(this.io_commits_info_7_mmio!=rhs_.io_commits_info_7_mmio) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_mmio=0x%0h while the rhs_.io_commits_info_7_mmio=0x%0h",this.io_commits_info_7_mmio,rhs_.io_commits_info_7_mmio),UVM_NONE)
        end

        if(this.io_commits_info_7_commitType!=rhs_.io_commits_info_7_commitType) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_commitType=0x%0h while the rhs_.io_commits_info_7_commitType=0x%0h",this.io_commits_info_7_commitType,rhs_.io_commits_info_7_commitType),UVM_NONE)
        end

        if(this.io_commits_info_7_ftqIdx_flag!=rhs_.io_commits_info_7_ftqIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_ftqIdx_flag=0x%0h while the rhs_.io_commits_info_7_ftqIdx_flag=0x%0h",this.io_commits_info_7_ftqIdx_flag,rhs_.io_commits_info_7_ftqIdx_flag),UVM_NONE)
        end

        if(this.io_commits_info_7_ftqIdx_value!=rhs_.io_commits_info_7_ftqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_ftqIdx_value=0x%0h while the rhs_.io_commits_info_7_ftqIdx_value=0x%0h",this.io_commits_info_7_ftqIdx_value,rhs_.io_commits_info_7_ftqIdx_value),UVM_NONE)
        end

        if(this.io_commits_info_7_ftqOffset!=rhs_.io_commits_info_7_ftqOffset) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_ftqOffset=0x%0h while the rhs_.io_commits_info_7_ftqOffset=0x%0h",this.io_commits_info_7_ftqOffset,rhs_.io_commits_info_7_ftqOffset),UVM_NONE)
        end

        if(this.io_commits_info_7_instrSize!=rhs_.io_commits_info_7_instrSize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_instrSize=0x%0h while the rhs_.io_commits_info_7_instrSize=0x%0h",this.io_commits_info_7_instrSize,rhs_.io_commits_info_7_instrSize),UVM_NONE)
        end

        if(this.io_commits_info_7_fpWen!=rhs_.io_commits_info_7_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_fpWen=0x%0h while the rhs_.io_commits_info_7_fpWen=0x%0h",this.io_commits_info_7_fpWen,rhs_.io_commits_info_7_fpWen),UVM_NONE)
        end

        if(this.io_commits_info_7_rfWen!=rhs_.io_commits_info_7_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_rfWen=0x%0h while the rhs_.io_commits_info_7_rfWen=0x%0h",this.io_commits_info_7_rfWen,rhs_.io_commits_info_7_rfWen),UVM_NONE)
        end

        if(this.io_commits_info_7_needFlush!=rhs_.io_commits_info_7_needFlush) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_needFlush=0x%0h while the rhs_.io_commits_info_7_needFlush=0x%0h",this.io_commits_info_7_needFlush,rhs_.io_commits_info_7_needFlush),UVM_NONE)
        end

        if(this.io_commits_info_7_traceBlockInPipe_itype!=rhs_.io_commits_info_7_traceBlockInPipe_itype) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_traceBlockInPipe_itype=0x%0h while the rhs_.io_commits_info_7_traceBlockInPipe_itype=0x%0h",this.io_commits_info_7_traceBlockInPipe_itype,rhs_.io_commits_info_7_traceBlockInPipe_itype),UVM_NONE)
        end

        if(this.io_commits_info_7_traceBlockInPipe_iretire!=rhs_.io_commits_info_7_traceBlockInPipe_iretire) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_traceBlockInPipe_iretire=0x%0h while the rhs_.io_commits_info_7_traceBlockInPipe_iretire=0x%0h",this.io_commits_info_7_traceBlockInPipe_iretire,rhs_.io_commits_info_7_traceBlockInPipe_iretire),UVM_NONE)
        end

        if(this.io_commits_info_7_traceBlockInPipe_ilastsize!=rhs_.io_commits_info_7_traceBlockInPipe_ilastsize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_traceBlockInPipe_ilastsize=0x%0h while the rhs_.io_commits_info_7_traceBlockInPipe_ilastsize=0x%0h",this.io_commits_info_7_traceBlockInPipe_ilastsize,rhs_.io_commits_info_7_traceBlockInPipe_ilastsize),UVM_NONE)
        end

        if(this.io_commits_info_7_debug_pc!=rhs_.io_commits_info_7_debug_pc) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_debug_pc=0x%0h while the rhs_.io_commits_info_7_debug_pc=0x%0h",this.io_commits_info_7_debug_pc,rhs_.io_commits_info_7_debug_pc),UVM_NONE)
        end

        if(this.io_commits_info_7_debug_instr!=rhs_.io_commits_info_7_debug_instr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_debug_instr=0x%0h while the rhs_.io_commits_info_7_debug_instr=0x%0h",this.io_commits_info_7_debug_instr,rhs_.io_commits_info_7_debug_instr),UVM_NONE)
        end

        if(this.io_commits_info_7_debug_ldest!=rhs_.io_commits_info_7_debug_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_debug_ldest=0x%0h while the rhs_.io_commits_info_7_debug_ldest=0x%0h",this.io_commits_info_7_debug_ldest,rhs_.io_commits_info_7_debug_ldest),UVM_NONE)
        end

        if(this.io_commits_info_7_debug_pdest!=rhs_.io_commits_info_7_debug_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_debug_pdest=0x%0h while the rhs_.io_commits_info_7_debug_pdest=0x%0h",this.io_commits_info_7_debug_pdest,rhs_.io_commits_info_7_debug_pdest),UVM_NONE)
        end

        if(this.io_commits_info_7_debug_otherPdest_0!=rhs_.io_commits_info_7_debug_otherPdest_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_debug_otherPdest_0=0x%0h while the rhs_.io_commits_info_7_debug_otherPdest_0=0x%0h",this.io_commits_info_7_debug_otherPdest_0,rhs_.io_commits_info_7_debug_otherPdest_0),UVM_NONE)
        end

        if(this.io_commits_info_7_debug_otherPdest_1!=rhs_.io_commits_info_7_debug_otherPdest_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_debug_otherPdest_1=0x%0h while the rhs_.io_commits_info_7_debug_otherPdest_1=0x%0h",this.io_commits_info_7_debug_otherPdest_1,rhs_.io_commits_info_7_debug_otherPdest_1),UVM_NONE)
        end

        if(this.io_commits_info_7_debug_otherPdest_2!=rhs_.io_commits_info_7_debug_otherPdest_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_debug_otherPdest_2=0x%0h while the rhs_.io_commits_info_7_debug_otherPdest_2=0x%0h",this.io_commits_info_7_debug_otherPdest_2,rhs_.io_commits_info_7_debug_otherPdest_2),UVM_NONE)
        end

        if(this.io_commits_info_7_debug_otherPdest_3!=rhs_.io_commits_info_7_debug_otherPdest_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_debug_otherPdest_3=0x%0h while the rhs_.io_commits_info_7_debug_otherPdest_3=0x%0h",this.io_commits_info_7_debug_otherPdest_3,rhs_.io_commits_info_7_debug_otherPdest_3),UVM_NONE)
        end

        if(this.io_commits_info_7_debug_otherPdest_4!=rhs_.io_commits_info_7_debug_otherPdest_4) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_debug_otherPdest_4=0x%0h while the rhs_.io_commits_info_7_debug_otherPdest_4=0x%0h",this.io_commits_info_7_debug_otherPdest_4,rhs_.io_commits_info_7_debug_otherPdest_4),UVM_NONE)
        end

        if(this.io_commits_info_7_debug_otherPdest_5!=rhs_.io_commits_info_7_debug_otherPdest_5) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_debug_otherPdest_5=0x%0h while the rhs_.io_commits_info_7_debug_otherPdest_5=0x%0h",this.io_commits_info_7_debug_otherPdest_5,rhs_.io_commits_info_7_debug_otherPdest_5),UVM_NONE)
        end

        if(this.io_commits_info_7_debug_otherPdest_6!=rhs_.io_commits_info_7_debug_otherPdest_6) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_debug_otherPdest_6=0x%0h while the rhs_.io_commits_info_7_debug_otherPdest_6=0x%0h",this.io_commits_info_7_debug_otherPdest_6,rhs_.io_commits_info_7_debug_otherPdest_6),UVM_NONE)
        end

        if(this.io_commits_info_7_debug_fuType!=rhs_.io_commits_info_7_debug_fuType) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_debug_fuType=0x%0h while the rhs_.io_commits_info_7_debug_fuType=0x%0h",this.io_commits_info_7_debug_fuType,rhs_.io_commits_info_7_debug_fuType),UVM_NONE)
        end

        if(this.io_commits_info_7_dirtyFs!=rhs_.io_commits_info_7_dirtyFs) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_dirtyFs=0x%0h while the rhs_.io_commits_info_7_dirtyFs=0x%0h",this.io_commits_info_7_dirtyFs,rhs_.io_commits_info_7_dirtyFs),UVM_NONE)
        end

        if(this.io_commits_info_7_dirtyVs!=rhs_.io_commits_info_7_dirtyVs) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_info_7_dirtyVs=0x%0h while the rhs_.io_commits_info_7_dirtyVs=0x%0h",this.io_commits_info_7_dirtyVs,rhs_.io_commits_info_7_dirtyVs),UVM_NONE)
        end

        if(this.io_commits_robIdx_0_flag!=rhs_.io_commits_robIdx_0_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_robIdx_0_flag=0x%0h while the rhs_.io_commits_robIdx_0_flag=0x%0h",this.io_commits_robIdx_0_flag,rhs_.io_commits_robIdx_0_flag),UVM_NONE)
        end

        if(this.io_commits_robIdx_0_value!=rhs_.io_commits_robIdx_0_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_robIdx_0_value=0x%0h while the rhs_.io_commits_robIdx_0_value=0x%0h",this.io_commits_robIdx_0_value,rhs_.io_commits_robIdx_0_value),UVM_NONE)
        end

        if(this.io_commits_robIdx_1_flag!=rhs_.io_commits_robIdx_1_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_robIdx_1_flag=0x%0h while the rhs_.io_commits_robIdx_1_flag=0x%0h",this.io_commits_robIdx_1_flag,rhs_.io_commits_robIdx_1_flag),UVM_NONE)
        end

        if(this.io_commits_robIdx_1_value!=rhs_.io_commits_robIdx_1_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_robIdx_1_value=0x%0h while the rhs_.io_commits_robIdx_1_value=0x%0h",this.io_commits_robIdx_1_value,rhs_.io_commits_robIdx_1_value),UVM_NONE)
        end

        if(this.io_commits_robIdx_2_flag!=rhs_.io_commits_robIdx_2_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_robIdx_2_flag=0x%0h while the rhs_.io_commits_robIdx_2_flag=0x%0h",this.io_commits_robIdx_2_flag,rhs_.io_commits_robIdx_2_flag),UVM_NONE)
        end

        if(this.io_commits_robIdx_2_value!=rhs_.io_commits_robIdx_2_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_robIdx_2_value=0x%0h while the rhs_.io_commits_robIdx_2_value=0x%0h",this.io_commits_robIdx_2_value,rhs_.io_commits_robIdx_2_value),UVM_NONE)
        end

        if(this.io_commits_robIdx_3_flag!=rhs_.io_commits_robIdx_3_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_robIdx_3_flag=0x%0h while the rhs_.io_commits_robIdx_3_flag=0x%0h",this.io_commits_robIdx_3_flag,rhs_.io_commits_robIdx_3_flag),UVM_NONE)
        end

        if(this.io_commits_robIdx_3_value!=rhs_.io_commits_robIdx_3_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_robIdx_3_value=0x%0h while the rhs_.io_commits_robIdx_3_value=0x%0h",this.io_commits_robIdx_3_value,rhs_.io_commits_robIdx_3_value),UVM_NONE)
        end

        if(this.io_commits_robIdx_4_flag!=rhs_.io_commits_robIdx_4_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_robIdx_4_flag=0x%0h while the rhs_.io_commits_robIdx_4_flag=0x%0h",this.io_commits_robIdx_4_flag,rhs_.io_commits_robIdx_4_flag),UVM_NONE)
        end

        if(this.io_commits_robIdx_4_value!=rhs_.io_commits_robIdx_4_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_robIdx_4_value=0x%0h while the rhs_.io_commits_robIdx_4_value=0x%0h",this.io_commits_robIdx_4_value,rhs_.io_commits_robIdx_4_value),UVM_NONE)
        end

        if(this.io_commits_robIdx_5_flag!=rhs_.io_commits_robIdx_5_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_robIdx_5_flag=0x%0h while the rhs_.io_commits_robIdx_5_flag=0x%0h",this.io_commits_robIdx_5_flag,rhs_.io_commits_robIdx_5_flag),UVM_NONE)
        end

        if(this.io_commits_robIdx_5_value!=rhs_.io_commits_robIdx_5_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_robIdx_5_value=0x%0h while the rhs_.io_commits_robIdx_5_value=0x%0h",this.io_commits_robIdx_5_value,rhs_.io_commits_robIdx_5_value),UVM_NONE)
        end

        if(this.io_commits_robIdx_6_flag!=rhs_.io_commits_robIdx_6_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_robIdx_6_flag=0x%0h while the rhs_.io_commits_robIdx_6_flag=0x%0h",this.io_commits_robIdx_6_flag,rhs_.io_commits_robIdx_6_flag),UVM_NONE)
        end

        if(this.io_commits_robIdx_6_value!=rhs_.io_commits_robIdx_6_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_robIdx_6_value=0x%0h while the rhs_.io_commits_robIdx_6_value=0x%0h",this.io_commits_robIdx_6_value,rhs_.io_commits_robIdx_6_value),UVM_NONE)
        end

        if(this.io_commits_robIdx_7_flag!=rhs_.io_commits_robIdx_7_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_robIdx_7_flag=0x%0h while the rhs_.io_commits_robIdx_7_flag=0x%0h",this.io_commits_robIdx_7_flag,rhs_.io_commits_robIdx_7_flag),UVM_NONE)
        end

        if(this.io_commits_robIdx_7_value!=rhs_.io_commits_robIdx_7_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_commits_robIdx_7_value=0x%0h while the rhs_.io_commits_robIdx_7_value=0x%0h",this.io_commits_robIdx_7_value,rhs_.io_commits_robIdx_7_value),UVM_NONE)
        end

        if(this.io_trace_blockCommit!=rhs_.io_trace_blockCommit) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_blockCommit=0x%0h while the rhs_.io_trace_blockCommit=0x%0h",this.io_trace_blockCommit,rhs_.io_trace_blockCommit),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_0_valid!=rhs_.io_trace_traceCommitInfo_blocks_0_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_0_valid=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_0_valid=0x%0h",this.io_trace_traceCommitInfo_blocks_0_valid,rhs_.io_trace_traceCommitInfo_blocks_0_valid),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value!=rhs_.io_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value=0x%0h",this.io_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value,rhs_.io_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_0_bits_ftqOffset!=rhs_.io_trace_traceCommitInfo_blocks_0_bits_ftqOffset) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_0_bits_ftqOffset=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_0_bits_ftqOffset=0x%0h",this.io_trace_traceCommitInfo_blocks_0_bits_ftqOffset,rhs_.io_trace_traceCommitInfo_blocks_0_bits_ftqOffset),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype!=rhs_.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype=0x%0h",this.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype,rhs_.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire!=rhs_.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire=0x%0h",this.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire,rhs_.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize!=rhs_.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize=0x%0h",this.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize,rhs_.io_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_1_valid!=rhs_.io_trace_traceCommitInfo_blocks_1_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_1_valid=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_1_valid=0x%0h",this.io_trace_traceCommitInfo_blocks_1_valid,rhs_.io_trace_traceCommitInfo_blocks_1_valid),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value!=rhs_.io_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value=0x%0h",this.io_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value,rhs_.io_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_1_bits_ftqOffset!=rhs_.io_trace_traceCommitInfo_blocks_1_bits_ftqOffset) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_1_bits_ftqOffset=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_1_bits_ftqOffset=0x%0h",this.io_trace_traceCommitInfo_blocks_1_bits_ftqOffset,rhs_.io_trace_traceCommitInfo_blocks_1_bits_ftqOffset),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype!=rhs_.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype=0x%0h",this.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype,rhs_.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire!=rhs_.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire=0x%0h",this.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire,rhs_.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize!=rhs_.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize=0x%0h",this.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize,rhs_.io_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_2_valid!=rhs_.io_trace_traceCommitInfo_blocks_2_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_2_valid=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_2_valid=0x%0h",this.io_trace_traceCommitInfo_blocks_2_valid,rhs_.io_trace_traceCommitInfo_blocks_2_valid),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value!=rhs_.io_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value=0x%0h",this.io_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value,rhs_.io_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_2_bits_ftqOffset!=rhs_.io_trace_traceCommitInfo_blocks_2_bits_ftqOffset) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_2_bits_ftqOffset=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_2_bits_ftqOffset=0x%0h",this.io_trace_traceCommitInfo_blocks_2_bits_ftqOffset,rhs_.io_trace_traceCommitInfo_blocks_2_bits_ftqOffset),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype!=rhs_.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype=0x%0h",this.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype,rhs_.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire!=rhs_.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire=0x%0h",this.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire,rhs_.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize!=rhs_.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize=0x%0h",this.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize,rhs_.io_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_3_valid!=rhs_.io_trace_traceCommitInfo_blocks_3_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_3_valid=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_3_valid=0x%0h",this.io_trace_traceCommitInfo_blocks_3_valid,rhs_.io_trace_traceCommitInfo_blocks_3_valid),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value!=rhs_.io_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value=0x%0h",this.io_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value,rhs_.io_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_3_bits_ftqOffset!=rhs_.io_trace_traceCommitInfo_blocks_3_bits_ftqOffset) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_3_bits_ftqOffset=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_3_bits_ftqOffset=0x%0h",this.io_trace_traceCommitInfo_blocks_3_bits_ftqOffset,rhs_.io_trace_traceCommitInfo_blocks_3_bits_ftqOffset),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype!=rhs_.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype=0x%0h",this.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype,rhs_.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire!=rhs_.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire=0x%0h",this.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire,rhs_.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize!=rhs_.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize=0x%0h",this.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize,rhs_.io_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_4_valid!=rhs_.io_trace_traceCommitInfo_blocks_4_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_4_valid=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_4_valid=0x%0h",this.io_trace_traceCommitInfo_blocks_4_valid,rhs_.io_trace_traceCommitInfo_blocks_4_valid),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value!=rhs_.io_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value=0x%0h",this.io_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value,rhs_.io_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_4_bits_ftqOffset!=rhs_.io_trace_traceCommitInfo_blocks_4_bits_ftqOffset) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_4_bits_ftqOffset=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_4_bits_ftqOffset=0x%0h",this.io_trace_traceCommitInfo_blocks_4_bits_ftqOffset,rhs_.io_trace_traceCommitInfo_blocks_4_bits_ftqOffset),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype!=rhs_.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype=0x%0h",this.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype,rhs_.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire!=rhs_.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire=0x%0h",this.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire,rhs_.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize!=rhs_.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize=0x%0h",this.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize,rhs_.io_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_5_valid!=rhs_.io_trace_traceCommitInfo_blocks_5_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_5_valid=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_5_valid=0x%0h",this.io_trace_traceCommitInfo_blocks_5_valid,rhs_.io_trace_traceCommitInfo_blocks_5_valid),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value!=rhs_.io_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value=0x%0h",this.io_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value,rhs_.io_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_5_bits_ftqOffset!=rhs_.io_trace_traceCommitInfo_blocks_5_bits_ftqOffset) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_5_bits_ftqOffset=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_5_bits_ftqOffset=0x%0h",this.io_trace_traceCommitInfo_blocks_5_bits_ftqOffset,rhs_.io_trace_traceCommitInfo_blocks_5_bits_ftqOffset),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype!=rhs_.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype=0x%0h",this.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype,rhs_.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire!=rhs_.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire=0x%0h",this.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire,rhs_.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize!=rhs_.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize=0x%0h",this.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize,rhs_.io_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_6_valid!=rhs_.io_trace_traceCommitInfo_blocks_6_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_6_valid=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_6_valid=0x%0h",this.io_trace_traceCommitInfo_blocks_6_valid,rhs_.io_trace_traceCommitInfo_blocks_6_valid),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value!=rhs_.io_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value=0x%0h",this.io_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value,rhs_.io_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_6_bits_ftqOffset!=rhs_.io_trace_traceCommitInfo_blocks_6_bits_ftqOffset) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_6_bits_ftqOffset=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_6_bits_ftqOffset=0x%0h",this.io_trace_traceCommitInfo_blocks_6_bits_ftqOffset,rhs_.io_trace_traceCommitInfo_blocks_6_bits_ftqOffset),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype!=rhs_.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype=0x%0h",this.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype,rhs_.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire!=rhs_.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire=0x%0h",this.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire,rhs_.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize!=rhs_.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize=0x%0h",this.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize,rhs_.io_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_7_valid!=rhs_.io_trace_traceCommitInfo_blocks_7_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_7_valid=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_7_valid=0x%0h",this.io_trace_traceCommitInfo_blocks_7_valid,rhs_.io_trace_traceCommitInfo_blocks_7_valid),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value!=rhs_.io_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value=0x%0h",this.io_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value,rhs_.io_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_7_bits_ftqOffset!=rhs_.io_trace_traceCommitInfo_blocks_7_bits_ftqOffset) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_7_bits_ftqOffset=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_7_bits_ftqOffset=0x%0h",this.io_trace_traceCommitInfo_blocks_7_bits_ftqOffset,rhs_.io_trace_traceCommitInfo_blocks_7_bits_ftqOffset),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype!=rhs_.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype=0x%0h",this.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype,rhs_.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire!=rhs_.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire=0x%0h",this.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire,rhs_.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire),UVM_NONE)
        end

        if(this.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize!=rhs_.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize=0x%0h while the rhs_.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize=0x%0h",this.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize,rhs_.io_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize),UVM_NONE)
        end

        if(this.io_rabCommits_isCommit!=rhs_.io_rabCommits_isCommit) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_isCommit=0x%0h while the rhs_.io_rabCommits_isCommit=0x%0h",this.io_rabCommits_isCommit,rhs_.io_rabCommits_isCommit),UVM_NONE)
        end

        if(this.io_rabCommits_commitValid_0!=rhs_.io_rabCommits_commitValid_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_commitValid_0=0x%0h while the rhs_.io_rabCommits_commitValid_0=0x%0h",this.io_rabCommits_commitValid_0,rhs_.io_rabCommits_commitValid_0),UVM_NONE)
        end

        if(this.io_rabCommits_commitValid_1!=rhs_.io_rabCommits_commitValid_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_commitValid_1=0x%0h while the rhs_.io_rabCommits_commitValid_1=0x%0h",this.io_rabCommits_commitValid_1,rhs_.io_rabCommits_commitValid_1),UVM_NONE)
        end

        if(this.io_rabCommits_commitValid_2!=rhs_.io_rabCommits_commitValid_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_commitValid_2=0x%0h while the rhs_.io_rabCommits_commitValid_2=0x%0h",this.io_rabCommits_commitValid_2,rhs_.io_rabCommits_commitValid_2),UVM_NONE)
        end

        if(this.io_rabCommits_commitValid_3!=rhs_.io_rabCommits_commitValid_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_commitValid_3=0x%0h while the rhs_.io_rabCommits_commitValid_3=0x%0h",this.io_rabCommits_commitValid_3,rhs_.io_rabCommits_commitValid_3),UVM_NONE)
        end

        if(this.io_rabCommits_commitValid_4!=rhs_.io_rabCommits_commitValid_4) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_commitValid_4=0x%0h while the rhs_.io_rabCommits_commitValid_4=0x%0h",this.io_rabCommits_commitValid_4,rhs_.io_rabCommits_commitValid_4),UVM_NONE)
        end

        if(this.io_rabCommits_commitValid_5!=rhs_.io_rabCommits_commitValid_5) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_commitValid_5=0x%0h while the rhs_.io_rabCommits_commitValid_5=0x%0h",this.io_rabCommits_commitValid_5,rhs_.io_rabCommits_commitValid_5),UVM_NONE)
        end

        if(this.io_rabCommits_isWalk!=rhs_.io_rabCommits_isWalk) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_isWalk=0x%0h while the rhs_.io_rabCommits_isWalk=0x%0h",this.io_rabCommits_isWalk,rhs_.io_rabCommits_isWalk),UVM_NONE)
        end

        if(this.io_rabCommits_walkValid_0!=rhs_.io_rabCommits_walkValid_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_walkValid_0=0x%0h while the rhs_.io_rabCommits_walkValid_0=0x%0h",this.io_rabCommits_walkValid_0,rhs_.io_rabCommits_walkValid_0),UVM_NONE)
        end

        if(this.io_rabCommits_walkValid_1!=rhs_.io_rabCommits_walkValid_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_walkValid_1=0x%0h while the rhs_.io_rabCommits_walkValid_1=0x%0h",this.io_rabCommits_walkValid_1,rhs_.io_rabCommits_walkValid_1),UVM_NONE)
        end

        if(this.io_rabCommits_walkValid_2!=rhs_.io_rabCommits_walkValid_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_walkValid_2=0x%0h while the rhs_.io_rabCommits_walkValid_2=0x%0h",this.io_rabCommits_walkValid_2,rhs_.io_rabCommits_walkValid_2),UVM_NONE)
        end

        if(this.io_rabCommits_walkValid_3!=rhs_.io_rabCommits_walkValid_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_walkValid_3=0x%0h while the rhs_.io_rabCommits_walkValid_3=0x%0h",this.io_rabCommits_walkValid_3,rhs_.io_rabCommits_walkValid_3),UVM_NONE)
        end

        if(this.io_rabCommits_walkValid_4!=rhs_.io_rabCommits_walkValid_4) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_walkValid_4=0x%0h while the rhs_.io_rabCommits_walkValid_4=0x%0h",this.io_rabCommits_walkValid_4,rhs_.io_rabCommits_walkValid_4),UVM_NONE)
        end

        if(this.io_rabCommits_walkValid_5!=rhs_.io_rabCommits_walkValid_5) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_walkValid_5=0x%0h while the rhs_.io_rabCommits_walkValid_5=0x%0h",this.io_rabCommits_walkValid_5,rhs_.io_rabCommits_walkValid_5),UVM_NONE)
        end

        if(this.io_rabCommits_info_0_ldest!=rhs_.io_rabCommits_info_0_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_0_ldest=0x%0h while the rhs_.io_rabCommits_info_0_ldest=0x%0h",this.io_rabCommits_info_0_ldest,rhs_.io_rabCommits_info_0_ldest),UVM_NONE)
        end

        if(this.io_rabCommits_info_0_pdest!=rhs_.io_rabCommits_info_0_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_0_pdest=0x%0h while the rhs_.io_rabCommits_info_0_pdest=0x%0h",this.io_rabCommits_info_0_pdest,rhs_.io_rabCommits_info_0_pdest),UVM_NONE)
        end

        if(this.io_rabCommits_info_0_rfWen!=rhs_.io_rabCommits_info_0_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_0_rfWen=0x%0h while the rhs_.io_rabCommits_info_0_rfWen=0x%0h",this.io_rabCommits_info_0_rfWen,rhs_.io_rabCommits_info_0_rfWen),UVM_NONE)
        end

        if(this.io_rabCommits_info_0_fpWen!=rhs_.io_rabCommits_info_0_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_0_fpWen=0x%0h while the rhs_.io_rabCommits_info_0_fpWen=0x%0h",this.io_rabCommits_info_0_fpWen,rhs_.io_rabCommits_info_0_fpWen),UVM_NONE)
        end

        if(this.io_rabCommits_info_0_vecWen!=rhs_.io_rabCommits_info_0_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_0_vecWen=0x%0h while the rhs_.io_rabCommits_info_0_vecWen=0x%0h",this.io_rabCommits_info_0_vecWen,rhs_.io_rabCommits_info_0_vecWen),UVM_NONE)
        end

        if(this.io_rabCommits_info_0_v0Wen!=rhs_.io_rabCommits_info_0_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_0_v0Wen=0x%0h while the rhs_.io_rabCommits_info_0_v0Wen=0x%0h",this.io_rabCommits_info_0_v0Wen,rhs_.io_rabCommits_info_0_v0Wen),UVM_NONE)
        end

        if(this.io_rabCommits_info_0_vlWen!=rhs_.io_rabCommits_info_0_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_0_vlWen=0x%0h while the rhs_.io_rabCommits_info_0_vlWen=0x%0h",this.io_rabCommits_info_0_vlWen,rhs_.io_rabCommits_info_0_vlWen),UVM_NONE)
        end

        if(this.io_rabCommits_info_0_isMove!=rhs_.io_rabCommits_info_0_isMove) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_0_isMove=0x%0h while the rhs_.io_rabCommits_info_0_isMove=0x%0h",this.io_rabCommits_info_0_isMove,rhs_.io_rabCommits_info_0_isMove),UVM_NONE)
        end

        if(this.io_rabCommits_info_1_ldest!=rhs_.io_rabCommits_info_1_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_1_ldest=0x%0h while the rhs_.io_rabCommits_info_1_ldest=0x%0h",this.io_rabCommits_info_1_ldest,rhs_.io_rabCommits_info_1_ldest),UVM_NONE)
        end

        if(this.io_rabCommits_info_1_pdest!=rhs_.io_rabCommits_info_1_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_1_pdest=0x%0h while the rhs_.io_rabCommits_info_1_pdest=0x%0h",this.io_rabCommits_info_1_pdest,rhs_.io_rabCommits_info_1_pdest),UVM_NONE)
        end

        if(this.io_rabCommits_info_1_rfWen!=rhs_.io_rabCommits_info_1_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_1_rfWen=0x%0h while the rhs_.io_rabCommits_info_1_rfWen=0x%0h",this.io_rabCommits_info_1_rfWen,rhs_.io_rabCommits_info_1_rfWen),UVM_NONE)
        end

        if(this.io_rabCommits_info_1_fpWen!=rhs_.io_rabCommits_info_1_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_1_fpWen=0x%0h while the rhs_.io_rabCommits_info_1_fpWen=0x%0h",this.io_rabCommits_info_1_fpWen,rhs_.io_rabCommits_info_1_fpWen),UVM_NONE)
        end

        if(this.io_rabCommits_info_1_vecWen!=rhs_.io_rabCommits_info_1_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_1_vecWen=0x%0h while the rhs_.io_rabCommits_info_1_vecWen=0x%0h",this.io_rabCommits_info_1_vecWen,rhs_.io_rabCommits_info_1_vecWen),UVM_NONE)
        end

        if(this.io_rabCommits_info_1_v0Wen!=rhs_.io_rabCommits_info_1_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_1_v0Wen=0x%0h while the rhs_.io_rabCommits_info_1_v0Wen=0x%0h",this.io_rabCommits_info_1_v0Wen,rhs_.io_rabCommits_info_1_v0Wen),UVM_NONE)
        end

        if(this.io_rabCommits_info_1_vlWen!=rhs_.io_rabCommits_info_1_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_1_vlWen=0x%0h while the rhs_.io_rabCommits_info_1_vlWen=0x%0h",this.io_rabCommits_info_1_vlWen,rhs_.io_rabCommits_info_1_vlWen),UVM_NONE)
        end

        if(this.io_rabCommits_info_1_isMove!=rhs_.io_rabCommits_info_1_isMove) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_1_isMove=0x%0h while the rhs_.io_rabCommits_info_1_isMove=0x%0h",this.io_rabCommits_info_1_isMove,rhs_.io_rabCommits_info_1_isMove),UVM_NONE)
        end

        if(this.io_rabCommits_info_2_ldest!=rhs_.io_rabCommits_info_2_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_2_ldest=0x%0h while the rhs_.io_rabCommits_info_2_ldest=0x%0h",this.io_rabCommits_info_2_ldest,rhs_.io_rabCommits_info_2_ldest),UVM_NONE)
        end

        if(this.io_rabCommits_info_2_pdest!=rhs_.io_rabCommits_info_2_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_2_pdest=0x%0h while the rhs_.io_rabCommits_info_2_pdest=0x%0h",this.io_rabCommits_info_2_pdest,rhs_.io_rabCommits_info_2_pdest),UVM_NONE)
        end

        if(this.io_rabCommits_info_2_rfWen!=rhs_.io_rabCommits_info_2_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_2_rfWen=0x%0h while the rhs_.io_rabCommits_info_2_rfWen=0x%0h",this.io_rabCommits_info_2_rfWen,rhs_.io_rabCommits_info_2_rfWen),UVM_NONE)
        end

        if(this.io_rabCommits_info_2_fpWen!=rhs_.io_rabCommits_info_2_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_2_fpWen=0x%0h while the rhs_.io_rabCommits_info_2_fpWen=0x%0h",this.io_rabCommits_info_2_fpWen,rhs_.io_rabCommits_info_2_fpWen),UVM_NONE)
        end

        if(this.io_rabCommits_info_2_vecWen!=rhs_.io_rabCommits_info_2_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_2_vecWen=0x%0h while the rhs_.io_rabCommits_info_2_vecWen=0x%0h",this.io_rabCommits_info_2_vecWen,rhs_.io_rabCommits_info_2_vecWen),UVM_NONE)
        end

        if(this.io_rabCommits_info_2_v0Wen!=rhs_.io_rabCommits_info_2_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_2_v0Wen=0x%0h while the rhs_.io_rabCommits_info_2_v0Wen=0x%0h",this.io_rabCommits_info_2_v0Wen,rhs_.io_rabCommits_info_2_v0Wen),UVM_NONE)
        end

        if(this.io_rabCommits_info_2_vlWen!=rhs_.io_rabCommits_info_2_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_2_vlWen=0x%0h while the rhs_.io_rabCommits_info_2_vlWen=0x%0h",this.io_rabCommits_info_2_vlWen,rhs_.io_rabCommits_info_2_vlWen),UVM_NONE)
        end

        if(this.io_rabCommits_info_2_isMove!=rhs_.io_rabCommits_info_2_isMove) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_2_isMove=0x%0h while the rhs_.io_rabCommits_info_2_isMove=0x%0h",this.io_rabCommits_info_2_isMove,rhs_.io_rabCommits_info_2_isMove),UVM_NONE)
        end

        if(this.io_rabCommits_info_3_ldest!=rhs_.io_rabCommits_info_3_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_3_ldest=0x%0h while the rhs_.io_rabCommits_info_3_ldest=0x%0h",this.io_rabCommits_info_3_ldest,rhs_.io_rabCommits_info_3_ldest),UVM_NONE)
        end

        if(this.io_rabCommits_info_3_pdest!=rhs_.io_rabCommits_info_3_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_3_pdest=0x%0h while the rhs_.io_rabCommits_info_3_pdest=0x%0h",this.io_rabCommits_info_3_pdest,rhs_.io_rabCommits_info_3_pdest),UVM_NONE)
        end

        if(this.io_rabCommits_info_3_rfWen!=rhs_.io_rabCommits_info_3_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_3_rfWen=0x%0h while the rhs_.io_rabCommits_info_3_rfWen=0x%0h",this.io_rabCommits_info_3_rfWen,rhs_.io_rabCommits_info_3_rfWen),UVM_NONE)
        end

        if(this.io_rabCommits_info_3_fpWen!=rhs_.io_rabCommits_info_3_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_3_fpWen=0x%0h while the rhs_.io_rabCommits_info_3_fpWen=0x%0h",this.io_rabCommits_info_3_fpWen,rhs_.io_rabCommits_info_3_fpWen),UVM_NONE)
        end

        if(this.io_rabCommits_info_3_vecWen!=rhs_.io_rabCommits_info_3_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_3_vecWen=0x%0h while the rhs_.io_rabCommits_info_3_vecWen=0x%0h",this.io_rabCommits_info_3_vecWen,rhs_.io_rabCommits_info_3_vecWen),UVM_NONE)
        end

        if(this.io_rabCommits_info_3_v0Wen!=rhs_.io_rabCommits_info_3_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_3_v0Wen=0x%0h while the rhs_.io_rabCommits_info_3_v0Wen=0x%0h",this.io_rabCommits_info_3_v0Wen,rhs_.io_rabCommits_info_3_v0Wen),UVM_NONE)
        end

        if(this.io_rabCommits_info_3_vlWen!=rhs_.io_rabCommits_info_3_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_3_vlWen=0x%0h while the rhs_.io_rabCommits_info_3_vlWen=0x%0h",this.io_rabCommits_info_3_vlWen,rhs_.io_rabCommits_info_3_vlWen),UVM_NONE)
        end

        if(this.io_rabCommits_info_3_isMove!=rhs_.io_rabCommits_info_3_isMove) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_3_isMove=0x%0h while the rhs_.io_rabCommits_info_3_isMove=0x%0h",this.io_rabCommits_info_3_isMove,rhs_.io_rabCommits_info_3_isMove),UVM_NONE)
        end

        if(this.io_rabCommits_info_4_ldest!=rhs_.io_rabCommits_info_4_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_4_ldest=0x%0h while the rhs_.io_rabCommits_info_4_ldest=0x%0h",this.io_rabCommits_info_4_ldest,rhs_.io_rabCommits_info_4_ldest),UVM_NONE)
        end

        if(this.io_rabCommits_info_4_pdest!=rhs_.io_rabCommits_info_4_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_4_pdest=0x%0h while the rhs_.io_rabCommits_info_4_pdest=0x%0h",this.io_rabCommits_info_4_pdest,rhs_.io_rabCommits_info_4_pdest),UVM_NONE)
        end

        if(this.io_rabCommits_info_4_rfWen!=rhs_.io_rabCommits_info_4_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_4_rfWen=0x%0h while the rhs_.io_rabCommits_info_4_rfWen=0x%0h",this.io_rabCommits_info_4_rfWen,rhs_.io_rabCommits_info_4_rfWen),UVM_NONE)
        end

        if(this.io_rabCommits_info_4_fpWen!=rhs_.io_rabCommits_info_4_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_4_fpWen=0x%0h while the rhs_.io_rabCommits_info_4_fpWen=0x%0h",this.io_rabCommits_info_4_fpWen,rhs_.io_rabCommits_info_4_fpWen),UVM_NONE)
        end

        if(this.io_rabCommits_info_4_vecWen!=rhs_.io_rabCommits_info_4_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_4_vecWen=0x%0h while the rhs_.io_rabCommits_info_4_vecWen=0x%0h",this.io_rabCommits_info_4_vecWen,rhs_.io_rabCommits_info_4_vecWen),UVM_NONE)
        end

        if(this.io_rabCommits_info_4_v0Wen!=rhs_.io_rabCommits_info_4_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_4_v0Wen=0x%0h while the rhs_.io_rabCommits_info_4_v0Wen=0x%0h",this.io_rabCommits_info_4_v0Wen,rhs_.io_rabCommits_info_4_v0Wen),UVM_NONE)
        end

        if(this.io_rabCommits_info_4_vlWen!=rhs_.io_rabCommits_info_4_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_4_vlWen=0x%0h while the rhs_.io_rabCommits_info_4_vlWen=0x%0h",this.io_rabCommits_info_4_vlWen,rhs_.io_rabCommits_info_4_vlWen),UVM_NONE)
        end

        if(this.io_rabCommits_info_4_isMove!=rhs_.io_rabCommits_info_4_isMove) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_4_isMove=0x%0h while the rhs_.io_rabCommits_info_4_isMove=0x%0h",this.io_rabCommits_info_4_isMove,rhs_.io_rabCommits_info_4_isMove),UVM_NONE)
        end

        if(this.io_rabCommits_info_5_ldest!=rhs_.io_rabCommits_info_5_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_5_ldest=0x%0h while the rhs_.io_rabCommits_info_5_ldest=0x%0h",this.io_rabCommits_info_5_ldest,rhs_.io_rabCommits_info_5_ldest),UVM_NONE)
        end

        if(this.io_rabCommits_info_5_pdest!=rhs_.io_rabCommits_info_5_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_5_pdest=0x%0h while the rhs_.io_rabCommits_info_5_pdest=0x%0h",this.io_rabCommits_info_5_pdest,rhs_.io_rabCommits_info_5_pdest),UVM_NONE)
        end

        if(this.io_rabCommits_info_5_rfWen!=rhs_.io_rabCommits_info_5_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_5_rfWen=0x%0h while the rhs_.io_rabCommits_info_5_rfWen=0x%0h",this.io_rabCommits_info_5_rfWen,rhs_.io_rabCommits_info_5_rfWen),UVM_NONE)
        end

        if(this.io_rabCommits_info_5_fpWen!=rhs_.io_rabCommits_info_5_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_5_fpWen=0x%0h while the rhs_.io_rabCommits_info_5_fpWen=0x%0h",this.io_rabCommits_info_5_fpWen,rhs_.io_rabCommits_info_5_fpWen),UVM_NONE)
        end

        if(this.io_rabCommits_info_5_vecWen!=rhs_.io_rabCommits_info_5_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_5_vecWen=0x%0h while the rhs_.io_rabCommits_info_5_vecWen=0x%0h",this.io_rabCommits_info_5_vecWen,rhs_.io_rabCommits_info_5_vecWen),UVM_NONE)
        end

        if(this.io_rabCommits_info_5_v0Wen!=rhs_.io_rabCommits_info_5_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_5_v0Wen=0x%0h while the rhs_.io_rabCommits_info_5_v0Wen=0x%0h",this.io_rabCommits_info_5_v0Wen,rhs_.io_rabCommits_info_5_v0Wen),UVM_NONE)
        end

        if(this.io_rabCommits_info_5_vlWen!=rhs_.io_rabCommits_info_5_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_5_vlWen=0x%0h while the rhs_.io_rabCommits_info_5_vlWen=0x%0h",this.io_rabCommits_info_5_vlWen,rhs_.io_rabCommits_info_5_vlWen),UVM_NONE)
        end

        if(this.io_rabCommits_info_5_isMove!=rhs_.io_rabCommits_info_5_isMove) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_rabCommits_info_5_isMove=0x%0h while the rhs_.io_rabCommits_info_5_isMove=0x%0h",this.io_rabCommits_info_5_isMove,rhs_.io_rabCommits_info_5_isMove),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_0!=rhs_.io_diffCommits_commitValid_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_0=0x%0h while the rhs_.io_diffCommits_commitValid_0=0x%0h",this.io_diffCommits_commitValid_0,rhs_.io_diffCommits_commitValid_0),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_1!=rhs_.io_diffCommits_commitValid_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_1=0x%0h while the rhs_.io_diffCommits_commitValid_1=0x%0h",this.io_diffCommits_commitValid_1,rhs_.io_diffCommits_commitValid_1),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_2!=rhs_.io_diffCommits_commitValid_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_2=0x%0h while the rhs_.io_diffCommits_commitValid_2=0x%0h",this.io_diffCommits_commitValid_2,rhs_.io_diffCommits_commitValid_2),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_3!=rhs_.io_diffCommits_commitValid_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_3=0x%0h while the rhs_.io_diffCommits_commitValid_3=0x%0h",this.io_diffCommits_commitValid_3,rhs_.io_diffCommits_commitValid_3),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_4!=rhs_.io_diffCommits_commitValid_4) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_4=0x%0h while the rhs_.io_diffCommits_commitValid_4=0x%0h",this.io_diffCommits_commitValid_4,rhs_.io_diffCommits_commitValid_4),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_5!=rhs_.io_diffCommits_commitValid_5) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_5=0x%0h while the rhs_.io_diffCommits_commitValid_5=0x%0h",this.io_diffCommits_commitValid_5,rhs_.io_diffCommits_commitValid_5),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_6!=rhs_.io_diffCommits_commitValid_6) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_6=0x%0h while the rhs_.io_diffCommits_commitValid_6=0x%0h",this.io_diffCommits_commitValid_6,rhs_.io_diffCommits_commitValid_6),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_7!=rhs_.io_diffCommits_commitValid_7) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_7=0x%0h while the rhs_.io_diffCommits_commitValid_7=0x%0h",this.io_diffCommits_commitValid_7,rhs_.io_diffCommits_commitValid_7),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_8!=rhs_.io_diffCommits_commitValid_8) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_8=0x%0h while the rhs_.io_diffCommits_commitValid_8=0x%0h",this.io_diffCommits_commitValid_8,rhs_.io_diffCommits_commitValid_8),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_9!=rhs_.io_diffCommits_commitValid_9) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_9=0x%0h while the rhs_.io_diffCommits_commitValid_9=0x%0h",this.io_diffCommits_commitValid_9,rhs_.io_diffCommits_commitValid_9),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_10!=rhs_.io_diffCommits_commitValid_10) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_10=0x%0h while the rhs_.io_diffCommits_commitValid_10=0x%0h",this.io_diffCommits_commitValid_10,rhs_.io_diffCommits_commitValid_10),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_11!=rhs_.io_diffCommits_commitValid_11) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_11=0x%0h while the rhs_.io_diffCommits_commitValid_11=0x%0h",this.io_diffCommits_commitValid_11,rhs_.io_diffCommits_commitValid_11),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_12!=rhs_.io_diffCommits_commitValid_12) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_12=0x%0h while the rhs_.io_diffCommits_commitValid_12=0x%0h",this.io_diffCommits_commitValid_12,rhs_.io_diffCommits_commitValid_12),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_13!=rhs_.io_diffCommits_commitValid_13) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_13=0x%0h while the rhs_.io_diffCommits_commitValid_13=0x%0h",this.io_diffCommits_commitValid_13,rhs_.io_diffCommits_commitValid_13),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_14!=rhs_.io_diffCommits_commitValid_14) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_14=0x%0h while the rhs_.io_diffCommits_commitValid_14=0x%0h",this.io_diffCommits_commitValid_14,rhs_.io_diffCommits_commitValid_14),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_15!=rhs_.io_diffCommits_commitValid_15) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_15=0x%0h while the rhs_.io_diffCommits_commitValid_15=0x%0h",this.io_diffCommits_commitValid_15,rhs_.io_diffCommits_commitValid_15),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_16!=rhs_.io_diffCommits_commitValid_16) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_16=0x%0h while the rhs_.io_diffCommits_commitValid_16=0x%0h",this.io_diffCommits_commitValid_16,rhs_.io_diffCommits_commitValid_16),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_17!=rhs_.io_diffCommits_commitValid_17) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_17=0x%0h while the rhs_.io_diffCommits_commitValid_17=0x%0h",this.io_diffCommits_commitValid_17,rhs_.io_diffCommits_commitValid_17),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_18!=rhs_.io_diffCommits_commitValid_18) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_18=0x%0h while the rhs_.io_diffCommits_commitValid_18=0x%0h",this.io_diffCommits_commitValid_18,rhs_.io_diffCommits_commitValid_18),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_19!=rhs_.io_diffCommits_commitValid_19) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_19=0x%0h while the rhs_.io_diffCommits_commitValid_19=0x%0h",this.io_diffCommits_commitValid_19,rhs_.io_diffCommits_commitValid_19),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_20!=rhs_.io_diffCommits_commitValid_20) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_20=0x%0h while the rhs_.io_diffCommits_commitValid_20=0x%0h",this.io_diffCommits_commitValid_20,rhs_.io_diffCommits_commitValid_20),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_21!=rhs_.io_diffCommits_commitValid_21) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_21=0x%0h while the rhs_.io_diffCommits_commitValid_21=0x%0h",this.io_diffCommits_commitValid_21,rhs_.io_diffCommits_commitValid_21),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_22!=rhs_.io_diffCommits_commitValid_22) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_22=0x%0h while the rhs_.io_diffCommits_commitValid_22=0x%0h",this.io_diffCommits_commitValid_22,rhs_.io_diffCommits_commitValid_22),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_23!=rhs_.io_diffCommits_commitValid_23) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_23=0x%0h while the rhs_.io_diffCommits_commitValid_23=0x%0h",this.io_diffCommits_commitValid_23,rhs_.io_diffCommits_commitValid_23),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_24!=rhs_.io_diffCommits_commitValid_24) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_24=0x%0h while the rhs_.io_diffCommits_commitValid_24=0x%0h",this.io_diffCommits_commitValid_24,rhs_.io_diffCommits_commitValid_24),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_25!=rhs_.io_diffCommits_commitValid_25) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_25=0x%0h while the rhs_.io_diffCommits_commitValid_25=0x%0h",this.io_diffCommits_commitValid_25,rhs_.io_diffCommits_commitValid_25),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_26!=rhs_.io_diffCommits_commitValid_26) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_26=0x%0h while the rhs_.io_diffCommits_commitValid_26=0x%0h",this.io_diffCommits_commitValid_26,rhs_.io_diffCommits_commitValid_26),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_27!=rhs_.io_diffCommits_commitValid_27) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_27=0x%0h while the rhs_.io_diffCommits_commitValid_27=0x%0h",this.io_diffCommits_commitValid_27,rhs_.io_diffCommits_commitValid_27),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_28!=rhs_.io_diffCommits_commitValid_28) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_28=0x%0h while the rhs_.io_diffCommits_commitValid_28=0x%0h",this.io_diffCommits_commitValid_28,rhs_.io_diffCommits_commitValid_28),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_29!=rhs_.io_diffCommits_commitValid_29) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_29=0x%0h while the rhs_.io_diffCommits_commitValid_29=0x%0h",this.io_diffCommits_commitValid_29,rhs_.io_diffCommits_commitValid_29),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_30!=rhs_.io_diffCommits_commitValid_30) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_30=0x%0h while the rhs_.io_diffCommits_commitValid_30=0x%0h",this.io_diffCommits_commitValid_30,rhs_.io_diffCommits_commitValid_30),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_31!=rhs_.io_diffCommits_commitValid_31) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_31=0x%0h while the rhs_.io_diffCommits_commitValid_31=0x%0h",this.io_diffCommits_commitValid_31,rhs_.io_diffCommits_commitValid_31),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_32!=rhs_.io_diffCommits_commitValid_32) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_32=0x%0h while the rhs_.io_diffCommits_commitValid_32=0x%0h",this.io_diffCommits_commitValid_32,rhs_.io_diffCommits_commitValid_32),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_33!=rhs_.io_diffCommits_commitValid_33) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_33=0x%0h while the rhs_.io_diffCommits_commitValid_33=0x%0h",this.io_diffCommits_commitValid_33,rhs_.io_diffCommits_commitValid_33),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_34!=rhs_.io_diffCommits_commitValid_34) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_34=0x%0h while the rhs_.io_diffCommits_commitValid_34=0x%0h",this.io_diffCommits_commitValid_34,rhs_.io_diffCommits_commitValid_34),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_35!=rhs_.io_diffCommits_commitValid_35) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_35=0x%0h while the rhs_.io_diffCommits_commitValid_35=0x%0h",this.io_diffCommits_commitValid_35,rhs_.io_diffCommits_commitValid_35),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_36!=rhs_.io_diffCommits_commitValid_36) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_36=0x%0h while the rhs_.io_diffCommits_commitValid_36=0x%0h",this.io_diffCommits_commitValid_36,rhs_.io_diffCommits_commitValid_36),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_37!=rhs_.io_diffCommits_commitValid_37) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_37=0x%0h while the rhs_.io_diffCommits_commitValid_37=0x%0h",this.io_diffCommits_commitValid_37,rhs_.io_diffCommits_commitValid_37),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_38!=rhs_.io_diffCommits_commitValid_38) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_38=0x%0h while the rhs_.io_diffCommits_commitValid_38=0x%0h",this.io_diffCommits_commitValid_38,rhs_.io_diffCommits_commitValid_38),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_39!=rhs_.io_diffCommits_commitValid_39) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_39=0x%0h while the rhs_.io_diffCommits_commitValid_39=0x%0h",this.io_diffCommits_commitValid_39,rhs_.io_diffCommits_commitValid_39),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_40!=rhs_.io_diffCommits_commitValid_40) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_40=0x%0h while the rhs_.io_diffCommits_commitValid_40=0x%0h",this.io_diffCommits_commitValid_40,rhs_.io_diffCommits_commitValid_40),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_41!=rhs_.io_diffCommits_commitValid_41) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_41=0x%0h while the rhs_.io_diffCommits_commitValid_41=0x%0h",this.io_diffCommits_commitValid_41,rhs_.io_diffCommits_commitValid_41),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_42!=rhs_.io_diffCommits_commitValid_42) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_42=0x%0h while the rhs_.io_diffCommits_commitValid_42=0x%0h",this.io_diffCommits_commitValid_42,rhs_.io_diffCommits_commitValid_42),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_43!=rhs_.io_diffCommits_commitValid_43) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_43=0x%0h while the rhs_.io_diffCommits_commitValid_43=0x%0h",this.io_diffCommits_commitValid_43,rhs_.io_diffCommits_commitValid_43),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_44!=rhs_.io_diffCommits_commitValid_44) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_44=0x%0h while the rhs_.io_diffCommits_commitValid_44=0x%0h",this.io_diffCommits_commitValid_44,rhs_.io_diffCommits_commitValid_44),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_45!=rhs_.io_diffCommits_commitValid_45) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_45=0x%0h while the rhs_.io_diffCommits_commitValid_45=0x%0h",this.io_diffCommits_commitValid_45,rhs_.io_diffCommits_commitValid_45),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_46!=rhs_.io_diffCommits_commitValid_46) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_46=0x%0h while the rhs_.io_diffCommits_commitValid_46=0x%0h",this.io_diffCommits_commitValid_46,rhs_.io_diffCommits_commitValid_46),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_47!=rhs_.io_diffCommits_commitValid_47) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_47=0x%0h while the rhs_.io_diffCommits_commitValid_47=0x%0h",this.io_diffCommits_commitValid_47,rhs_.io_diffCommits_commitValid_47),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_48!=rhs_.io_diffCommits_commitValid_48) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_48=0x%0h while the rhs_.io_diffCommits_commitValid_48=0x%0h",this.io_diffCommits_commitValid_48,rhs_.io_diffCommits_commitValid_48),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_49!=rhs_.io_diffCommits_commitValid_49) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_49=0x%0h while the rhs_.io_diffCommits_commitValid_49=0x%0h",this.io_diffCommits_commitValid_49,rhs_.io_diffCommits_commitValid_49),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_50!=rhs_.io_diffCommits_commitValid_50) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_50=0x%0h while the rhs_.io_diffCommits_commitValid_50=0x%0h",this.io_diffCommits_commitValid_50,rhs_.io_diffCommits_commitValid_50),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_51!=rhs_.io_diffCommits_commitValid_51) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_51=0x%0h while the rhs_.io_diffCommits_commitValid_51=0x%0h",this.io_diffCommits_commitValid_51,rhs_.io_diffCommits_commitValid_51),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_52!=rhs_.io_diffCommits_commitValid_52) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_52=0x%0h while the rhs_.io_diffCommits_commitValid_52=0x%0h",this.io_diffCommits_commitValid_52,rhs_.io_diffCommits_commitValid_52),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_53!=rhs_.io_diffCommits_commitValid_53) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_53=0x%0h while the rhs_.io_diffCommits_commitValid_53=0x%0h",this.io_diffCommits_commitValid_53,rhs_.io_diffCommits_commitValid_53),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_54!=rhs_.io_diffCommits_commitValid_54) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_54=0x%0h while the rhs_.io_diffCommits_commitValid_54=0x%0h",this.io_diffCommits_commitValid_54,rhs_.io_diffCommits_commitValid_54),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_55!=rhs_.io_diffCommits_commitValid_55) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_55=0x%0h while the rhs_.io_diffCommits_commitValid_55=0x%0h",this.io_diffCommits_commitValid_55,rhs_.io_diffCommits_commitValid_55),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_56!=rhs_.io_diffCommits_commitValid_56) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_56=0x%0h while the rhs_.io_diffCommits_commitValid_56=0x%0h",this.io_diffCommits_commitValid_56,rhs_.io_diffCommits_commitValid_56),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_57!=rhs_.io_diffCommits_commitValid_57) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_57=0x%0h while the rhs_.io_diffCommits_commitValid_57=0x%0h",this.io_diffCommits_commitValid_57,rhs_.io_diffCommits_commitValid_57),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_58!=rhs_.io_diffCommits_commitValid_58) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_58=0x%0h while the rhs_.io_diffCommits_commitValid_58=0x%0h",this.io_diffCommits_commitValid_58,rhs_.io_diffCommits_commitValid_58),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_59!=rhs_.io_diffCommits_commitValid_59) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_59=0x%0h while the rhs_.io_diffCommits_commitValid_59=0x%0h",this.io_diffCommits_commitValid_59,rhs_.io_diffCommits_commitValid_59),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_60!=rhs_.io_diffCommits_commitValid_60) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_60=0x%0h while the rhs_.io_diffCommits_commitValid_60=0x%0h",this.io_diffCommits_commitValid_60,rhs_.io_diffCommits_commitValid_60),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_61!=rhs_.io_diffCommits_commitValid_61) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_61=0x%0h while the rhs_.io_diffCommits_commitValid_61=0x%0h",this.io_diffCommits_commitValid_61,rhs_.io_diffCommits_commitValid_61),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_62!=rhs_.io_diffCommits_commitValid_62) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_62=0x%0h while the rhs_.io_diffCommits_commitValid_62=0x%0h",this.io_diffCommits_commitValid_62,rhs_.io_diffCommits_commitValid_62),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_63!=rhs_.io_diffCommits_commitValid_63) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_63=0x%0h while the rhs_.io_diffCommits_commitValid_63=0x%0h",this.io_diffCommits_commitValid_63,rhs_.io_diffCommits_commitValid_63),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_64!=rhs_.io_diffCommits_commitValid_64) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_64=0x%0h while the rhs_.io_diffCommits_commitValid_64=0x%0h",this.io_diffCommits_commitValid_64,rhs_.io_diffCommits_commitValid_64),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_65!=rhs_.io_diffCommits_commitValid_65) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_65=0x%0h while the rhs_.io_diffCommits_commitValid_65=0x%0h",this.io_diffCommits_commitValid_65,rhs_.io_diffCommits_commitValid_65),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_66!=rhs_.io_diffCommits_commitValid_66) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_66=0x%0h while the rhs_.io_diffCommits_commitValid_66=0x%0h",this.io_diffCommits_commitValid_66,rhs_.io_diffCommits_commitValid_66),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_67!=rhs_.io_diffCommits_commitValid_67) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_67=0x%0h while the rhs_.io_diffCommits_commitValid_67=0x%0h",this.io_diffCommits_commitValid_67,rhs_.io_diffCommits_commitValid_67),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_68!=rhs_.io_diffCommits_commitValid_68) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_68=0x%0h while the rhs_.io_diffCommits_commitValid_68=0x%0h",this.io_diffCommits_commitValid_68,rhs_.io_diffCommits_commitValid_68),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_69!=rhs_.io_diffCommits_commitValid_69) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_69=0x%0h while the rhs_.io_diffCommits_commitValid_69=0x%0h",this.io_diffCommits_commitValid_69,rhs_.io_diffCommits_commitValid_69),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_70!=rhs_.io_diffCommits_commitValid_70) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_70=0x%0h while the rhs_.io_diffCommits_commitValid_70=0x%0h",this.io_diffCommits_commitValid_70,rhs_.io_diffCommits_commitValid_70),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_71!=rhs_.io_diffCommits_commitValid_71) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_71=0x%0h while the rhs_.io_diffCommits_commitValid_71=0x%0h",this.io_diffCommits_commitValid_71,rhs_.io_diffCommits_commitValid_71),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_72!=rhs_.io_diffCommits_commitValid_72) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_72=0x%0h while the rhs_.io_diffCommits_commitValid_72=0x%0h",this.io_diffCommits_commitValid_72,rhs_.io_diffCommits_commitValid_72),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_73!=rhs_.io_diffCommits_commitValid_73) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_73=0x%0h while the rhs_.io_diffCommits_commitValid_73=0x%0h",this.io_diffCommits_commitValid_73,rhs_.io_diffCommits_commitValid_73),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_74!=rhs_.io_diffCommits_commitValid_74) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_74=0x%0h while the rhs_.io_diffCommits_commitValid_74=0x%0h",this.io_diffCommits_commitValid_74,rhs_.io_diffCommits_commitValid_74),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_75!=rhs_.io_diffCommits_commitValid_75) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_75=0x%0h while the rhs_.io_diffCommits_commitValid_75=0x%0h",this.io_diffCommits_commitValid_75,rhs_.io_diffCommits_commitValid_75),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_76!=rhs_.io_diffCommits_commitValid_76) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_76=0x%0h while the rhs_.io_diffCommits_commitValid_76=0x%0h",this.io_diffCommits_commitValid_76,rhs_.io_diffCommits_commitValid_76),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_77!=rhs_.io_diffCommits_commitValid_77) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_77=0x%0h while the rhs_.io_diffCommits_commitValid_77=0x%0h",this.io_diffCommits_commitValid_77,rhs_.io_diffCommits_commitValid_77),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_78!=rhs_.io_diffCommits_commitValid_78) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_78=0x%0h while the rhs_.io_diffCommits_commitValid_78=0x%0h",this.io_diffCommits_commitValid_78,rhs_.io_diffCommits_commitValid_78),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_79!=rhs_.io_diffCommits_commitValid_79) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_79=0x%0h while the rhs_.io_diffCommits_commitValid_79=0x%0h",this.io_diffCommits_commitValid_79,rhs_.io_diffCommits_commitValid_79),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_80!=rhs_.io_diffCommits_commitValid_80) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_80=0x%0h while the rhs_.io_diffCommits_commitValid_80=0x%0h",this.io_diffCommits_commitValid_80,rhs_.io_diffCommits_commitValid_80),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_81!=rhs_.io_diffCommits_commitValid_81) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_81=0x%0h while the rhs_.io_diffCommits_commitValid_81=0x%0h",this.io_diffCommits_commitValid_81,rhs_.io_diffCommits_commitValid_81),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_82!=rhs_.io_diffCommits_commitValid_82) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_82=0x%0h while the rhs_.io_diffCommits_commitValid_82=0x%0h",this.io_diffCommits_commitValid_82,rhs_.io_diffCommits_commitValid_82),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_83!=rhs_.io_diffCommits_commitValid_83) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_83=0x%0h while the rhs_.io_diffCommits_commitValid_83=0x%0h",this.io_diffCommits_commitValid_83,rhs_.io_diffCommits_commitValid_83),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_84!=rhs_.io_diffCommits_commitValid_84) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_84=0x%0h while the rhs_.io_diffCommits_commitValid_84=0x%0h",this.io_diffCommits_commitValid_84,rhs_.io_diffCommits_commitValid_84),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_85!=rhs_.io_diffCommits_commitValid_85) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_85=0x%0h while the rhs_.io_diffCommits_commitValid_85=0x%0h",this.io_diffCommits_commitValid_85,rhs_.io_diffCommits_commitValid_85),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_86!=rhs_.io_diffCommits_commitValid_86) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_86=0x%0h while the rhs_.io_diffCommits_commitValid_86=0x%0h",this.io_diffCommits_commitValid_86,rhs_.io_diffCommits_commitValid_86),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_87!=rhs_.io_diffCommits_commitValid_87) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_87=0x%0h while the rhs_.io_diffCommits_commitValid_87=0x%0h",this.io_diffCommits_commitValid_87,rhs_.io_diffCommits_commitValid_87),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_88!=rhs_.io_diffCommits_commitValid_88) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_88=0x%0h while the rhs_.io_diffCommits_commitValid_88=0x%0h",this.io_diffCommits_commitValid_88,rhs_.io_diffCommits_commitValid_88),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_89!=rhs_.io_diffCommits_commitValid_89) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_89=0x%0h while the rhs_.io_diffCommits_commitValid_89=0x%0h",this.io_diffCommits_commitValid_89,rhs_.io_diffCommits_commitValid_89),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_90!=rhs_.io_diffCommits_commitValid_90) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_90=0x%0h while the rhs_.io_diffCommits_commitValid_90=0x%0h",this.io_diffCommits_commitValid_90,rhs_.io_diffCommits_commitValid_90),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_91!=rhs_.io_diffCommits_commitValid_91) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_91=0x%0h while the rhs_.io_diffCommits_commitValid_91=0x%0h",this.io_diffCommits_commitValid_91,rhs_.io_diffCommits_commitValid_91),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_92!=rhs_.io_diffCommits_commitValid_92) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_92=0x%0h while the rhs_.io_diffCommits_commitValid_92=0x%0h",this.io_diffCommits_commitValid_92,rhs_.io_diffCommits_commitValid_92),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_93!=rhs_.io_diffCommits_commitValid_93) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_93=0x%0h while the rhs_.io_diffCommits_commitValid_93=0x%0h",this.io_diffCommits_commitValid_93,rhs_.io_diffCommits_commitValid_93),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_94!=rhs_.io_diffCommits_commitValid_94) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_94=0x%0h while the rhs_.io_diffCommits_commitValid_94=0x%0h",this.io_diffCommits_commitValid_94,rhs_.io_diffCommits_commitValid_94),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_95!=rhs_.io_diffCommits_commitValid_95) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_95=0x%0h while the rhs_.io_diffCommits_commitValid_95=0x%0h",this.io_diffCommits_commitValid_95,rhs_.io_diffCommits_commitValid_95),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_96!=rhs_.io_diffCommits_commitValid_96) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_96=0x%0h while the rhs_.io_diffCommits_commitValid_96=0x%0h",this.io_diffCommits_commitValid_96,rhs_.io_diffCommits_commitValid_96),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_97!=rhs_.io_diffCommits_commitValid_97) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_97=0x%0h while the rhs_.io_diffCommits_commitValid_97=0x%0h",this.io_diffCommits_commitValid_97,rhs_.io_diffCommits_commitValid_97),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_98!=rhs_.io_diffCommits_commitValid_98) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_98=0x%0h while the rhs_.io_diffCommits_commitValid_98=0x%0h",this.io_diffCommits_commitValid_98,rhs_.io_diffCommits_commitValid_98),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_99!=rhs_.io_diffCommits_commitValid_99) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_99=0x%0h while the rhs_.io_diffCommits_commitValid_99=0x%0h",this.io_diffCommits_commitValid_99,rhs_.io_diffCommits_commitValid_99),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_100!=rhs_.io_diffCommits_commitValid_100) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_100=0x%0h while the rhs_.io_diffCommits_commitValid_100=0x%0h",this.io_diffCommits_commitValid_100,rhs_.io_diffCommits_commitValid_100),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_101!=rhs_.io_diffCommits_commitValid_101) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_101=0x%0h while the rhs_.io_diffCommits_commitValid_101=0x%0h",this.io_diffCommits_commitValid_101,rhs_.io_diffCommits_commitValid_101),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_102!=rhs_.io_diffCommits_commitValid_102) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_102=0x%0h while the rhs_.io_diffCommits_commitValid_102=0x%0h",this.io_diffCommits_commitValid_102,rhs_.io_diffCommits_commitValid_102),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_103!=rhs_.io_diffCommits_commitValid_103) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_103=0x%0h while the rhs_.io_diffCommits_commitValid_103=0x%0h",this.io_diffCommits_commitValid_103,rhs_.io_diffCommits_commitValid_103),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_104!=rhs_.io_diffCommits_commitValid_104) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_104=0x%0h while the rhs_.io_diffCommits_commitValid_104=0x%0h",this.io_diffCommits_commitValid_104,rhs_.io_diffCommits_commitValid_104),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_105!=rhs_.io_diffCommits_commitValid_105) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_105=0x%0h while the rhs_.io_diffCommits_commitValid_105=0x%0h",this.io_diffCommits_commitValid_105,rhs_.io_diffCommits_commitValid_105),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_106!=rhs_.io_diffCommits_commitValid_106) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_106=0x%0h while the rhs_.io_diffCommits_commitValid_106=0x%0h",this.io_diffCommits_commitValid_106,rhs_.io_diffCommits_commitValid_106),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_107!=rhs_.io_diffCommits_commitValid_107) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_107=0x%0h while the rhs_.io_diffCommits_commitValid_107=0x%0h",this.io_diffCommits_commitValid_107,rhs_.io_diffCommits_commitValid_107),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_108!=rhs_.io_diffCommits_commitValid_108) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_108=0x%0h while the rhs_.io_diffCommits_commitValid_108=0x%0h",this.io_diffCommits_commitValid_108,rhs_.io_diffCommits_commitValid_108),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_109!=rhs_.io_diffCommits_commitValid_109) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_109=0x%0h while the rhs_.io_diffCommits_commitValid_109=0x%0h",this.io_diffCommits_commitValid_109,rhs_.io_diffCommits_commitValid_109),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_110!=rhs_.io_diffCommits_commitValid_110) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_110=0x%0h while the rhs_.io_diffCommits_commitValid_110=0x%0h",this.io_diffCommits_commitValid_110,rhs_.io_diffCommits_commitValid_110),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_111!=rhs_.io_diffCommits_commitValid_111) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_111=0x%0h while the rhs_.io_diffCommits_commitValid_111=0x%0h",this.io_diffCommits_commitValid_111,rhs_.io_diffCommits_commitValid_111),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_112!=rhs_.io_diffCommits_commitValid_112) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_112=0x%0h while the rhs_.io_diffCommits_commitValid_112=0x%0h",this.io_diffCommits_commitValid_112,rhs_.io_diffCommits_commitValid_112),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_113!=rhs_.io_diffCommits_commitValid_113) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_113=0x%0h while the rhs_.io_diffCommits_commitValid_113=0x%0h",this.io_diffCommits_commitValid_113,rhs_.io_diffCommits_commitValid_113),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_114!=rhs_.io_diffCommits_commitValid_114) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_114=0x%0h while the rhs_.io_diffCommits_commitValid_114=0x%0h",this.io_diffCommits_commitValid_114,rhs_.io_diffCommits_commitValid_114),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_115!=rhs_.io_diffCommits_commitValid_115) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_115=0x%0h while the rhs_.io_diffCommits_commitValid_115=0x%0h",this.io_diffCommits_commitValid_115,rhs_.io_diffCommits_commitValid_115),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_116!=rhs_.io_diffCommits_commitValid_116) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_116=0x%0h while the rhs_.io_diffCommits_commitValid_116=0x%0h",this.io_diffCommits_commitValid_116,rhs_.io_diffCommits_commitValid_116),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_117!=rhs_.io_diffCommits_commitValid_117) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_117=0x%0h while the rhs_.io_diffCommits_commitValid_117=0x%0h",this.io_diffCommits_commitValid_117,rhs_.io_diffCommits_commitValid_117),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_118!=rhs_.io_diffCommits_commitValid_118) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_118=0x%0h while the rhs_.io_diffCommits_commitValid_118=0x%0h",this.io_diffCommits_commitValid_118,rhs_.io_diffCommits_commitValid_118),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_119!=rhs_.io_diffCommits_commitValid_119) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_119=0x%0h while the rhs_.io_diffCommits_commitValid_119=0x%0h",this.io_diffCommits_commitValid_119,rhs_.io_diffCommits_commitValid_119),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_120!=rhs_.io_diffCommits_commitValid_120) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_120=0x%0h while the rhs_.io_diffCommits_commitValid_120=0x%0h",this.io_diffCommits_commitValid_120,rhs_.io_diffCommits_commitValid_120),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_121!=rhs_.io_diffCommits_commitValid_121) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_121=0x%0h while the rhs_.io_diffCommits_commitValid_121=0x%0h",this.io_diffCommits_commitValid_121,rhs_.io_diffCommits_commitValid_121),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_122!=rhs_.io_diffCommits_commitValid_122) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_122=0x%0h while the rhs_.io_diffCommits_commitValid_122=0x%0h",this.io_diffCommits_commitValid_122,rhs_.io_diffCommits_commitValid_122),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_123!=rhs_.io_diffCommits_commitValid_123) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_123=0x%0h while the rhs_.io_diffCommits_commitValid_123=0x%0h",this.io_diffCommits_commitValid_123,rhs_.io_diffCommits_commitValid_123),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_124!=rhs_.io_diffCommits_commitValid_124) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_124=0x%0h while the rhs_.io_diffCommits_commitValid_124=0x%0h",this.io_diffCommits_commitValid_124,rhs_.io_diffCommits_commitValid_124),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_125!=rhs_.io_diffCommits_commitValid_125) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_125=0x%0h while the rhs_.io_diffCommits_commitValid_125=0x%0h",this.io_diffCommits_commitValid_125,rhs_.io_diffCommits_commitValid_125),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_126!=rhs_.io_diffCommits_commitValid_126) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_126=0x%0h while the rhs_.io_diffCommits_commitValid_126=0x%0h",this.io_diffCommits_commitValid_126,rhs_.io_diffCommits_commitValid_126),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_127!=rhs_.io_diffCommits_commitValid_127) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_127=0x%0h while the rhs_.io_diffCommits_commitValid_127=0x%0h",this.io_diffCommits_commitValid_127,rhs_.io_diffCommits_commitValid_127),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_128!=rhs_.io_diffCommits_commitValid_128) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_128=0x%0h while the rhs_.io_diffCommits_commitValid_128=0x%0h",this.io_diffCommits_commitValid_128,rhs_.io_diffCommits_commitValid_128),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_129!=rhs_.io_diffCommits_commitValid_129) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_129=0x%0h while the rhs_.io_diffCommits_commitValid_129=0x%0h",this.io_diffCommits_commitValid_129,rhs_.io_diffCommits_commitValid_129),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_130!=rhs_.io_diffCommits_commitValid_130) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_130=0x%0h while the rhs_.io_diffCommits_commitValid_130=0x%0h",this.io_diffCommits_commitValid_130,rhs_.io_diffCommits_commitValid_130),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_131!=rhs_.io_diffCommits_commitValid_131) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_131=0x%0h while the rhs_.io_diffCommits_commitValid_131=0x%0h",this.io_diffCommits_commitValid_131,rhs_.io_diffCommits_commitValid_131),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_132!=rhs_.io_diffCommits_commitValid_132) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_132=0x%0h while the rhs_.io_diffCommits_commitValid_132=0x%0h",this.io_diffCommits_commitValid_132,rhs_.io_diffCommits_commitValid_132),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_133!=rhs_.io_diffCommits_commitValid_133) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_133=0x%0h while the rhs_.io_diffCommits_commitValid_133=0x%0h",this.io_diffCommits_commitValid_133,rhs_.io_diffCommits_commitValid_133),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_134!=rhs_.io_diffCommits_commitValid_134) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_134=0x%0h while the rhs_.io_diffCommits_commitValid_134=0x%0h",this.io_diffCommits_commitValid_134,rhs_.io_diffCommits_commitValid_134),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_135!=rhs_.io_diffCommits_commitValid_135) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_135=0x%0h while the rhs_.io_diffCommits_commitValid_135=0x%0h",this.io_diffCommits_commitValid_135,rhs_.io_diffCommits_commitValid_135),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_136!=rhs_.io_diffCommits_commitValid_136) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_136=0x%0h while the rhs_.io_diffCommits_commitValid_136=0x%0h",this.io_diffCommits_commitValid_136,rhs_.io_diffCommits_commitValid_136),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_137!=rhs_.io_diffCommits_commitValid_137) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_137=0x%0h while the rhs_.io_diffCommits_commitValid_137=0x%0h",this.io_diffCommits_commitValid_137,rhs_.io_diffCommits_commitValid_137),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_138!=rhs_.io_diffCommits_commitValid_138) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_138=0x%0h while the rhs_.io_diffCommits_commitValid_138=0x%0h",this.io_diffCommits_commitValid_138,rhs_.io_diffCommits_commitValid_138),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_139!=rhs_.io_diffCommits_commitValid_139) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_139=0x%0h while the rhs_.io_diffCommits_commitValid_139=0x%0h",this.io_diffCommits_commitValid_139,rhs_.io_diffCommits_commitValid_139),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_140!=rhs_.io_diffCommits_commitValid_140) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_140=0x%0h while the rhs_.io_diffCommits_commitValid_140=0x%0h",this.io_diffCommits_commitValid_140,rhs_.io_diffCommits_commitValid_140),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_141!=rhs_.io_diffCommits_commitValid_141) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_141=0x%0h while the rhs_.io_diffCommits_commitValid_141=0x%0h",this.io_diffCommits_commitValid_141,rhs_.io_diffCommits_commitValid_141),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_142!=rhs_.io_diffCommits_commitValid_142) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_142=0x%0h while the rhs_.io_diffCommits_commitValid_142=0x%0h",this.io_diffCommits_commitValid_142,rhs_.io_diffCommits_commitValid_142),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_143!=rhs_.io_diffCommits_commitValid_143) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_143=0x%0h while the rhs_.io_diffCommits_commitValid_143=0x%0h",this.io_diffCommits_commitValid_143,rhs_.io_diffCommits_commitValid_143),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_144!=rhs_.io_diffCommits_commitValid_144) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_144=0x%0h while the rhs_.io_diffCommits_commitValid_144=0x%0h",this.io_diffCommits_commitValid_144,rhs_.io_diffCommits_commitValid_144),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_145!=rhs_.io_diffCommits_commitValid_145) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_145=0x%0h while the rhs_.io_diffCommits_commitValid_145=0x%0h",this.io_diffCommits_commitValid_145,rhs_.io_diffCommits_commitValid_145),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_146!=rhs_.io_diffCommits_commitValid_146) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_146=0x%0h while the rhs_.io_diffCommits_commitValid_146=0x%0h",this.io_diffCommits_commitValid_146,rhs_.io_diffCommits_commitValid_146),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_147!=rhs_.io_diffCommits_commitValid_147) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_147=0x%0h while the rhs_.io_diffCommits_commitValid_147=0x%0h",this.io_diffCommits_commitValid_147,rhs_.io_diffCommits_commitValid_147),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_148!=rhs_.io_diffCommits_commitValid_148) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_148=0x%0h while the rhs_.io_diffCommits_commitValid_148=0x%0h",this.io_diffCommits_commitValid_148,rhs_.io_diffCommits_commitValid_148),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_149!=rhs_.io_diffCommits_commitValid_149) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_149=0x%0h while the rhs_.io_diffCommits_commitValid_149=0x%0h",this.io_diffCommits_commitValid_149,rhs_.io_diffCommits_commitValid_149),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_150!=rhs_.io_diffCommits_commitValid_150) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_150=0x%0h while the rhs_.io_diffCommits_commitValid_150=0x%0h",this.io_diffCommits_commitValid_150,rhs_.io_diffCommits_commitValid_150),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_151!=rhs_.io_diffCommits_commitValid_151) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_151=0x%0h while the rhs_.io_diffCommits_commitValid_151=0x%0h",this.io_diffCommits_commitValid_151,rhs_.io_diffCommits_commitValid_151),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_152!=rhs_.io_diffCommits_commitValid_152) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_152=0x%0h while the rhs_.io_diffCommits_commitValid_152=0x%0h",this.io_diffCommits_commitValid_152,rhs_.io_diffCommits_commitValid_152),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_153!=rhs_.io_diffCommits_commitValid_153) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_153=0x%0h while the rhs_.io_diffCommits_commitValid_153=0x%0h",this.io_diffCommits_commitValid_153,rhs_.io_diffCommits_commitValid_153),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_154!=rhs_.io_diffCommits_commitValid_154) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_154=0x%0h while the rhs_.io_diffCommits_commitValid_154=0x%0h",this.io_diffCommits_commitValid_154,rhs_.io_diffCommits_commitValid_154),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_155!=rhs_.io_diffCommits_commitValid_155) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_155=0x%0h while the rhs_.io_diffCommits_commitValid_155=0x%0h",this.io_diffCommits_commitValid_155,rhs_.io_diffCommits_commitValid_155),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_156!=rhs_.io_diffCommits_commitValid_156) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_156=0x%0h while the rhs_.io_diffCommits_commitValid_156=0x%0h",this.io_diffCommits_commitValid_156,rhs_.io_diffCommits_commitValid_156),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_157!=rhs_.io_diffCommits_commitValid_157) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_157=0x%0h while the rhs_.io_diffCommits_commitValid_157=0x%0h",this.io_diffCommits_commitValid_157,rhs_.io_diffCommits_commitValid_157),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_158!=rhs_.io_diffCommits_commitValid_158) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_158=0x%0h while the rhs_.io_diffCommits_commitValid_158=0x%0h",this.io_diffCommits_commitValid_158,rhs_.io_diffCommits_commitValid_158),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_159!=rhs_.io_diffCommits_commitValid_159) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_159=0x%0h while the rhs_.io_diffCommits_commitValid_159=0x%0h",this.io_diffCommits_commitValid_159,rhs_.io_diffCommits_commitValid_159),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_160!=rhs_.io_diffCommits_commitValid_160) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_160=0x%0h while the rhs_.io_diffCommits_commitValid_160=0x%0h",this.io_diffCommits_commitValid_160,rhs_.io_diffCommits_commitValid_160),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_161!=rhs_.io_diffCommits_commitValid_161) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_161=0x%0h while the rhs_.io_diffCommits_commitValid_161=0x%0h",this.io_diffCommits_commitValid_161,rhs_.io_diffCommits_commitValid_161),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_162!=rhs_.io_diffCommits_commitValid_162) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_162=0x%0h while the rhs_.io_diffCommits_commitValid_162=0x%0h",this.io_diffCommits_commitValid_162,rhs_.io_diffCommits_commitValid_162),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_163!=rhs_.io_diffCommits_commitValid_163) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_163=0x%0h while the rhs_.io_diffCommits_commitValid_163=0x%0h",this.io_diffCommits_commitValid_163,rhs_.io_diffCommits_commitValid_163),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_164!=rhs_.io_diffCommits_commitValid_164) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_164=0x%0h while the rhs_.io_diffCommits_commitValid_164=0x%0h",this.io_diffCommits_commitValid_164,rhs_.io_diffCommits_commitValid_164),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_165!=rhs_.io_diffCommits_commitValid_165) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_165=0x%0h while the rhs_.io_diffCommits_commitValid_165=0x%0h",this.io_diffCommits_commitValid_165,rhs_.io_diffCommits_commitValid_165),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_166!=rhs_.io_diffCommits_commitValid_166) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_166=0x%0h while the rhs_.io_diffCommits_commitValid_166=0x%0h",this.io_diffCommits_commitValid_166,rhs_.io_diffCommits_commitValid_166),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_167!=rhs_.io_diffCommits_commitValid_167) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_167=0x%0h while the rhs_.io_diffCommits_commitValid_167=0x%0h",this.io_diffCommits_commitValid_167,rhs_.io_diffCommits_commitValid_167),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_168!=rhs_.io_diffCommits_commitValid_168) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_168=0x%0h while the rhs_.io_diffCommits_commitValid_168=0x%0h",this.io_diffCommits_commitValid_168,rhs_.io_diffCommits_commitValid_168),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_169!=rhs_.io_diffCommits_commitValid_169) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_169=0x%0h while the rhs_.io_diffCommits_commitValid_169=0x%0h",this.io_diffCommits_commitValid_169,rhs_.io_diffCommits_commitValid_169),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_170!=rhs_.io_diffCommits_commitValid_170) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_170=0x%0h while the rhs_.io_diffCommits_commitValid_170=0x%0h",this.io_diffCommits_commitValid_170,rhs_.io_diffCommits_commitValid_170),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_171!=rhs_.io_diffCommits_commitValid_171) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_171=0x%0h while the rhs_.io_diffCommits_commitValid_171=0x%0h",this.io_diffCommits_commitValid_171,rhs_.io_diffCommits_commitValid_171),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_172!=rhs_.io_diffCommits_commitValid_172) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_172=0x%0h while the rhs_.io_diffCommits_commitValid_172=0x%0h",this.io_diffCommits_commitValid_172,rhs_.io_diffCommits_commitValid_172),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_173!=rhs_.io_diffCommits_commitValid_173) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_173=0x%0h while the rhs_.io_diffCommits_commitValid_173=0x%0h",this.io_diffCommits_commitValid_173,rhs_.io_diffCommits_commitValid_173),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_174!=rhs_.io_diffCommits_commitValid_174) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_174=0x%0h while the rhs_.io_diffCommits_commitValid_174=0x%0h",this.io_diffCommits_commitValid_174,rhs_.io_diffCommits_commitValid_174),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_175!=rhs_.io_diffCommits_commitValid_175) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_175=0x%0h while the rhs_.io_diffCommits_commitValid_175=0x%0h",this.io_diffCommits_commitValid_175,rhs_.io_diffCommits_commitValid_175),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_176!=rhs_.io_diffCommits_commitValid_176) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_176=0x%0h while the rhs_.io_diffCommits_commitValid_176=0x%0h",this.io_diffCommits_commitValid_176,rhs_.io_diffCommits_commitValid_176),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_177!=rhs_.io_diffCommits_commitValid_177) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_177=0x%0h while the rhs_.io_diffCommits_commitValid_177=0x%0h",this.io_diffCommits_commitValid_177,rhs_.io_diffCommits_commitValid_177),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_178!=rhs_.io_diffCommits_commitValid_178) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_178=0x%0h while the rhs_.io_diffCommits_commitValid_178=0x%0h",this.io_diffCommits_commitValid_178,rhs_.io_diffCommits_commitValid_178),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_179!=rhs_.io_diffCommits_commitValid_179) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_179=0x%0h while the rhs_.io_diffCommits_commitValid_179=0x%0h",this.io_diffCommits_commitValid_179,rhs_.io_diffCommits_commitValid_179),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_180!=rhs_.io_diffCommits_commitValid_180) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_180=0x%0h while the rhs_.io_diffCommits_commitValid_180=0x%0h",this.io_diffCommits_commitValid_180,rhs_.io_diffCommits_commitValid_180),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_181!=rhs_.io_diffCommits_commitValid_181) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_181=0x%0h while the rhs_.io_diffCommits_commitValid_181=0x%0h",this.io_diffCommits_commitValid_181,rhs_.io_diffCommits_commitValid_181),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_182!=rhs_.io_diffCommits_commitValid_182) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_182=0x%0h while the rhs_.io_diffCommits_commitValid_182=0x%0h",this.io_diffCommits_commitValid_182,rhs_.io_diffCommits_commitValid_182),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_183!=rhs_.io_diffCommits_commitValid_183) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_183=0x%0h while the rhs_.io_diffCommits_commitValid_183=0x%0h",this.io_diffCommits_commitValid_183,rhs_.io_diffCommits_commitValid_183),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_184!=rhs_.io_diffCommits_commitValid_184) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_184=0x%0h while the rhs_.io_diffCommits_commitValid_184=0x%0h",this.io_diffCommits_commitValid_184,rhs_.io_diffCommits_commitValid_184),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_185!=rhs_.io_diffCommits_commitValid_185) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_185=0x%0h while the rhs_.io_diffCommits_commitValid_185=0x%0h",this.io_diffCommits_commitValid_185,rhs_.io_diffCommits_commitValid_185),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_186!=rhs_.io_diffCommits_commitValid_186) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_186=0x%0h while the rhs_.io_diffCommits_commitValid_186=0x%0h",this.io_diffCommits_commitValid_186,rhs_.io_diffCommits_commitValid_186),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_187!=rhs_.io_diffCommits_commitValid_187) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_187=0x%0h while the rhs_.io_diffCommits_commitValid_187=0x%0h",this.io_diffCommits_commitValid_187,rhs_.io_diffCommits_commitValid_187),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_188!=rhs_.io_diffCommits_commitValid_188) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_188=0x%0h while the rhs_.io_diffCommits_commitValid_188=0x%0h",this.io_diffCommits_commitValid_188,rhs_.io_diffCommits_commitValid_188),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_189!=rhs_.io_diffCommits_commitValid_189) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_189=0x%0h while the rhs_.io_diffCommits_commitValid_189=0x%0h",this.io_diffCommits_commitValid_189,rhs_.io_diffCommits_commitValid_189),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_190!=rhs_.io_diffCommits_commitValid_190) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_190=0x%0h while the rhs_.io_diffCommits_commitValid_190=0x%0h",this.io_diffCommits_commitValid_190,rhs_.io_diffCommits_commitValid_190),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_191!=rhs_.io_diffCommits_commitValid_191) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_191=0x%0h while the rhs_.io_diffCommits_commitValid_191=0x%0h",this.io_diffCommits_commitValid_191,rhs_.io_diffCommits_commitValid_191),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_192!=rhs_.io_diffCommits_commitValid_192) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_192=0x%0h while the rhs_.io_diffCommits_commitValid_192=0x%0h",this.io_diffCommits_commitValid_192,rhs_.io_diffCommits_commitValid_192),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_193!=rhs_.io_diffCommits_commitValid_193) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_193=0x%0h while the rhs_.io_diffCommits_commitValid_193=0x%0h",this.io_diffCommits_commitValid_193,rhs_.io_diffCommits_commitValid_193),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_194!=rhs_.io_diffCommits_commitValid_194) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_194=0x%0h while the rhs_.io_diffCommits_commitValid_194=0x%0h",this.io_diffCommits_commitValid_194,rhs_.io_diffCommits_commitValid_194),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_195!=rhs_.io_diffCommits_commitValid_195) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_195=0x%0h while the rhs_.io_diffCommits_commitValid_195=0x%0h",this.io_diffCommits_commitValid_195,rhs_.io_diffCommits_commitValid_195),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_196!=rhs_.io_diffCommits_commitValid_196) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_196=0x%0h while the rhs_.io_diffCommits_commitValid_196=0x%0h",this.io_diffCommits_commitValid_196,rhs_.io_diffCommits_commitValid_196),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_197!=rhs_.io_diffCommits_commitValid_197) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_197=0x%0h while the rhs_.io_diffCommits_commitValid_197=0x%0h",this.io_diffCommits_commitValid_197,rhs_.io_diffCommits_commitValid_197),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_198!=rhs_.io_diffCommits_commitValid_198) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_198=0x%0h while the rhs_.io_diffCommits_commitValid_198=0x%0h",this.io_diffCommits_commitValid_198,rhs_.io_diffCommits_commitValid_198),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_199!=rhs_.io_diffCommits_commitValid_199) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_199=0x%0h while the rhs_.io_diffCommits_commitValid_199=0x%0h",this.io_diffCommits_commitValid_199,rhs_.io_diffCommits_commitValid_199),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_200!=rhs_.io_diffCommits_commitValid_200) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_200=0x%0h while the rhs_.io_diffCommits_commitValid_200=0x%0h",this.io_diffCommits_commitValid_200,rhs_.io_diffCommits_commitValid_200),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_201!=rhs_.io_diffCommits_commitValid_201) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_201=0x%0h while the rhs_.io_diffCommits_commitValid_201=0x%0h",this.io_diffCommits_commitValid_201,rhs_.io_diffCommits_commitValid_201),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_202!=rhs_.io_diffCommits_commitValid_202) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_202=0x%0h while the rhs_.io_diffCommits_commitValid_202=0x%0h",this.io_diffCommits_commitValid_202,rhs_.io_diffCommits_commitValid_202),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_203!=rhs_.io_diffCommits_commitValid_203) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_203=0x%0h while the rhs_.io_diffCommits_commitValid_203=0x%0h",this.io_diffCommits_commitValid_203,rhs_.io_diffCommits_commitValid_203),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_204!=rhs_.io_diffCommits_commitValid_204) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_204=0x%0h while the rhs_.io_diffCommits_commitValid_204=0x%0h",this.io_diffCommits_commitValid_204,rhs_.io_diffCommits_commitValid_204),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_205!=rhs_.io_diffCommits_commitValid_205) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_205=0x%0h while the rhs_.io_diffCommits_commitValid_205=0x%0h",this.io_diffCommits_commitValid_205,rhs_.io_diffCommits_commitValid_205),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_206!=rhs_.io_diffCommits_commitValid_206) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_206=0x%0h while the rhs_.io_diffCommits_commitValid_206=0x%0h",this.io_diffCommits_commitValid_206,rhs_.io_diffCommits_commitValid_206),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_207!=rhs_.io_diffCommits_commitValid_207) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_207=0x%0h while the rhs_.io_diffCommits_commitValid_207=0x%0h",this.io_diffCommits_commitValid_207,rhs_.io_diffCommits_commitValid_207),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_208!=rhs_.io_diffCommits_commitValid_208) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_208=0x%0h while the rhs_.io_diffCommits_commitValid_208=0x%0h",this.io_diffCommits_commitValid_208,rhs_.io_diffCommits_commitValid_208),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_209!=rhs_.io_diffCommits_commitValid_209) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_209=0x%0h while the rhs_.io_diffCommits_commitValid_209=0x%0h",this.io_diffCommits_commitValid_209,rhs_.io_diffCommits_commitValid_209),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_210!=rhs_.io_diffCommits_commitValid_210) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_210=0x%0h while the rhs_.io_diffCommits_commitValid_210=0x%0h",this.io_diffCommits_commitValid_210,rhs_.io_diffCommits_commitValid_210),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_211!=rhs_.io_diffCommits_commitValid_211) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_211=0x%0h while the rhs_.io_diffCommits_commitValid_211=0x%0h",this.io_diffCommits_commitValid_211,rhs_.io_diffCommits_commitValid_211),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_212!=rhs_.io_diffCommits_commitValid_212) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_212=0x%0h while the rhs_.io_diffCommits_commitValid_212=0x%0h",this.io_diffCommits_commitValid_212,rhs_.io_diffCommits_commitValid_212),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_213!=rhs_.io_diffCommits_commitValid_213) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_213=0x%0h while the rhs_.io_diffCommits_commitValid_213=0x%0h",this.io_diffCommits_commitValid_213,rhs_.io_diffCommits_commitValid_213),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_214!=rhs_.io_diffCommits_commitValid_214) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_214=0x%0h while the rhs_.io_diffCommits_commitValid_214=0x%0h",this.io_diffCommits_commitValid_214,rhs_.io_diffCommits_commitValid_214),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_215!=rhs_.io_diffCommits_commitValid_215) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_215=0x%0h while the rhs_.io_diffCommits_commitValid_215=0x%0h",this.io_diffCommits_commitValid_215,rhs_.io_diffCommits_commitValid_215),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_216!=rhs_.io_diffCommits_commitValid_216) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_216=0x%0h while the rhs_.io_diffCommits_commitValid_216=0x%0h",this.io_diffCommits_commitValid_216,rhs_.io_diffCommits_commitValid_216),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_217!=rhs_.io_diffCommits_commitValid_217) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_217=0x%0h while the rhs_.io_diffCommits_commitValid_217=0x%0h",this.io_diffCommits_commitValid_217,rhs_.io_diffCommits_commitValid_217),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_218!=rhs_.io_diffCommits_commitValid_218) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_218=0x%0h while the rhs_.io_diffCommits_commitValid_218=0x%0h",this.io_diffCommits_commitValid_218,rhs_.io_diffCommits_commitValid_218),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_219!=rhs_.io_diffCommits_commitValid_219) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_219=0x%0h while the rhs_.io_diffCommits_commitValid_219=0x%0h",this.io_diffCommits_commitValid_219,rhs_.io_diffCommits_commitValid_219),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_220!=rhs_.io_diffCommits_commitValid_220) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_220=0x%0h while the rhs_.io_diffCommits_commitValid_220=0x%0h",this.io_diffCommits_commitValid_220,rhs_.io_diffCommits_commitValid_220),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_221!=rhs_.io_diffCommits_commitValid_221) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_221=0x%0h while the rhs_.io_diffCommits_commitValid_221=0x%0h",this.io_diffCommits_commitValid_221,rhs_.io_diffCommits_commitValid_221),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_222!=rhs_.io_diffCommits_commitValid_222) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_222=0x%0h while the rhs_.io_diffCommits_commitValid_222=0x%0h",this.io_diffCommits_commitValid_222,rhs_.io_diffCommits_commitValid_222),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_223!=rhs_.io_diffCommits_commitValid_223) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_223=0x%0h while the rhs_.io_diffCommits_commitValid_223=0x%0h",this.io_diffCommits_commitValid_223,rhs_.io_diffCommits_commitValid_223),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_224!=rhs_.io_diffCommits_commitValid_224) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_224=0x%0h while the rhs_.io_diffCommits_commitValid_224=0x%0h",this.io_diffCommits_commitValid_224,rhs_.io_diffCommits_commitValid_224),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_225!=rhs_.io_diffCommits_commitValid_225) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_225=0x%0h while the rhs_.io_diffCommits_commitValid_225=0x%0h",this.io_diffCommits_commitValid_225,rhs_.io_diffCommits_commitValid_225),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_226!=rhs_.io_diffCommits_commitValid_226) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_226=0x%0h while the rhs_.io_diffCommits_commitValid_226=0x%0h",this.io_diffCommits_commitValid_226,rhs_.io_diffCommits_commitValid_226),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_227!=rhs_.io_diffCommits_commitValid_227) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_227=0x%0h while the rhs_.io_diffCommits_commitValid_227=0x%0h",this.io_diffCommits_commitValid_227,rhs_.io_diffCommits_commitValid_227),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_228!=rhs_.io_diffCommits_commitValid_228) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_228=0x%0h while the rhs_.io_diffCommits_commitValid_228=0x%0h",this.io_diffCommits_commitValid_228,rhs_.io_diffCommits_commitValid_228),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_229!=rhs_.io_diffCommits_commitValid_229) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_229=0x%0h while the rhs_.io_diffCommits_commitValid_229=0x%0h",this.io_diffCommits_commitValid_229,rhs_.io_diffCommits_commitValid_229),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_230!=rhs_.io_diffCommits_commitValid_230) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_230=0x%0h while the rhs_.io_diffCommits_commitValid_230=0x%0h",this.io_diffCommits_commitValid_230,rhs_.io_diffCommits_commitValid_230),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_231!=rhs_.io_diffCommits_commitValid_231) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_231=0x%0h while the rhs_.io_diffCommits_commitValid_231=0x%0h",this.io_diffCommits_commitValid_231,rhs_.io_diffCommits_commitValid_231),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_232!=rhs_.io_diffCommits_commitValid_232) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_232=0x%0h while the rhs_.io_diffCommits_commitValid_232=0x%0h",this.io_diffCommits_commitValid_232,rhs_.io_diffCommits_commitValid_232),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_233!=rhs_.io_diffCommits_commitValid_233) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_233=0x%0h while the rhs_.io_diffCommits_commitValid_233=0x%0h",this.io_diffCommits_commitValid_233,rhs_.io_diffCommits_commitValid_233),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_234!=rhs_.io_diffCommits_commitValid_234) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_234=0x%0h while the rhs_.io_diffCommits_commitValid_234=0x%0h",this.io_diffCommits_commitValid_234,rhs_.io_diffCommits_commitValid_234),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_235!=rhs_.io_diffCommits_commitValid_235) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_235=0x%0h while the rhs_.io_diffCommits_commitValid_235=0x%0h",this.io_diffCommits_commitValid_235,rhs_.io_diffCommits_commitValid_235),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_236!=rhs_.io_diffCommits_commitValid_236) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_236=0x%0h while the rhs_.io_diffCommits_commitValid_236=0x%0h",this.io_diffCommits_commitValid_236,rhs_.io_diffCommits_commitValid_236),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_237!=rhs_.io_diffCommits_commitValid_237) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_237=0x%0h while the rhs_.io_diffCommits_commitValid_237=0x%0h",this.io_diffCommits_commitValid_237,rhs_.io_diffCommits_commitValid_237),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_238!=rhs_.io_diffCommits_commitValid_238) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_238=0x%0h while the rhs_.io_diffCommits_commitValid_238=0x%0h",this.io_diffCommits_commitValid_238,rhs_.io_diffCommits_commitValid_238),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_239!=rhs_.io_diffCommits_commitValid_239) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_239=0x%0h while the rhs_.io_diffCommits_commitValid_239=0x%0h",this.io_diffCommits_commitValid_239,rhs_.io_diffCommits_commitValid_239),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_240!=rhs_.io_diffCommits_commitValid_240) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_240=0x%0h while the rhs_.io_diffCommits_commitValid_240=0x%0h",this.io_diffCommits_commitValid_240,rhs_.io_diffCommits_commitValid_240),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_241!=rhs_.io_diffCommits_commitValid_241) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_241=0x%0h while the rhs_.io_diffCommits_commitValid_241=0x%0h",this.io_diffCommits_commitValid_241,rhs_.io_diffCommits_commitValid_241),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_242!=rhs_.io_diffCommits_commitValid_242) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_242=0x%0h while the rhs_.io_diffCommits_commitValid_242=0x%0h",this.io_diffCommits_commitValid_242,rhs_.io_diffCommits_commitValid_242),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_243!=rhs_.io_diffCommits_commitValid_243) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_243=0x%0h while the rhs_.io_diffCommits_commitValid_243=0x%0h",this.io_diffCommits_commitValid_243,rhs_.io_diffCommits_commitValid_243),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_244!=rhs_.io_diffCommits_commitValid_244) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_244=0x%0h while the rhs_.io_diffCommits_commitValid_244=0x%0h",this.io_diffCommits_commitValid_244,rhs_.io_diffCommits_commitValid_244),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_245!=rhs_.io_diffCommits_commitValid_245) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_245=0x%0h while the rhs_.io_diffCommits_commitValid_245=0x%0h",this.io_diffCommits_commitValid_245,rhs_.io_diffCommits_commitValid_245),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_246!=rhs_.io_diffCommits_commitValid_246) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_246=0x%0h while the rhs_.io_diffCommits_commitValid_246=0x%0h",this.io_diffCommits_commitValid_246,rhs_.io_diffCommits_commitValid_246),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_247!=rhs_.io_diffCommits_commitValid_247) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_247=0x%0h while the rhs_.io_diffCommits_commitValid_247=0x%0h",this.io_diffCommits_commitValid_247,rhs_.io_diffCommits_commitValid_247),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_248!=rhs_.io_diffCommits_commitValid_248) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_248=0x%0h while the rhs_.io_diffCommits_commitValid_248=0x%0h",this.io_diffCommits_commitValid_248,rhs_.io_diffCommits_commitValid_248),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_249!=rhs_.io_diffCommits_commitValid_249) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_249=0x%0h while the rhs_.io_diffCommits_commitValid_249=0x%0h",this.io_diffCommits_commitValid_249,rhs_.io_diffCommits_commitValid_249),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_250!=rhs_.io_diffCommits_commitValid_250) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_250=0x%0h while the rhs_.io_diffCommits_commitValid_250=0x%0h",this.io_diffCommits_commitValid_250,rhs_.io_diffCommits_commitValid_250),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_251!=rhs_.io_diffCommits_commitValid_251) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_251=0x%0h while the rhs_.io_diffCommits_commitValid_251=0x%0h",this.io_diffCommits_commitValid_251,rhs_.io_diffCommits_commitValid_251),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_252!=rhs_.io_diffCommits_commitValid_252) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_252=0x%0h while the rhs_.io_diffCommits_commitValid_252=0x%0h",this.io_diffCommits_commitValid_252,rhs_.io_diffCommits_commitValid_252),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_253!=rhs_.io_diffCommits_commitValid_253) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_253=0x%0h while the rhs_.io_diffCommits_commitValid_253=0x%0h",this.io_diffCommits_commitValid_253,rhs_.io_diffCommits_commitValid_253),UVM_NONE)
        end

        if(this.io_diffCommits_commitValid_254!=rhs_.io_diffCommits_commitValid_254) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_commitValid_254=0x%0h while the rhs_.io_diffCommits_commitValid_254=0x%0h",this.io_diffCommits_commitValid_254,rhs_.io_diffCommits_commitValid_254),UVM_NONE)
        end

        if(this.io_diffCommits_info_0_ldest!=rhs_.io_diffCommits_info_0_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_0_ldest=0x%0h while the rhs_.io_diffCommits_info_0_ldest=0x%0h",this.io_diffCommits_info_0_ldest,rhs_.io_diffCommits_info_0_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_0_pdest!=rhs_.io_diffCommits_info_0_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_0_pdest=0x%0h while the rhs_.io_diffCommits_info_0_pdest=0x%0h",this.io_diffCommits_info_0_pdest,rhs_.io_diffCommits_info_0_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_0_rfWen!=rhs_.io_diffCommits_info_0_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_0_rfWen=0x%0h while the rhs_.io_diffCommits_info_0_rfWen=0x%0h",this.io_diffCommits_info_0_rfWen,rhs_.io_diffCommits_info_0_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_0_fpWen!=rhs_.io_diffCommits_info_0_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_0_fpWen=0x%0h while the rhs_.io_diffCommits_info_0_fpWen=0x%0h",this.io_diffCommits_info_0_fpWen,rhs_.io_diffCommits_info_0_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_0_vecWen!=rhs_.io_diffCommits_info_0_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_0_vecWen=0x%0h while the rhs_.io_diffCommits_info_0_vecWen=0x%0h",this.io_diffCommits_info_0_vecWen,rhs_.io_diffCommits_info_0_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_0_v0Wen!=rhs_.io_diffCommits_info_0_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_0_v0Wen=0x%0h while the rhs_.io_diffCommits_info_0_v0Wen=0x%0h",this.io_diffCommits_info_0_v0Wen,rhs_.io_diffCommits_info_0_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_0_vlWen!=rhs_.io_diffCommits_info_0_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_0_vlWen=0x%0h while the rhs_.io_diffCommits_info_0_vlWen=0x%0h",this.io_diffCommits_info_0_vlWen,rhs_.io_diffCommits_info_0_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_1_ldest!=rhs_.io_diffCommits_info_1_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_1_ldest=0x%0h while the rhs_.io_diffCommits_info_1_ldest=0x%0h",this.io_diffCommits_info_1_ldest,rhs_.io_diffCommits_info_1_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_1_pdest!=rhs_.io_diffCommits_info_1_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_1_pdest=0x%0h while the rhs_.io_diffCommits_info_1_pdest=0x%0h",this.io_diffCommits_info_1_pdest,rhs_.io_diffCommits_info_1_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_1_rfWen!=rhs_.io_diffCommits_info_1_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_1_rfWen=0x%0h while the rhs_.io_diffCommits_info_1_rfWen=0x%0h",this.io_diffCommits_info_1_rfWen,rhs_.io_diffCommits_info_1_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_1_fpWen!=rhs_.io_diffCommits_info_1_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_1_fpWen=0x%0h while the rhs_.io_diffCommits_info_1_fpWen=0x%0h",this.io_diffCommits_info_1_fpWen,rhs_.io_diffCommits_info_1_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_1_vecWen!=rhs_.io_diffCommits_info_1_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_1_vecWen=0x%0h while the rhs_.io_diffCommits_info_1_vecWen=0x%0h",this.io_diffCommits_info_1_vecWen,rhs_.io_diffCommits_info_1_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_1_v0Wen!=rhs_.io_diffCommits_info_1_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_1_v0Wen=0x%0h while the rhs_.io_diffCommits_info_1_v0Wen=0x%0h",this.io_diffCommits_info_1_v0Wen,rhs_.io_diffCommits_info_1_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_1_vlWen!=rhs_.io_diffCommits_info_1_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_1_vlWen=0x%0h while the rhs_.io_diffCommits_info_1_vlWen=0x%0h",this.io_diffCommits_info_1_vlWen,rhs_.io_diffCommits_info_1_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_2_ldest!=rhs_.io_diffCommits_info_2_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_2_ldest=0x%0h while the rhs_.io_diffCommits_info_2_ldest=0x%0h",this.io_diffCommits_info_2_ldest,rhs_.io_diffCommits_info_2_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_2_pdest!=rhs_.io_diffCommits_info_2_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_2_pdest=0x%0h while the rhs_.io_diffCommits_info_2_pdest=0x%0h",this.io_diffCommits_info_2_pdest,rhs_.io_diffCommits_info_2_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_2_rfWen!=rhs_.io_diffCommits_info_2_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_2_rfWen=0x%0h while the rhs_.io_diffCommits_info_2_rfWen=0x%0h",this.io_diffCommits_info_2_rfWen,rhs_.io_diffCommits_info_2_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_2_fpWen!=rhs_.io_diffCommits_info_2_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_2_fpWen=0x%0h while the rhs_.io_diffCommits_info_2_fpWen=0x%0h",this.io_diffCommits_info_2_fpWen,rhs_.io_diffCommits_info_2_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_2_vecWen!=rhs_.io_diffCommits_info_2_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_2_vecWen=0x%0h while the rhs_.io_diffCommits_info_2_vecWen=0x%0h",this.io_diffCommits_info_2_vecWen,rhs_.io_diffCommits_info_2_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_2_v0Wen!=rhs_.io_diffCommits_info_2_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_2_v0Wen=0x%0h while the rhs_.io_diffCommits_info_2_v0Wen=0x%0h",this.io_diffCommits_info_2_v0Wen,rhs_.io_diffCommits_info_2_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_2_vlWen!=rhs_.io_diffCommits_info_2_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_2_vlWen=0x%0h while the rhs_.io_diffCommits_info_2_vlWen=0x%0h",this.io_diffCommits_info_2_vlWen,rhs_.io_diffCommits_info_2_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_3_ldest!=rhs_.io_diffCommits_info_3_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_3_ldest=0x%0h while the rhs_.io_diffCommits_info_3_ldest=0x%0h",this.io_diffCommits_info_3_ldest,rhs_.io_diffCommits_info_3_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_3_pdest!=rhs_.io_diffCommits_info_3_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_3_pdest=0x%0h while the rhs_.io_diffCommits_info_3_pdest=0x%0h",this.io_diffCommits_info_3_pdest,rhs_.io_diffCommits_info_3_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_3_rfWen!=rhs_.io_diffCommits_info_3_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_3_rfWen=0x%0h while the rhs_.io_diffCommits_info_3_rfWen=0x%0h",this.io_diffCommits_info_3_rfWen,rhs_.io_diffCommits_info_3_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_3_fpWen!=rhs_.io_diffCommits_info_3_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_3_fpWen=0x%0h while the rhs_.io_diffCommits_info_3_fpWen=0x%0h",this.io_diffCommits_info_3_fpWen,rhs_.io_diffCommits_info_3_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_3_vecWen!=rhs_.io_diffCommits_info_3_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_3_vecWen=0x%0h while the rhs_.io_diffCommits_info_3_vecWen=0x%0h",this.io_diffCommits_info_3_vecWen,rhs_.io_diffCommits_info_3_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_3_v0Wen!=rhs_.io_diffCommits_info_3_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_3_v0Wen=0x%0h while the rhs_.io_diffCommits_info_3_v0Wen=0x%0h",this.io_diffCommits_info_3_v0Wen,rhs_.io_diffCommits_info_3_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_3_vlWen!=rhs_.io_diffCommits_info_3_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_3_vlWen=0x%0h while the rhs_.io_diffCommits_info_3_vlWen=0x%0h",this.io_diffCommits_info_3_vlWen,rhs_.io_diffCommits_info_3_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_4_ldest!=rhs_.io_diffCommits_info_4_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_4_ldest=0x%0h while the rhs_.io_diffCommits_info_4_ldest=0x%0h",this.io_diffCommits_info_4_ldest,rhs_.io_diffCommits_info_4_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_4_pdest!=rhs_.io_diffCommits_info_4_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_4_pdest=0x%0h while the rhs_.io_diffCommits_info_4_pdest=0x%0h",this.io_diffCommits_info_4_pdest,rhs_.io_diffCommits_info_4_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_4_rfWen!=rhs_.io_diffCommits_info_4_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_4_rfWen=0x%0h while the rhs_.io_diffCommits_info_4_rfWen=0x%0h",this.io_diffCommits_info_4_rfWen,rhs_.io_diffCommits_info_4_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_4_fpWen!=rhs_.io_diffCommits_info_4_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_4_fpWen=0x%0h while the rhs_.io_diffCommits_info_4_fpWen=0x%0h",this.io_diffCommits_info_4_fpWen,rhs_.io_diffCommits_info_4_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_4_vecWen!=rhs_.io_diffCommits_info_4_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_4_vecWen=0x%0h while the rhs_.io_diffCommits_info_4_vecWen=0x%0h",this.io_diffCommits_info_4_vecWen,rhs_.io_diffCommits_info_4_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_4_v0Wen!=rhs_.io_diffCommits_info_4_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_4_v0Wen=0x%0h while the rhs_.io_diffCommits_info_4_v0Wen=0x%0h",this.io_diffCommits_info_4_v0Wen,rhs_.io_diffCommits_info_4_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_4_vlWen!=rhs_.io_diffCommits_info_4_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_4_vlWen=0x%0h while the rhs_.io_diffCommits_info_4_vlWen=0x%0h",this.io_diffCommits_info_4_vlWen,rhs_.io_diffCommits_info_4_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_5_ldest!=rhs_.io_diffCommits_info_5_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_5_ldest=0x%0h while the rhs_.io_diffCommits_info_5_ldest=0x%0h",this.io_diffCommits_info_5_ldest,rhs_.io_diffCommits_info_5_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_5_pdest!=rhs_.io_diffCommits_info_5_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_5_pdest=0x%0h while the rhs_.io_diffCommits_info_5_pdest=0x%0h",this.io_diffCommits_info_5_pdest,rhs_.io_diffCommits_info_5_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_5_rfWen!=rhs_.io_diffCommits_info_5_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_5_rfWen=0x%0h while the rhs_.io_diffCommits_info_5_rfWen=0x%0h",this.io_diffCommits_info_5_rfWen,rhs_.io_diffCommits_info_5_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_5_fpWen!=rhs_.io_diffCommits_info_5_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_5_fpWen=0x%0h while the rhs_.io_diffCommits_info_5_fpWen=0x%0h",this.io_diffCommits_info_5_fpWen,rhs_.io_diffCommits_info_5_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_5_vecWen!=rhs_.io_diffCommits_info_5_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_5_vecWen=0x%0h while the rhs_.io_diffCommits_info_5_vecWen=0x%0h",this.io_diffCommits_info_5_vecWen,rhs_.io_diffCommits_info_5_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_5_v0Wen!=rhs_.io_diffCommits_info_5_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_5_v0Wen=0x%0h while the rhs_.io_diffCommits_info_5_v0Wen=0x%0h",this.io_diffCommits_info_5_v0Wen,rhs_.io_diffCommits_info_5_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_5_vlWen!=rhs_.io_diffCommits_info_5_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_5_vlWen=0x%0h while the rhs_.io_diffCommits_info_5_vlWen=0x%0h",this.io_diffCommits_info_5_vlWen,rhs_.io_diffCommits_info_5_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_6_ldest!=rhs_.io_diffCommits_info_6_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_6_ldest=0x%0h while the rhs_.io_diffCommits_info_6_ldest=0x%0h",this.io_diffCommits_info_6_ldest,rhs_.io_diffCommits_info_6_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_6_pdest!=rhs_.io_diffCommits_info_6_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_6_pdest=0x%0h while the rhs_.io_diffCommits_info_6_pdest=0x%0h",this.io_diffCommits_info_6_pdest,rhs_.io_diffCommits_info_6_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_6_rfWen!=rhs_.io_diffCommits_info_6_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_6_rfWen=0x%0h while the rhs_.io_diffCommits_info_6_rfWen=0x%0h",this.io_diffCommits_info_6_rfWen,rhs_.io_diffCommits_info_6_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_6_fpWen!=rhs_.io_diffCommits_info_6_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_6_fpWen=0x%0h while the rhs_.io_diffCommits_info_6_fpWen=0x%0h",this.io_diffCommits_info_6_fpWen,rhs_.io_diffCommits_info_6_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_6_vecWen!=rhs_.io_diffCommits_info_6_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_6_vecWen=0x%0h while the rhs_.io_diffCommits_info_6_vecWen=0x%0h",this.io_diffCommits_info_6_vecWen,rhs_.io_diffCommits_info_6_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_6_v0Wen!=rhs_.io_diffCommits_info_6_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_6_v0Wen=0x%0h while the rhs_.io_diffCommits_info_6_v0Wen=0x%0h",this.io_diffCommits_info_6_v0Wen,rhs_.io_diffCommits_info_6_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_6_vlWen!=rhs_.io_diffCommits_info_6_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_6_vlWen=0x%0h while the rhs_.io_diffCommits_info_6_vlWen=0x%0h",this.io_diffCommits_info_6_vlWen,rhs_.io_diffCommits_info_6_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_7_ldest!=rhs_.io_diffCommits_info_7_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_7_ldest=0x%0h while the rhs_.io_diffCommits_info_7_ldest=0x%0h",this.io_diffCommits_info_7_ldest,rhs_.io_diffCommits_info_7_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_7_pdest!=rhs_.io_diffCommits_info_7_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_7_pdest=0x%0h while the rhs_.io_diffCommits_info_7_pdest=0x%0h",this.io_diffCommits_info_7_pdest,rhs_.io_diffCommits_info_7_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_7_rfWen!=rhs_.io_diffCommits_info_7_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_7_rfWen=0x%0h while the rhs_.io_diffCommits_info_7_rfWen=0x%0h",this.io_diffCommits_info_7_rfWen,rhs_.io_diffCommits_info_7_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_7_fpWen!=rhs_.io_diffCommits_info_7_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_7_fpWen=0x%0h while the rhs_.io_diffCommits_info_7_fpWen=0x%0h",this.io_diffCommits_info_7_fpWen,rhs_.io_diffCommits_info_7_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_7_vecWen!=rhs_.io_diffCommits_info_7_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_7_vecWen=0x%0h while the rhs_.io_diffCommits_info_7_vecWen=0x%0h",this.io_diffCommits_info_7_vecWen,rhs_.io_diffCommits_info_7_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_7_v0Wen!=rhs_.io_diffCommits_info_7_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_7_v0Wen=0x%0h while the rhs_.io_diffCommits_info_7_v0Wen=0x%0h",this.io_diffCommits_info_7_v0Wen,rhs_.io_diffCommits_info_7_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_7_vlWen!=rhs_.io_diffCommits_info_7_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_7_vlWen=0x%0h while the rhs_.io_diffCommits_info_7_vlWen=0x%0h",this.io_diffCommits_info_7_vlWen,rhs_.io_diffCommits_info_7_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_8_ldest!=rhs_.io_diffCommits_info_8_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_8_ldest=0x%0h while the rhs_.io_diffCommits_info_8_ldest=0x%0h",this.io_diffCommits_info_8_ldest,rhs_.io_diffCommits_info_8_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_8_pdest!=rhs_.io_diffCommits_info_8_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_8_pdest=0x%0h while the rhs_.io_diffCommits_info_8_pdest=0x%0h",this.io_diffCommits_info_8_pdest,rhs_.io_diffCommits_info_8_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_8_rfWen!=rhs_.io_diffCommits_info_8_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_8_rfWen=0x%0h while the rhs_.io_diffCommits_info_8_rfWen=0x%0h",this.io_diffCommits_info_8_rfWen,rhs_.io_diffCommits_info_8_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_8_fpWen!=rhs_.io_diffCommits_info_8_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_8_fpWen=0x%0h while the rhs_.io_diffCommits_info_8_fpWen=0x%0h",this.io_diffCommits_info_8_fpWen,rhs_.io_diffCommits_info_8_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_8_vecWen!=rhs_.io_diffCommits_info_8_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_8_vecWen=0x%0h while the rhs_.io_diffCommits_info_8_vecWen=0x%0h",this.io_diffCommits_info_8_vecWen,rhs_.io_diffCommits_info_8_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_8_v0Wen!=rhs_.io_diffCommits_info_8_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_8_v0Wen=0x%0h while the rhs_.io_diffCommits_info_8_v0Wen=0x%0h",this.io_diffCommits_info_8_v0Wen,rhs_.io_diffCommits_info_8_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_8_vlWen!=rhs_.io_diffCommits_info_8_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_8_vlWen=0x%0h while the rhs_.io_diffCommits_info_8_vlWen=0x%0h",this.io_diffCommits_info_8_vlWen,rhs_.io_diffCommits_info_8_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_9_ldest!=rhs_.io_diffCommits_info_9_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_9_ldest=0x%0h while the rhs_.io_diffCommits_info_9_ldest=0x%0h",this.io_diffCommits_info_9_ldest,rhs_.io_diffCommits_info_9_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_9_pdest!=rhs_.io_diffCommits_info_9_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_9_pdest=0x%0h while the rhs_.io_diffCommits_info_9_pdest=0x%0h",this.io_diffCommits_info_9_pdest,rhs_.io_diffCommits_info_9_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_9_rfWen!=rhs_.io_diffCommits_info_9_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_9_rfWen=0x%0h while the rhs_.io_diffCommits_info_9_rfWen=0x%0h",this.io_diffCommits_info_9_rfWen,rhs_.io_diffCommits_info_9_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_9_fpWen!=rhs_.io_diffCommits_info_9_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_9_fpWen=0x%0h while the rhs_.io_diffCommits_info_9_fpWen=0x%0h",this.io_diffCommits_info_9_fpWen,rhs_.io_diffCommits_info_9_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_9_vecWen!=rhs_.io_diffCommits_info_9_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_9_vecWen=0x%0h while the rhs_.io_diffCommits_info_9_vecWen=0x%0h",this.io_diffCommits_info_9_vecWen,rhs_.io_diffCommits_info_9_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_9_v0Wen!=rhs_.io_diffCommits_info_9_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_9_v0Wen=0x%0h while the rhs_.io_diffCommits_info_9_v0Wen=0x%0h",this.io_diffCommits_info_9_v0Wen,rhs_.io_diffCommits_info_9_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_9_vlWen!=rhs_.io_diffCommits_info_9_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_9_vlWen=0x%0h while the rhs_.io_diffCommits_info_9_vlWen=0x%0h",this.io_diffCommits_info_9_vlWen,rhs_.io_diffCommits_info_9_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_10_ldest!=rhs_.io_diffCommits_info_10_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_10_ldest=0x%0h while the rhs_.io_diffCommits_info_10_ldest=0x%0h",this.io_diffCommits_info_10_ldest,rhs_.io_diffCommits_info_10_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_10_pdest!=rhs_.io_diffCommits_info_10_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_10_pdest=0x%0h while the rhs_.io_diffCommits_info_10_pdest=0x%0h",this.io_diffCommits_info_10_pdest,rhs_.io_diffCommits_info_10_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_10_rfWen!=rhs_.io_diffCommits_info_10_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_10_rfWen=0x%0h while the rhs_.io_diffCommits_info_10_rfWen=0x%0h",this.io_diffCommits_info_10_rfWen,rhs_.io_diffCommits_info_10_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_10_fpWen!=rhs_.io_diffCommits_info_10_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_10_fpWen=0x%0h while the rhs_.io_diffCommits_info_10_fpWen=0x%0h",this.io_diffCommits_info_10_fpWen,rhs_.io_diffCommits_info_10_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_10_vecWen!=rhs_.io_diffCommits_info_10_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_10_vecWen=0x%0h while the rhs_.io_diffCommits_info_10_vecWen=0x%0h",this.io_diffCommits_info_10_vecWen,rhs_.io_diffCommits_info_10_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_10_v0Wen!=rhs_.io_diffCommits_info_10_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_10_v0Wen=0x%0h while the rhs_.io_diffCommits_info_10_v0Wen=0x%0h",this.io_diffCommits_info_10_v0Wen,rhs_.io_diffCommits_info_10_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_10_vlWen!=rhs_.io_diffCommits_info_10_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_10_vlWen=0x%0h while the rhs_.io_diffCommits_info_10_vlWen=0x%0h",this.io_diffCommits_info_10_vlWen,rhs_.io_diffCommits_info_10_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_11_ldest!=rhs_.io_diffCommits_info_11_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_11_ldest=0x%0h while the rhs_.io_diffCommits_info_11_ldest=0x%0h",this.io_diffCommits_info_11_ldest,rhs_.io_diffCommits_info_11_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_11_pdest!=rhs_.io_diffCommits_info_11_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_11_pdest=0x%0h while the rhs_.io_diffCommits_info_11_pdest=0x%0h",this.io_diffCommits_info_11_pdest,rhs_.io_diffCommits_info_11_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_11_rfWen!=rhs_.io_diffCommits_info_11_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_11_rfWen=0x%0h while the rhs_.io_diffCommits_info_11_rfWen=0x%0h",this.io_diffCommits_info_11_rfWen,rhs_.io_diffCommits_info_11_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_11_fpWen!=rhs_.io_diffCommits_info_11_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_11_fpWen=0x%0h while the rhs_.io_diffCommits_info_11_fpWen=0x%0h",this.io_diffCommits_info_11_fpWen,rhs_.io_diffCommits_info_11_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_11_vecWen!=rhs_.io_diffCommits_info_11_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_11_vecWen=0x%0h while the rhs_.io_diffCommits_info_11_vecWen=0x%0h",this.io_diffCommits_info_11_vecWen,rhs_.io_diffCommits_info_11_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_11_v0Wen!=rhs_.io_diffCommits_info_11_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_11_v0Wen=0x%0h while the rhs_.io_diffCommits_info_11_v0Wen=0x%0h",this.io_diffCommits_info_11_v0Wen,rhs_.io_diffCommits_info_11_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_11_vlWen!=rhs_.io_diffCommits_info_11_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_11_vlWen=0x%0h while the rhs_.io_diffCommits_info_11_vlWen=0x%0h",this.io_diffCommits_info_11_vlWen,rhs_.io_diffCommits_info_11_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_12_ldest!=rhs_.io_diffCommits_info_12_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_12_ldest=0x%0h while the rhs_.io_diffCommits_info_12_ldest=0x%0h",this.io_diffCommits_info_12_ldest,rhs_.io_diffCommits_info_12_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_12_pdest!=rhs_.io_diffCommits_info_12_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_12_pdest=0x%0h while the rhs_.io_diffCommits_info_12_pdest=0x%0h",this.io_diffCommits_info_12_pdest,rhs_.io_diffCommits_info_12_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_12_rfWen!=rhs_.io_diffCommits_info_12_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_12_rfWen=0x%0h while the rhs_.io_diffCommits_info_12_rfWen=0x%0h",this.io_diffCommits_info_12_rfWen,rhs_.io_diffCommits_info_12_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_12_fpWen!=rhs_.io_diffCommits_info_12_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_12_fpWen=0x%0h while the rhs_.io_diffCommits_info_12_fpWen=0x%0h",this.io_diffCommits_info_12_fpWen,rhs_.io_diffCommits_info_12_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_12_vecWen!=rhs_.io_diffCommits_info_12_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_12_vecWen=0x%0h while the rhs_.io_diffCommits_info_12_vecWen=0x%0h",this.io_diffCommits_info_12_vecWen,rhs_.io_diffCommits_info_12_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_12_v0Wen!=rhs_.io_diffCommits_info_12_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_12_v0Wen=0x%0h while the rhs_.io_diffCommits_info_12_v0Wen=0x%0h",this.io_diffCommits_info_12_v0Wen,rhs_.io_diffCommits_info_12_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_12_vlWen!=rhs_.io_diffCommits_info_12_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_12_vlWen=0x%0h while the rhs_.io_diffCommits_info_12_vlWen=0x%0h",this.io_diffCommits_info_12_vlWen,rhs_.io_diffCommits_info_12_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_13_ldest!=rhs_.io_diffCommits_info_13_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_13_ldest=0x%0h while the rhs_.io_diffCommits_info_13_ldest=0x%0h",this.io_diffCommits_info_13_ldest,rhs_.io_diffCommits_info_13_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_13_pdest!=rhs_.io_diffCommits_info_13_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_13_pdest=0x%0h while the rhs_.io_diffCommits_info_13_pdest=0x%0h",this.io_diffCommits_info_13_pdest,rhs_.io_diffCommits_info_13_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_13_rfWen!=rhs_.io_diffCommits_info_13_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_13_rfWen=0x%0h while the rhs_.io_diffCommits_info_13_rfWen=0x%0h",this.io_diffCommits_info_13_rfWen,rhs_.io_diffCommits_info_13_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_13_fpWen!=rhs_.io_diffCommits_info_13_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_13_fpWen=0x%0h while the rhs_.io_diffCommits_info_13_fpWen=0x%0h",this.io_diffCommits_info_13_fpWen,rhs_.io_diffCommits_info_13_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_13_vecWen!=rhs_.io_diffCommits_info_13_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_13_vecWen=0x%0h while the rhs_.io_diffCommits_info_13_vecWen=0x%0h",this.io_diffCommits_info_13_vecWen,rhs_.io_diffCommits_info_13_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_13_v0Wen!=rhs_.io_diffCommits_info_13_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_13_v0Wen=0x%0h while the rhs_.io_diffCommits_info_13_v0Wen=0x%0h",this.io_diffCommits_info_13_v0Wen,rhs_.io_diffCommits_info_13_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_13_vlWen!=rhs_.io_diffCommits_info_13_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_13_vlWen=0x%0h while the rhs_.io_diffCommits_info_13_vlWen=0x%0h",this.io_diffCommits_info_13_vlWen,rhs_.io_diffCommits_info_13_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_14_ldest!=rhs_.io_diffCommits_info_14_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_14_ldest=0x%0h while the rhs_.io_diffCommits_info_14_ldest=0x%0h",this.io_diffCommits_info_14_ldest,rhs_.io_diffCommits_info_14_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_14_pdest!=rhs_.io_diffCommits_info_14_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_14_pdest=0x%0h while the rhs_.io_diffCommits_info_14_pdest=0x%0h",this.io_diffCommits_info_14_pdest,rhs_.io_diffCommits_info_14_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_14_rfWen!=rhs_.io_diffCommits_info_14_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_14_rfWen=0x%0h while the rhs_.io_diffCommits_info_14_rfWen=0x%0h",this.io_diffCommits_info_14_rfWen,rhs_.io_diffCommits_info_14_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_14_fpWen!=rhs_.io_diffCommits_info_14_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_14_fpWen=0x%0h while the rhs_.io_diffCommits_info_14_fpWen=0x%0h",this.io_diffCommits_info_14_fpWen,rhs_.io_diffCommits_info_14_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_14_vecWen!=rhs_.io_diffCommits_info_14_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_14_vecWen=0x%0h while the rhs_.io_diffCommits_info_14_vecWen=0x%0h",this.io_diffCommits_info_14_vecWen,rhs_.io_diffCommits_info_14_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_14_v0Wen!=rhs_.io_diffCommits_info_14_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_14_v0Wen=0x%0h while the rhs_.io_diffCommits_info_14_v0Wen=0x%0h",this.io_diffCommits_info_14_v0Wen,rhs_.io_diffCommits_info_14_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_14_vlWen!=rhs_.io_diffCommits_info_14_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_14_vlWen=0x%0h while the rhs_.io_diffCommits_info_14_vlWen=0x%0h",this.io_diffCommits_info_14_vlWen,rhs_.io_diffCommits_info_14_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_15_ldest!=rhs_.io_diffCommits_info_15_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_15_ldest=0x%0h while the rhs_.io_diffCommits_info_15_ldest=0x%0h",this.io_diffCommits_info_15_ldest,rhs_.io_diffCommits_info_15_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_15_pdest!=rhs_.io_diffCommits_info_15_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_15_pdest=0x%0h while the rhs_.io_diffCommits_info_15_pdest=0x%0h",this.io_diffCommits_info_15_pdest,rhs_.io_diffCommits_info_15_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_15_rfWen!=rhs_.io_diffCommits_info_15_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_15_rfWen=0x%0h while the rhs_.io_diffCommits_info_15_rfWen=0x%0h",this.io_diffCommits_info_15_rfWen,rhs_.io_diffCommits_info_15_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_15_fpWen!=rhs_.io_diffCommits_info_15_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_15_fpWen=0x%0h while the rhs_.io_diffCommits_info_15_fpWen=0x%0h",this.io_diffCommits_info_15_fpWen,rhs_.io_diffCommits_info_15_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_15_vecWen!=rhs_.io_diffCommits_info_15_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_15_vecWen=0x%0h while the rhs_.io_diffCommits_info_15_vecWen=0x%0h",this.io_diffCommits_info_15_vecWen,rhs_.io_diffCommits_info_15_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_15_v0Wen!=rhs_.io_diffCommits_info_15_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_15_v0Wen=0x%0h while the rhs_.io_diffCommits_info_15_v0Wen=0x%0h",this.io_diffCommits_info_15_v0Wen,rhs_.io_diffCommits_info_15_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_15_vlWen!=rhs_.io_diffCommits_info_15_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_15_vlWen=0x%0h while the rhs_.io_diffCommits_info_15_vlWen=0x%0h",this.io_diffCommits_info_15_vlWen,rhs_.io_diffCommits_info_15_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_16_ldest!=rhs_.io_diffCommits_info_16_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_16_ldest=0x%0h while the rhs_.io_diffCommits_info_16_ldest=0x%0h",this.io_diffCommits_info_16_ldest,rhs_.io_diffCommits_info_16_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_16_pdest!=rhs_.io_diffCommits_info_16_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_16_pdest=0x%0h while the rhs_.io_diffCommits_info_16_pdest=0x%0h",this.io_diffCommits_info_16_pdest,rhs_.io_diffCommits_info_16_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_16_rfWen!=rhs_.io_diffCommits_info_16_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_16_rfWen=0x%0h while the rhs_.io_diffCommits_info_16_rfWen=0x%0h",this.io_diffCommits_info_16_rfWen,rhs_.io_diffCommits_info_16_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_16_fpWen!=rhs_.io_diffCommits_info_16_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_16_fpWen=0x%0h while the rhs_.io_diffCommits_info_16_fpWen=0x%0h",this.io_diffCommits_info_16_fpWen,rhs_.io_diffCommits_info_16_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_16_vecWen!=rhs_.io_diffCommits_info_16_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_16_vecWen=0x%0h while the rhs_.io_diffCommits_info_16_vecWen=0x%0h",this.io_diffCommits_info_16_vecWen,rhs_.io_diffCommits_info_16_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_16_v0Wen!=rhs_.io_diffCommits_info_16_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_16_v0Wen=0x%0h while the rhs_.io_diffCommits_info_16_v0Wen=0x%0h",this.io_diffCommits_info_16_v0Wen,rhs_.io_diffCommits_info_16_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_16_vlWen!=rhs_.io_diffCommits_info_16_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_16_vlWen=0x%0h while the rhs_.io_diffCommits_info_16_vlWen=0x%0h",this.io_diffCommits_info_16_vlWen,rhs_.io_diffCommits_info_16_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_17_ldest!=rhs_.io_diffCommits_info_17_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_17_ldest=0x%0h while the rhs_.io_diffCommits_info_17_ldest=0x%0h",this.io_diffCommits_info_17_ldest,rhs_.io_diffCommits_info_17_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_17_pdest!=rhs_.io_diffCommits_info_17_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_17_pdest=0x%0h while the rhs_.io_diffCommits_info_17_pdest=0x%0h",this.io_diffCommits_info_17_pdest,rhs_.io_diffCommits_info_17_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_17_rfWen!=rhs_.io_diffCommits_info_17_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_17_rfWen=0x%0h while the rhs_.io_diffCommits_info_17_rfWen=0x%0h",this.io_diffCommits_info_17_rfWen,rhs_.io_diffCommits_info_17_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_17_fpWen!=rhs_.io_diffCommits_info_17_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_17_fpWen=0x%0h while the rhs_.io_diffCommits_info_17_fpWen=0x%0h",this.io_diffCommits_info_17_fpWen,rhs_.io_diffCommits_info_17_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_17_vecWen!=rhs_.io_diffCommits_info_17_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_17_vecWen=0x%0h while the rhs_.io_diffCommits_info_17_vecWen=0x%0h",this.io_diffCommits_info_17_vecWen,rhs_.io_diffCommits_info_17_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_17_v0Wen!=rhs_.io_diffCommits_info_17_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_17_v0Wen=0x%0h while the rhs_.io_diffCommits_info_17_v0Wen=0x%0h",this.io_diffCommits_info_17_v0Wen,rhs_.io_diffCommits_info_17_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_17_vlWen!=rhs_.io_diffCommits_info_17_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_17_vlWen=0x%0h while the rhs_.io_diffCommits_info_17_vlWen=0x%0h",this.io_diffCommits_info_17_vlWen,rhs_.io_diffCommits_info_17_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_18_ldest!=rhs_.io_diffCommits_info_18_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_18_ldest=0x%0h while the rhs_.io_diffCommits_info_18_ldest=0x%0h",this.io_diffCommits_info_18_ldest,rhs_.io_diffCommits_info_18_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_18_pdest!=rhs_.io_diffCommits_info_18_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_18_pdest=0x%0h while the rhs_.io_diffCommits_info_18_pdest=0x%0h",this.io_diffCommits_info_18_pdest,rhs_.io_diffCommits_info_18_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_18_rfWen!=rhs_.io_diffCommits_info_18_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_18_rfWen=0x%0h while the rhs_.io_diffCommits_info_18_rfWen=0x%0h",this.io_diffCommits_info_18_rfWen,rhs_.io_diffCommits_info_18_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_18_fpWen!=rhs_.io_diffCommits_info_18_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_18_fpWen=0x%0h while the rhs_.io_diffCommits_info_18_fpWen=0x%0h",this.io_diffCommits_info_18_fpWen,rhs_.io_diffCommits_info_18_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_18_vecWen!=rhs_.io_diffCommits_info_18_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_18_vecWen=0x%0h while the rhs_.io_diffCommits_info_18_vecWen=0x%0h",this.io_diffCommits_info_18_vecWen,rhs_.io_diffCommits_info_18_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_18_v0Wen!=rhs_.io_diffCommits_info_18_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_18_v0Wen=0x%0h while the rhs_.io_diffCommits_info_18_v0Wen=0x%0h",this.io_diffCommits_info_18_v0Wen,rhs_.io_diffCommits_info_18_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_18_vlWen!=rhs_.io_diffCommits_info_18_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_18_vlWen=0x%0h while the rhs_.io_diffCommits_info_18_vlWen=0x%0h",this.io_diffCommits_info_18_vlWen,rhs_.io_diffCommits_info_18_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_19_ldest!=rhs_.io_diffCommits_info_19_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_19_ldest=0x%0h while the rhs_.io_diffCommits_info_19_ldest=0x%0h",this.io_diffCommits_info_19_ldest,rhs_.io_diffCommits_info_19_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_19_pdest!=rhs_.io_diffCommits_info_19_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_19_pdest=0x%0h while the rhs_.io_diffCommits_info_19_pdest=0x%0h",this.io_diffCommits_info_19_pdest,rhs_.io_diffCommits_info_19_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_19_rfWen!=rhs_.io_diffCommits_info_19_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_19_rfWen=0x%0h while the rhs_.io_diffCommits_info_19_rfWen=0x%0h",this.io_diffCommits_info_19_rfWen,rhs_.io_diffCommits_info_19_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_19_fpWen!=rhs_.io_diffCommits_info_19_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_19_fpWen=0x%0h while the rhs_.io_diffCommits_info_19_fpWen=0x%0h",this.io_diffCommits_info_19_fpWen,rhs_.io_diffCommits_info_19_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_19_vecWen!=rhs_.io_diffCommits_info_19_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_19_vecWen=0x%0h while the rhs_.io_diffCommits_info_19_vecWen=0x%0h",this.io_diffCommits_info_19_vecWen,rhs_.io_diffCommits_info_19_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_19_v0Wen!=rhs_.io_diffCommits_info_19_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_19_v0Wen=0x%0h while the rhs_.io_diffCommits_info_19_v0Wen=0x%0h",this.io_diffCommits_info_19_v0Wen,rhs_.io_diffCommits_info_19_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_19_vlWen!=rhs_.io_diffCommits_info_19_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_19_vlWen=0x%0h while the rhs_.io_diffCommits_info_19_vlWen=0x%0h",this.io_diffCommits_info_19_vlWen,rhs_.io_diffCommits_info_19_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_20_ldest!=rhs_.io_diffCommits_info_20_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_20_ldest=0x%0h while the rhs_.io_diffCommits_info_20_ldest=0x%0h",this.io_diffCommits_info_20_ldest,rhs_.io_diffCommits_info_20_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_20_pdest!=rhs_.io_diffCommits_info_20_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_20_pdest=0x%0h while the rhs_.io_diffCommits_info_20_pdest=0x%0h",this.io_diffCommits_info_20_pdest,rhs_.io_diffCommits_info_20_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_20_rfWen!=rhs_.io_diffCommits_info_20_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_20_rfWen=0x%0h while the rhs_.io_diffCommits_info_20_rfWen=0x%0h",this.io_diffCommits_info_20_rfWen,rhs_.io_diffCommits_info_20_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_20_fpWen!=rhs_.io_diffCommits_info_20_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_20_fpWen=0x%0h while the rhs_.io_diffCommits_info_20_fpWen=0x%0h",this.io_diffCommits_info_20_fpWen,rhs_.io_diffCommits_info_20_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_20_vecWen!=rhs_.io_diffCommits_info_20_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_20_vecWen=0x%0h while the rhs_.io_diffCommits_info_20_vecWen=0x%0h",this.io_diffCommits_info_20_vecWen,rhs_.io_diffCommits_info_20_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_20_v0Wen!=rhs_.io_diffCommits_info_20_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_20_v0Wen=0x%0h while the rhs_.io_diffCommits_info_20_v0Wen=0x%0h",this.io_diffCommits_info_20_v0Wen,rhs_.io_diffCommits_info_20_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_20_vlWen!=rhs_.io_diffCommits_info_20_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_20_vlWen=0x%0h while the rhs_.io_diffCommits_info_20_vlWen=0x%0h",this.io_diffCommits_info_20_vlWen,rhs_.io_diffCommits_info_20_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_21_ldest!=rhs_.io_diffCommits_info_21_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_21_ldest=0x%0h while the rhs_.io_diffCommits_info_21_ldest=0x%0h",this.io_diffCommits_info_21_ldest,rhs_.io_diffCommits_info_21_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_21_pdest!=rhs_.io_diffCommits_info_21_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_21_pdest=0x%0h while the rhs_.io_diffCommits_info_21_pdest=0x%0h",this.io_diffCommits_info_21_pdest,rhs_.io_diffCommits_info_21_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_21_rfWen!=rhs_.io_diffCommits_info_21_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_21_rfWen=0x%0h while the rhs_.io_diffCommits_info_21_rfWen=0x%0h",this.io_diffCommits_info_21_rfWen,rhs_.io_diffCommits_info_21_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_21_fpWen!=rhs_.io_diffCommits_info_21_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_21_fpWen=0x%0h while the rhs_.io_diffCommits_info_21_fpWen=0x%0h",this.io_diffCommits_info_21_fpWen,rhs_.io_diffCommits_info_21_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_21_vecWen!=rhs_.io_diffCommits_info_21_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_21_vecWen=0x%0h while the rhs_.io_diffCommits_info_21_vecWen=0x%0h",this.io_diffCommits_info_21_vecWen,rhs_.io_diffCommits_info_21_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_21_v0Wen!=rhs_.io_diffCommits_info_21_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_21_v0Wen=0x%0h while the rhs_.io_diffCommits_info_21_v0Wen=0x%0h",this.io_diffCommits_info_21_v0Wen,rhs_.io_diffCommits_info_21_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_21_vlWen!=rhs_.io_diffCommits_info_21_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_21_vlWen=0x%0h while the rhs_.io_diffCommits_info_21_vlWen=0x%0h",this.io_diffCommits_info_21_vlWen,rhs_.io_diffCommits_info_21_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_22_ldest!=rhs_.io_diffCommits_info_22_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_22_ldest=0x%0h while the rhs_.io_diffCommits_info_22_ldest=0x%0h",this.io_diffCommits_info_22_ldest,rhs_.io_diffCommits_info_22_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_22_pdest!=rhs_.io_diffCommits_info_22_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_22_pdest=0x%0h while the rhs_.io_diffCommits_info_22_pdest=0x%0h",this.io_diffCommits_info_22_pdest,rhs_.io_diffCommits_info_22_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_22_rfWen!=rhs_.io_diffCommits_info_22_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_22_rfWen=0x%0h while the rhs_.io_diffCommits_info_22_rfWen=0x%0h",this.io_diffCommits_info_22_rfWen,rhs_.io_diffCommits_info_22_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_22_fpWen!=rhs_.io_diffCommits_info_22_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_22_fpWen=0x%0h while the rhs_.io_diffCommits_info_22_fpWen=0x%0h",this.io_diffCommits_info_22_fpWen,rhs_.io_diffCommits_info_22_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_22_vecWen!=rhs_.io_diffCommits_info_22_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_22_vecWen=0x%0h while the rhs_.io_diffCommits_info_22_vecWen=0x%0h",this.io_diffCommits_info_22_vecWen,rhs_.io_diffCommits_info_22_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_22_v0Wen!=rhs_.io_diffCommits_info_22_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_22_v0Wen=0x%0h while the rhs_.io_diffCommits_info_22_v0Wen=0x%0h",this.io_diffCommits_info_22_v0Wen,rhs_.io_diffCommits_info_22_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_22_vlWen!=rhs_.io_diffCommits_info_22_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_22_vlWen=0x%0h while the rhs_.io_diffCommits_info_22_vlWen=0x%0h",this.io_diffCommits_info_22_vlWen,rhs_.io_diffCommits_info_22_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_23_ldest!=rhs_.io_diffCommits_info_23_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_23_ldest=0x%0h while the rhs_.io_diffCommits_info_23_ldest=0x%0h",this.io_diffCommits_info_23_ldest,rhs_.io_diffCommits_info_23_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_23_pdest!=rhs_.io_diffCommits_info_23_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_23_pdest=0x%0h while the rhs_.io_diffCommits_info_23_pdest=0x%0h",this.io_diffCommits_info_23_pdest,rhs_.io_diffCommits_info_23_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_23_rfWen!=rhs_.io_diffCommits_info_23_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_23_rfWen=0x%0h while the rhs_.io_diffCommits_info_23_rfWen=0x%0h",this.io_diffCommits_info_23_rfWen,rhs_.io_diffCommits_info_23_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_23_fpWen!=rhs_.io_diffCommits_info_23_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_23_fpWen=0x%0h while the rhs_.io_diffCommits_info_23_fpWen=0x%0h",this.io_diffCommits_info_23_fpWen,rhs_.io_diffCommits_info_23_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_23_vecWen!=rhs_.io_diffCommits_info_23_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_23_vecWen=0x%0h while the rhs_.io_diffCommits_info_23_vecWen=0x%0h",this.io_diffCommits_info_23_vecWen,rhs_.io_diffCommits_info_23_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_23_v0Wen!=rhs_.io_diffCommits_info_23_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_23_v0Wen=0x%0h while the rhs_.io_diffCommits_info_23_v0Wen=0x%0h",this.io_diffCommits_info_23_v0Wen,rhs_.io_diffCommits_info_23_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_23_vlWen!=rhs_.io_diffCommits_info_23_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_23_vlWen=0x%0h while the rhs_.io_diffCommits_info_23_vlWen=0x%0h",this.io_diffCommits_info_23_vlWen,rhs_.io_diffCommits_info_23_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_24_ldest!=rhs_.io_diffCommits_info_24_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_24_ldest=0x%0h while the rhs_.io_diffCommits_info_24_ldest=0x%0h",this.io_diffCommits_info_24_ldest,rhs_.io_diffCommits_info_24_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_24_pdest!=rhs_.io_diffCommits_info_24_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_24_pdest=0x%0h while the rhs_.io_diffCommits_info_24_pdest=0x%0h",this.io_diffCommits_info_24_pdest,rhs_.io_diffCommits_info_24_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_24_rfWen!=rhs_.io_diffCommits_info_24_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_24_rfWen=0x%0h while the rhs_.io_diffCommits_info_24_rfWen=0x%0h",this.io_diffCommits_info_24_rfWen,rhs_.io_diffCommits_info_24_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_24_fpWen!=rhs_.io_diffCommits_info_24_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_24_fpWen=0x%0h while the rhs_.io_diffCommits_info_24_fpWen=0x%0h",this.io_diffCommits_info_24_fpWen,rhs_.io_diffCommits_info_24_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_24_vecWen!=rhs_.io_diffCommits_info_24_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_24_vecWen=0x%0h while the rhs_.io_diffCommits_info_24_vecWen=0x%0h",this.io_diffCommits_info_24_vecWen,rhs_.io_diffCommits_info_24_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_24_v0Wen!=rhs_.io_diffCommits_info_24_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_24_v0Wen=0x%0h while the rhs_.io_diffCommits_info_24_v0Wen=0x%0h",this.io_diffCommits_info_24_v0Wen,rhs_.io_diffCommits_info_24_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_24_vlWen!=rhs_.io_diffCommits_info_24_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_24_vlWen=0x%0h while the rhs_.io_diffCommits_info_24_vlWen=0x%0h",this.io_diffCommits_info_24_vlWen,rhs_.io_diffCommits_info_24_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_25_ldest!=rhs_.io_diffCommits_info_25_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_25_ldest=0x%0h while the rhs_.io_diffCommits_info_25_ldest=0x%0h",this.io_diffCommits_info_25_ldest,rhs_.io_diffCommits_info_25_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_25_pdest!=rhs_.io_diffCommits_info_25_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_25_pdest=0x%0h while the rhs_.io_diffCommits_info_25_pdest=0x%0h",this.io_diffCommits_info_25_pdest,rhs_.io_diffCommits_info_25_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_25_rfWen!=rhs_.io_diffCommits_info_25_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_25_rfWen=0x%0h while the rhs_.io_diffCommits_info_25_rfWen=0x%0h",this.io_diffCommits_info_25_rfWen,rhs_.io_diffCommits_info_25_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_25_fpWen!=rhs_.io_diffCommits_info_25_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_25_fpWen=0x%0h while the rhs_.io_diffCommits_info_25_fpWen=0x%0h",this.io_diffCommits_info_25_fpWen,rhs_.io_diffCommits_info_25_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_25_vecWen!=rhs_.io_diffCommits_info_25_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_25_vecWen=0x%0h while the rhs_.io_diffCommits_info_25_vecWen=0x%0h",this.io_diffCommits_info_25_vecWen,rhs_.io_diffCommits_info_25_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_25_v0Wen!=rhs_.io_diffCommits_info_25_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_25_v0Wen=0x%0h while the rhs_.io_diffCommits_info_25_v0Wen=0x%0h",this.io_diffCommits_info_25_v0Wen,rhs_.io_diffCommits_info_25_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_25_vlWen!=rhs_.io_diffCommits_info_25_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_25_vlWen=0x%0h while the rhs_.io_diffCommits_info_25_vlWen=0x%0h",this.io_diffCommits_info_25_vlWen,rhs_.io_diffCommits_info_25_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_26_ldest!=rhs_.io_diffCommits_info_26_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_26_ldest=0x%0h while the rhs_.io_diffCommits_info_26_ldest=0x%0h",this.io_diffCommits_info_26_ldest,rhs_.io_diffCommits_info_26_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_26_pdest!=rhs_.io_diffCommits_info_26_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_26_pdest=0x%0h while the rhs_.io_diffCommits_info_26_pdest=0x%0h",this.io_diffCommits_info_26_pdest,rhs_.io_diffCommits_info_26_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_26_rfWen!=rhs_.io_diffCommits_info_26_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_26_rfWen=0x%0h while the rhs_.io_diffCommits_info_26_rfWen=0x%0h",this.io_diffCommits_info_26_rfWen,rhs_.io_diffCommits_info_26_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_26_fpWen!=rhs_.io_diffCommits_info_26_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_26_fpWen=0x%0h while the rhs_.io_diffCommits_info_26_fpWen=0x%0h",this.io_diffCommits_info_26_fpWen,rhs_.io_diffCommits_info_26_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_26_vecWen!=rhs_.io_diffCommits_info_26_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_26_vecWen=0x%0h while the rhs_.io_diffCommits_info_26_vecWen=0x%0h",this.io_diffCommits_info_26_vecWen,rhs_.io_diffCommits_info_26_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_26_v0Wen!=rhs_.io_diffCommits_info_26_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_26_v0Wen=0x%0h while the rhs_.io_diffCommits_info_26_v0Wen=0x%0h",this.io_diffCommits_info_26_v0Wen,rhs_.io_diffCommits_info_26_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_26_vlWen!=rhs_.io_diffCommits_info_26_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_26_vlWen=0x%0h while the rhs_.io_diffCommits_info_26_vlWen=0x%0h",this.io_diffCommits_info_26_vlWen,rhs_.io_diffCommits_info_26_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_27_ldest!=rhs_.io_diffCommits_info_27_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_27_ldest=0x%0h while the rhs_.io_diffCommits_info_27_ldest=0x%0h",this.io_diffCommits_info_27_ldest,rhs_.io_diffCommits_info_27_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_27_pdest!=rhs_.io_diffCommits_info_27_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_27_pdest=0x%0h while the rhs_.io_diffCommits_info_27_pdest=0x%0h",this.io_diffCommits_info_27_pdest,rhs_.io_diffCommits_info_27_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_27_rfWen!=rhs_.io_diffCommits_info_27_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_27_rfWen=0x%0h while the rhs_.io_diffCommits_info_27_rfWen=0x%0h",this.io_diffCommits_info_27_rfWen,rhs_.io_diffCommits_info_27_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_27_fpWen!=rhs_.io_diffCommits_info_27_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_27_fpWen=0x%0h while the rhs_.io_diffCommits_info_27_fpWen=0x%0h",this.io_diffCommits_info_27_fpWen,rhs_.io_diffCommits_info_27_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_27_vecWen!=rhs_.io_diffCommits_info_27_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_27_vecWen=0x%0h while the rhs_.io_diffCommits_info_27_vecWen=0x%0h",this.io_diffCommits_info_27_vecWen,rhs_.io_diffCommits_info_27_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_27_v0Wen!=rhs_.io_diffCommits_info_27_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_27_v0Wen=0x%0h while the rhs_.io_diffCommits_info_27_v0Wen=0x%0h",this.io_diffCommits_info_27_v0Wen,rhs_.io_diffCommits_info_27_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_27_vlWen!=rhs_.io_diffCommits_info_27_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_27_vlWen=0x%0h while the rhs_.io_diffCommits_info_27_vlWen=0x%0h",this.io_diffCommits_info_27_vlWen,rhs_.io_diffCommits_info_27_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_28_ldest!=rhs_.io_diffCommits_info_28_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_28_ldest=0x%0h while the rhs_.io_diffCommits_info_28_ldest=0x%0h",this.io_diffCommits_info_28_ldest,rhs_.io_diffCommits_info_28_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_28_pdest!=rhs_.io_diffCommits_info_28_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_28_pdest=0x%0h while the rhs_.io_diffCommits_info_28_pdest=0x%0h",this.io_diffCommits_info_28_pdest,rhs_.io_diffCommits_info_28_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_28_rfWen!=rhs_.io_diffCommits_info_28_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_28_rfWen=0x%0h while the rhs_.io_diffCommits_info_28_rfWen=0x%0h",this.io_diffCommits_info_28_rfWen,rhs_.io_diffCommits_info_28_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_28_fpWen!=rhs_.io_diffCommits_info_28_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_28_fpWen=0x%0h while the rhs_.io_diffCommits_info_28_fpWen=0x%0h",this.io_diffCommits_info_28_fpWen,rhs_.io_diffCommits_info_28_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_28_vecWen!=rhs_.io_diffCommits_info_28_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_28_vecWen=0x%0h while the rhs_.io_diffCommits_info_28_vecWen=0x%0h",this.io_diffCommits_info_28_vecWen,rhs_.io_diffCommits_info_28_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_28_v0Wen!=rhs_.io_diffCommits_info_28_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_28_v0Wen=0x%0h while the rhs_.io_diffCommits_info_28_v0Wen=0x%0h",this.io_diffCommits_info_28_v0Wen,rhs_.io_diffCommits_info_28_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_28_vlWen!=rhs_.io_diffCommits_info_28_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_28_vlWen=0x%0h while the rhs_.io_diffCommits_info_28_vlWen=0x%0h",this.io_diffCommits_info_28_vlWen,rhs_.io_diffCommits_info_28_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_29_ldest!=rhs_.io_diffCommits_info_29_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_29_ldest=0x%0h while the rhs_.io_diffCommits_info_29_ldest=0x%0h",this.io_diffCommits_info_29_ldest,rhs_.io_diffCommits_info_29_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_29_pdest!=rhs_.io_diffCommits_info_29_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_29_pdest=0x%0h while the rhs_.io_diffCommits_info_29_pdest=0x%0h",this.io_diffCommits_info_29_pdest,rhs_.io_diffCommits_info_29_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_29_rfWen!=rhs_.io_diffCommits_info_29_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_29_rfWen=0x%0h while the rhs_.io_diffCommits_info_29_rfWen=0x%0h",this.io_diffCommits_info_29_rfWen,rhs_.io_diffCommits_info_29_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_29_fpWen!=rhs_.io_diffCommits_info_29_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_29_fpWen=0x%0h while the rhs_.io_diffCommits_info_29_fpWen=0x%0h",this.io_diffCommits_info_29_fpWen,rhs_.io_diffCommits_info_29_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_29_vecWen!=rhs_.io_diffCommits_info_29_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_29_vecWen=0x%0h while the rhs_.io_diffCommits_info_29_vecWen=0x%0h",this.io_diffCommits_info_29_vecWen,rhs_.io_diffCommits_info_29_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_29_v0Wen!=rhs_.io_diffCommits_info_29_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_29_v0Wen=0x%0h while the rhs_.io_diffCommits_info_29_v0Wen=0x%0h",this.io_diffCommits_info_29_v0Wen,rhs_.io_diffCommits_info_29_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_29_vlWen!=rhs_.io_diffCommits_info_29_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_29_vlWen=0x%0h while the rhs_.io_diffCommits_info_29_vlWen=0x%0h",this.io_diffCommits_info_29_vlWen,rhs_.io_diffCommits_info_29_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_30_ldest!=rhs_.io_diffCommits_info_30_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_30_ldest=0x%0h while the rhs_.io_diffCommits_info_30_ldest=0x%0h",this.io_diffCommits_info_30_ldest,rhs_.io_diffCommits_info_30_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_30_pdest!=rhs_.io_diffCommits_info_30_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_30_pdest=0x%0h while the rhs_.io_diffCommits_info_30_pdest=0x%0h",this.io_diffCommits_info_30_pdest,rhs_.io_diffCommits_info_30_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_30_rfWen!=rhs_.io_diffCommits_info_30_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_30_rfWen=0x%0h while the rhs_.io_diffCommits_info_30_rfWen=0x%0h",this.io_diffCommits_info_30_rfWen,rhs_.io_diffCommits_info_30_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_30_fpWen!=rhs_.io_diffCommits_info_30_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_30_fpWen=0x%0h while the rhs_.io_diffCommits_info_30_fpWen=0x%0h",this.io_diffCommits_info_30_fpWen,rhs_.io_diffCommits_info_30_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_30_vecWen!=rhs_.io_diffCommits_info_30_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_30_vecWen=0x%0h while the rhs_.io_diffCommits_info_30_vecWen=0x%0h",this.io_diffCommits_info_30_vecWen,rhs_.io_diffCommits_info_30_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_30_v0Wen!=rhs_.io_diffCommits_info_30_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_30_v0Wen=0x%0h while the rhs_.io_diffCommits_info_30_v0Wen=0x%0h",this.io_diffCommits_info_30_v0Wen,rhs_.io_diffCommits_info_30_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_30_vlWen!=rhs_.io_diffCommits_info_30_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_30_vlWen=0x%0h while the rhs_.io_diffCommits_info_30_vlWen=0x%0h",this.io_diffCommits_info_30_vlWen,rhs_.io_diffCommits_info_30_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_31_ldest!=rhs_.io_diffCommits_info_31_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_31_ldest=0x%0h while the rhs_.io_diffCommits_info_31_ldest=0x%0h",this.io_diffCommits_info_31_ldest,rhs_.io_diffCommits_info_31_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_31_pdest!=rhs_.io_diffCommits_info_31_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_31_pdest=0x%0h while the rhs_.io_diffCommits_info_31_pdest=0x%0h",this.io_diffCommits_info_31_pdest,rhs_.io_diffCommits_info_31_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_31_rfWen!=rhs_.io_diffCommits_info_31_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_31_rfWen=0x%0h while the rhs_.io_diffCommits_info_31_rfWen=0x%0h",this.io_diffCommits_info_31_rfWen,rhs_.io_diffCommits_info_31_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_31_fpWen!=rhs_.io_diffCommits_info_31_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_31_fpWen=0x%0h while the rhs_.io_diffCommits_info_31_fpWen=0x%0h",this.io_diffCommits_info_31_fpWen,rhs_.io_diffCommits_info_31_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_31_vecWen!=rhs_.io_diffCommits_info_31_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_31_vecWen=0x%0h while the rhs_.io_diffCommits_info_31_vecWen=0x%0h",this.io_diffCommits_info_31_vecWen,rhs_.io_diffCommits_info_31_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_31_v0Wen!=rhs_.io_diffCommits_info_31_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_31_v0Wen=0x%0h while the rhs_.io_diffCommits_info_31_v0Wen=0x%0h",this.io_diffCommits_info_31_v0Wen,rhs_.io_diffCommits_info_31_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_31_vlWen!=rhs_.io_diffCommits_info_31_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_31_vlWen=0x%0h while the rhs_.io_diffCommits_info_31_vlWen=0x%0h",this.io_diffCommits_info_31_vlWen,rhs_.io_diffCommits_info_31_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_32_ldest!=rhs_.io_diffCommits_info_32_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_32_ldest=0x%0h while the rhs_.io_diffCommits_info_32_ldest=0x%0h",this.io_diffCommits_info_32_ldest,rhs_.io_diffCommits_info_32_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_32_pdest!=rhs_.io_diffCommits_info_32_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_32_pdest=0x%0h while the rhs_.io_diffCommits_info_32_pdest=0x%0h",this.io_diffCommits_info_32_pdest,rhs_.io_diffCommits_info_32_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_32_rfWen!=rhs_.io_diffCommits_info_32_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_32_rfWen=0x%0h while the rhs_.io_diffCommits_info_32_rfWen=0x%0h",this.io_diffCommits_info_32_rfWen,rhs_.io_diffCommits_info_32_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_32_fpWen!=rhs_.io_diffCommits_info_32_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_32_fpWen=0x%0h while the rhs_.io_diffCommits_info_32_fpWen=0x%0h",this.io_diffCommits_info_32_fpWen,rhs_.io_diffCommits_info_32_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_32_vecWen!=rhs_.io_diffCommits_info_32_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_32_vecWen=0x%0h while the rhs_.io_diffCommits_info_32_vecWen=0x%0h",this.io_diffCommits_info_32_vecWen,rhs_.io_diffCommits_info_32_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_32_v0Wen!=rhs_.io_diffCommits_info_32_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_32_v0Wen=0x%0h while the rhs_.io_diffCommits_info_32_v0Wen=0x%0h",this.io_diffCommits_info_32_v0Wen,rhs_.io_diffCommits_info_32_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_32_vlWen!=rhs_.io_diffCommits_info_32_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_32_vlWen=0x%0h while the rhs_.io_diffCommits_info_32_vlWen=0x%0h",this.io_diffCommits_info_32_vlWen,rhs_.io_diffCommits_info_32_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_33_ldest!=rhs_.io_diffCommits_info_33_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_33_ldest=0x%0h while the rhs_.io_diffCommits_info_33_ldest=0x%0h",this.io_diffCommits_info_33_ldest,rhs_.io_diffCommits_info_33_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_33_pdest!=rhs_.io_diffCommits_info_33_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_33_pdest=0x%0h while the rhs_.io_diffCommits_info_33_pdest=0x%0h",this.io_diffCommits_info_33_pdest,rhs_.io_diffCommits_info_33_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_33_rfWen!=rhs_.io_diffCommits_info_33_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_33_rfWen=0x%0h while the rhs_.io_diffCommits_info_33_rfWen=0x%0h",this.io_diffCommits_info_33_rfWen,rhs_.io_diffCommits_info_33_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_33_fpWen!=rhs_.io_diffCommits_info_33_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_33_fpWen=0x%0h while the rhs_.io_diffCommits_info_33_fpWen=0x%0h",this.io_diffCommits_info_33_fpWen,rhs_.io_diffCommits_info_33_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_33_vecWen!=rhs_.io_diffCommits_info_33_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_33_vecWen=0x%0h while the rhs_.io_diffCommits_info_33_vecWen=0x%0h",this.io_diffCommits_info_33_vecWen,rhs_.io_diffCommits_info_33_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_33_v0Wen!=rhs_.io_diffCommits_info_33_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_33_v0Wen=0x%0h while the rhs_.io_diffCommits_info_33_v0Wen=0x%0h",this.io_diffCommits_info_33_v0Wen,rhs_.io_diffCommits_info_33_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_33_vlWen!=rhs_.io_diffCommits_info_33_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_33_vlWen=0x%0h while the rhs_.io_diffCommits_info_33_vlWen=0x%0h",this.io_diffCommits_info_33_vlWen,rhs_.io_diffCommits_info_33_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_34_ldest!=rhs_.io_diffCommits_info_34_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_34_ldest=0x%0h while the rhs_.io_diffCommits_info_34_ldest=0x%0h",this.io_diffCommits_info_34_ldest,rhs_.io_diffCommits_info_34_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_34_pdest!=rhs_.io_diffCommits_info_34_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_34_pdest=0x%0h while the rhs_.io_diffCommits_info_34_pdest=0x%0h",this.io_diffCommits_info_34_pdest,rhs_.io_diffCommits_info_34_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_34_rfWen!=rhs_.io_diffCommits_info_34_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_34_rfWen=0x%0h while the rhs_.io_diffCommits_info_34_rfWen=0x%0h",this.io_diffCommits_info_34_rfWen,rhs_.io_diffCommits_info_34_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_34_fpWen!=rhs_.io_diffCommits_info_34_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_34_fpWen=0x%0h while the rhs_.io_diffCommits_info_34_fpWen=0x%0h",this.io_diffCommits_info_34_fpWen,rhs_.io_diffCommits_info_34_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_34_vecWen!=rhs_.io_diffCommits_info_34_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_34_vecWen=0x%0h while the rhs_.io_diffCommits_info_34_vecWen=0x%0h",this.io_diffCommits_info_34_vecWen,rhs_.io_diffCommits_info_34_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_34_v0Wen!=rhs_.io_diffCommits_info_34_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_34_v0Wen=0x%0h while the rhs_.io_diffCommits_info_34_v0Wen=0x%0h",this.io_diffCommits_info_34_v0Wen,rhs_.io_diffCommits_info_34_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_34_vlWen!=rhs_.io_diffCommits_info_34_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_34_vlWen=0x%0h while the rhs_.io_diffCommits_info_34_vlWen=0x%0h",this.io_diffCommits_info_34_vlWen,rhs_.io_diffCommits_info_34_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_35_ldest!=rhs_.io_diffCommits_info_35_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_35_ldest=0x%0h while the rhs_.io_diffCommits_info_35_ldest=0x%0h",this.io_diffCommits_info_35_ldest,rhs_.io_diffCommits_info_35_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_35_pdest!=rhs_.io_diffCommits_info_35_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_35_pdest=0x%0h while the rhs_.io_diffCommits_info_35_pdest=0x%0h",this.io_diffCommits_info_35_pdest,rhs_.io_diffCommits_info_35_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_35_rfWen!=rhs_.io_diffCommits_info_35_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_35_rfWen=0x%0h while the rhs_.io_diffCommits_info_35_rfWen=0x%0h",this.io_diffCommits_info_35_rfWen,rhs_.io_diffCommits_info_35_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_35_fpWen!=rhs_.io_diffCommits_info_35_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_35_fpWen=0x%0h while the rhs_.io_diffCommits_info_35_fpWen=0x%0h",this.io_diffCommits_info_35_fpWen,rhs_.io_diffCommits_info_35_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_35_vecWen!=rhs_.io_diffCommits_info_35_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_35_vecWen=0x%0h while the rhs_.io_diffCommits_info_35_vecWen=0x%0h",this.io_diffCommits_info_35_vecWen,rhs_.io_diffCommits_info_35_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_35_v0Wen!=rhs_.io_diffCommits_info_35_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_35_v0Wen=0x%0h while the rhs_.io_diffCommits_info_35_v0Wen=0x%0h",this.io_diffCommits_info_35_v0Wen,rhs_.io_diffCommits_info_35_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_35_vlWen!=rhs_.io_diffCommits_info_35_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_35_vlWen=0x%0h while the rhs_.io_diffCommits_info_35_vlWen=0x%0h",this.io_diffCommits_info_35_vlWen,rhs_.io_diffCommits_info_35_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_36_ldest!=rhs_.io_diffCommits_info_36_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_36_ldest=0x%0h while the rhs_.io_diffCommits_info_36_ldest=0x%0h",this.io_diffCommits_info_36_ldest,rhs_.io_diffCommits_info_36_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_36_pdest!=rhs_.io_diffCommits_info_36_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_36_pdest=0x%0h while the rhs_.io_diffCommits_info_36_pdest=0x%0h",this.io_diffCommits_info_36_pdest,rhs_.io_diffCommits_info_36_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_36_rfWen!=rhs_.io_diffCommits_info_36_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_36_rfWen=0x%0h while the rhs_.io_diffCommits_info_36_rfWen=0x%0h",this.io_diffCommits_info_36_rfWen,rhs_.io_diffCommits_info_36_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_36_fpWen!=rhs_.io_diffCommits_info_36_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_36_fpWen=0x%0h while the rhs_.io_diffCommits_info_36_fpWen=0x%0h",this.io_diffCommits_info_36_fpWen,rhs_.io_diffCommits_info_36_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_36_vecWen!=rhs_.io_diffCommits_info_36_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_36_vecWen=0x%0h while the rhs_.io_diffCommits_info_36_vecWen=0x%0h",this.io_diffCommits_info_36_vecWen,rhs_.io_diffCommits_info_36_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_36_v0Wen!=rhs_.io_diffCommits_info_36_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_36_v0Wen=0x%0h while the rhs_.io_diffCommits_info_36_v0Wen=0x%0h",this.io_diffCommits_info_36_v0Wen,rhs_.io_diffCommits_info_36_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_36_vlWen!=rhs_.io_diffCommits_info_36_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_36_vlWen=0x%0h while the rhs_.io_diffCommits_info_36_vlWen=0x%0h",this.io_diffCommits_info_36_vlWen,rhs_.io_diffCommits_info_36_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_37_ldest!=rhs_.io_diffCommits_info_37_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_37_ldest=0x%0h while the rhs_.io_diffCommits_info_37_ldest=0x%0h",this.io_diffCommits_info_37_ldest,rhs_.io_diffCommits_info_37_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_37_pdest!=rhs_.io_diffCommits_info_37_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_37_pdest=0x%0h while the rhs_.io_diffCommits_info_37_pdest=0x%0h",this.io_diffCommits_info_37_pdest,rhs_.io_diffCommits_info_37_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_37_rfWen!=rhs_.io_diffCommits_info_37_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_37_rfWen=0x%0h while the rhs_.io_diffCommits_info_37_rfWen=0x%0h",this.io_diffCommits_info_37_rfWen,rhs_.io_diffCommits_info_37_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_37_fpWen!=rhs_.io_diffCommits_info_37_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_37_fpWen=0x%0h while the rhs_.io_diffCommits_info_37_fpWen=0x%0h",this.io_diffCommits_info_37_fpWen,rhs_.io_diffCommits_info_37_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_37_vecWen!=rhs_.io_diffCommits_info_37_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_37_vecWen=0x%0h while the rhs_.io_diffCommits_info_37_vecWen=0x%0h",this.io_diffCommits_info_37_vecWen,rhs_.io_diffCommits_info_37_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_37_v0Wen!=rhs_.io_diffCommits_info_37_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_37_v0Wen=0x%0h while the rhs_.io_diffCommits_info_37_v0Wen=0x%0h",this.io_diffCommits_info_37_v0Wen,rhs_.io_diffCommits_info_37_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_37_vlWen!=rhs_.io_diffCommits_info_37_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_37_vlWen=0x%0h while the rhs_.io_diffCommits_info_37_vlWen=0x%0h",this.io_diffCommits_info_37_vlWen,rhs_.io_diffCommits_info_37_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_38_ldest!=rhs_.io_diffCommits_info_38_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_38_ldest=0x%0h while the rhs_.io_diffCommits_info_38_ldest=0x%0h",this.io_diffCommits_info_38_ldest,rhs_.io_diffCommits_info_38_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_38_pdest!=rhs_.io_diffCommits_info_38_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_38_pdest=0x%0h while the rhs_.io_diffCommits_info_38_pdest=0x%0h",this.io_diffCommits_info_38_pdest,rhs_.io_diffCommits_info_38_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_38_rfWen!=rhs_.io_diffCommits_info_38_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_38_rfWen=0x%0h while the rhs_.io_diffCommits_info_38_rfWen=0x%0h",this.io_diffCommits_info_38_rfWen,rhs_.io_diffCommits_info_38_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_38_fpWen!=rhs_.io_diffCommits_info_38_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_38_fpWen=0x%0h while the rhs_.io_diffCommits_info_38_fpWen=0x%0h",this.io_diffCommits_info_38_fpWen,rhs_.io_diffCommits_info_38_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_38_vecWen!=rhs_.io_diffCommits_info_38_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_38_vecWen=0x%0h while the rhs_.io_diffCommits_info_38_vecWen=0x%0h",this.io_diffCommits_info_38_vecWen,rhs_.io_diffCommits_info_38_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_38_v0Wen!=rhs_.io_diffCommits_info_38_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_38_v0Wen=0x%0h while the rhs_.io_diffCommits_info_38_v0Wen=0x%0h",this.io_diffCommits_info_38_v0Wen,rhs_.io_diffCommits_info_38_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_38_vlWen!=rhs_.io_diffCommits_info_38_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_38_vlWen=0x%0h while the rhs_.io_diffCommits_info_38_vlWen=0x%0h",this.io_diffCommits_info_38_vlWen,rhs_.io_diffCommits_info_38_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_39_ldest!=rhs_.io_diffCommits_info_39_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_39_ldest=0x%0h while the rhs_.io_diffCommits_info_39_ldest=0x%0h",this.io_diffCommits_info_39_ldest,rhs_.io_diffCommits_info_39_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_39_pdest!=rhs_.io_diffCommits_info_39_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_39_pdest=0x%0h while the rhs_.io_diffCommits_info_39_pdest=0x%0h",this.io_diffCommits_info_39_pdest,rhs_.io_diffCommits_info_39_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_39_rfWen!=rhs_.io_diffCommits_info_39_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_39_rfWen=0x%0h while the rhs_.io_diffCommits_info_39_rfWen=0x%0h",this.io_diffCommits_info_39_rfWen,rhs_.io_diffCommits_info_39_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_39_fpWen!=rhs_.io_diffCommits_info_39_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_39_fpWen=0x%0h while the rhs_.io_diffCommits_info_39_fpWen=0x%0h",this.io_diffCommits_info_39_fpWen,rhs_.io_diffCommits_info_39_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_39_vecWen!=rhs_.io_diffCommits_info_39_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_39_vecWen=0x%0h while the rhs_.io_diffCommits_info_39_vecWen=0x%0h",this.io_diffCommits_info_39_vecWen,rhs_.io_diffCommits_info_39_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_39_v0Wen!=rhs_.io_diffCommits_info_39_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_39_v0Wen=0x%0h while the rhs_.io_diffCommits_info_39_v0Wen=0x%0h",this.io_diffCommits_info_39_v0Wen,rhs_.io_diffCommits_info_39_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_39_vlWen!=rhs_.io_diffCommits_info_39_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_39_vlWen=0x%0h while the rhs_.io_diffCommits_info_39_vlWen=0x%0h",this.io_diffCommits_info_39_vlWen,rhs_.io_diffCommits_info_39_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_40_ldest!=rhs_.io_diffCommits_info_40_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_40_ldest=0x%0h while the rhs_.io_diffCommits_info_40_ldest=0x%0h",this.io_diffCommits_info_40_ldest,rhs_.io_diffCommits_info_40_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_40_pdest!=rhs_.io_diffCommits_info_40_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_40_pdest=0x%0h while the rhs_.io_diffCommits_info_40_pdest=0x%0h",this.io_diffCommits_info_40_pdest,rhs_.io_diffCommits_info_40_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_40_rfWen!=rhs_.io_diffCommits_info_40_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_40_rfWen=0x%0h while the rhs_.io_diffCommits_info_40_rfWen=0x%0h",this.io_diffCommits_info_40_rfWen,rhs_.io_diffCommits_info_40_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_40_fpWen!=rhs_.io_diffCommits_info_40_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_40_fpWen=0x%0h while the rhs_.io_diffCommits_info_40_fpWen=0x%0h",this.io_diffCommits_info_40_fpWen,rhs_.io_diffCommits_info_40_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_40_vecWen!=rhs_.io_diffCommits_info_40_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_40_vecWen=0x%0h while the rhs_.io_diffCommits_info_40_vecWen=0x%0h",this.io_diffCommits_info_40_vecWen,rhs_.io_diffCommits_info_40_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_40_v0Wen!=rhs_.io_diffCommits_info_40_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_40_v0Wen=0x%0h while the rhs_.io_diffCommits_info_40_v0Wen=0x%0h",this.io_diffCommits_info_40_v0Wen,rhs_.io_diffCommits_info_40_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_40_vlWen!=rhs_.io_diffCommits_info_40_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_40_vlWen=0x%0h while the rhs_.io_diffCommits_info_40_vlWen=0x%0h",this.io_diffCommits_info_40_vlWen,rhs_.io_diffCommits_info_40_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_41_ldest!=rhs_.io_diffCommits_info_41_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_41_ldest=0x%0h while the rhs_.io_diffCommits_info_41_ldest=0x%0h",this.io_diffCommits_info_41_ldest,rhs_.io_diffCommits_info_41_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_41_pdest!=rhs_.io_diffCommits_info_41_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_41_pdest=0x%0h while the rhs_.io_diffCommits_info_41_pdest=0x%0h",this.io_diffCommits_info_41_pdest,rhs_.io_diffCommits_info_41_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_41_rfWen!=rhs_.io_diffCommits_info_41_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_41_rfWen=0x%0h while the rhs_.io_diffCommits_info_41_rfWen=0x%0h",this.io_diffCommits_info_41_rfWen,rhs_.io_diffCommits_info_41_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_41_fpWen!=rhs_.io_diffCommits_info_41_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_41_fpWen=0x%0h while the rhs_.io_diffCommits_info_41_fpWen=0x%0h",this.io_diffCommits_info_41_fpWen,rhs_.io_diffCommits_info_41_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_41_vecWen!=rhs_.io_diffCommits_info_41_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_41_vecWen=0x%0h while the rhs_.io_diffCommits_info_41_vecWen=0x%0h",this.io_diffCommits_info_41_vecWen,rhs_.io_diffCommits_info_41_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_41_v0Wen!=rhs_.io_diffCommits_info_41_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_41_v0Wen=0x%0h while the rhs_.io_diffCommits_info_41_v0Wen=0x%0h",this.io_diffCommits_info_41_v0Wen,rhs_.io_diffCommits_info_41_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_41_vlWen!=rhs_.io_diffCommits_info_41_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_41_vlWen=0x%0h while the rhs_.io_diffCommits_info_41_vlWen=0x%0h",this.io_diffCommits_info_41_vlWen,rhs_.io_diffCommits_info_41_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_42_ldest!=rhs_.io_diffCommits_info_42_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_42_ldest=0x%0h while the rhs_.io_diffCommits_info_42_ldest=0x%0h",this.io_diffCommits_info_42_ldest,rhs_.io_diffCommits_info_42_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_42_pdest!=rhs_.io_diffCommits_info_42_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_42_pdest=0x%0h while the rhs_.io_diffCommits_info_42_pdest=0x%0h",this.io_diffCommits_info_42_pdest,rhs_.io_diffCommits_info_42_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_42_rfWen!=rhs_.io_diffCommits_info_42_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_42_rfWen=0x%0h while the rhs_.io_diffCommits_info_42_rfWen=0x%0h",this.io_diffCommits_info_42_rfWen,rhs_.io_diffCommits_info_42_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_42_fpWen!=rhs_.io_diffCommits_info_42_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_42_fpWen=0x%0h while the rhs_.io_diffCommits_info_42_fpWen=0x%0h",this.io_diffCommits_info_42_fpWen,rhs_.io_diffCommits_info_42_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_42_vecWen!=rhs_.io_diffCommits_info_42_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_42_vecWen=0x%0h while the rhs_.io_diffCommits_info_42_vecWen=0x%0h",this.io_diffCommits_info_42_vecWen,rhs_.io_diffCommits_info_42_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_42_v0Wen!=rhs_.io_diffCommits_info_42_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_42_v0Wen=0x%0h while the rhs_.io_diffCommits_info_42_v0Wen=0x%0h",this.io_diffCommits_info_42_v0Wen,rhs_.io_diffCommits_info_42_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_42_vlWen!=rhs_.io_diffCommits_info_42_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_42_vlWen=0x%0h while the rhs_.io_diffCommits_info_42_vlWen=0x%0h",this.io_diffCommits_info_42_vlWen,rhs_.io_diffCommits_info_42_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_43_ldest!=rhs_.io_diffCommits_info_43_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_43_ldest=0x%0h while the rhs_.io_diffCommits_info_43_ldest=0x%0h",this.io_diffCommits_info_43_ldest,rhs_.io_diffCommits_info_43_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_43_pdest!=rhs_.io_diffCommits_info_43_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_43_pdest=0x%0h while the rhs_.io_diffCommits_info_43_pdest=0x%0h",this.io_diffCommits_info_43_pdest,rhs_.io_diffCommits_info_43_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_43_rfWen!=rhs_.io_diffCommits_info_43_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_43_rfWen=0x%0h while the rhs_.io_diffCommits_info_43_rfWen=0x%0h",this.io_diffCommits_info_43_rfWen,rhs_.io_diffCommits_info_43_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_43_fpWen!=rhs_.io_diffCommits_info_43_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_43_fpWen=0x%0h while the rhs_.io_diffCommits_info_43_fpWen=0x%0h",this.io_diffCommits_info_43_fpWen,rhs_.io_diffCommits_info_43_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_43_vecWen!=rhs_.io_diffCommits_info_43_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_43_vecWen=0x%0h while the rhs_.io_diffCommits_info_43_vecWen=0x%0h",this.io_diffCommits_info_43_vecWen,rhs_.io_diffCommits_info_43_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_43_v0Wen!=rhs_.io_diffCommits_info_43_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_43_v0Wen=0x%0h while the rhs_.io_diffCommits_info_43_v0Wen=0x%0h",this.io_diffCommits_info_43_v0Wen,rhs_.io_diffCommits_info_43_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_43_vlWen!=rhs_.io_diffCommits_info_43_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_43_vlWen=0x%0h while the rhs_.io_diffCommits_info_43_vlWen=0x%0h",this.io_diffCommits_info_43_vlWen,rhs_.io_diffCommits_info_43_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_44_ldest!=rhs_.io_diffCommits_info_44_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_44_ldest=0x%0h while the rhs_.io_diffCommits_info_44_ldest=0x%0h",this.io_diffCommits_info_44_ldest,rhs_.io_diffCommits_info_44_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_44_pdest!=rhs_.io_diffCommits_info_44_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_44_pdest=0x%0h while the rhs_.io_diffCommits_info_44_pdest=0x%0h",this.io_diffCommits_info_44_pdest,rhs_.io_diffCommits_info_44_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_44_rfWen!=rhs_.io_diffCommits_info_44_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_44_rfWen=0x%0h while the rhs_.io_diffCommits_info_44_rfWen=0x%0h",this.io_diffCommits_info_44_rfWen,rhs_.io_diffCommits_info_44_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_44_fpWen!=rhs_.io_diffCommits_info_44_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_44_fpWen=0x%0h while the rhs_.io_diffCommits_info_44_fpWen=0x%0h",this.io_diffCommits_info_44_fpWen,rhs_.io_diffCommits_info_44_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_44_vecWen!=rhs_.io_diffCommits_info_44_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_44_vecWen=0x%0h while the rhs_.io_diffCommits_info_44_vecWen=0x%0h",this.io_diffCommits_info_44_vecWen,rhs_.io_diffCommits_info_44_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_44_v0Wen!=rhs_.io_diffCommits_info_44_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_44_v0Wen=0x%0h while the rhs_.io_diffCommits_info_44_v0Wen=0x%0h",this.io_diffCommits_info_44_v0Wen,rhs_.io_diffCommits_info_44_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_44_vlWen!=rhs_.io_diffCommits_info_44_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_44_vlWen=0x%0h while the rhs_.io_diffCommits_info_44_vlWen=0x%0h",this.io_diffCommits_info_44_vlWen,rhs_.io_diffCommits_info_44_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_45_ldest!=rhs_.io_diffCommits_info_45_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_45_ldest=0x%0h while the rhs_.io_diffCommits_info_45_ldest=0x%0h",this.io_diffCommits_info_45_ldest,rhs_.io_diffCommits_info_45_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_45_pdest!=rhs_.io_diffCommits_info_45_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_45_pdest=0x%0h while the rhs_.io_diffCommits_info_45_pdest=0x%0h",this.io_diffCommits_info_45_pdest,rhs_.io_diffCommits_info_45_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_45_rfWen!=rhs_.io_diffCommits_info_45_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_45_rfWen=0x%0h while the rhs_.io_diffCommits_info_45_rfWen=0x%0h",this.io_diffCommits_info_45_rfWen,rhs_.io_diffCommits_info_45_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_45_fpWen!=rhs_.io_diffCommits_info_45_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_45_fpWen=0x%0h while the rhs_.io_diffCommits_info_45_fpWen=0x%0h",this.io_diffCommits_info_45_fpWen,rhs_.io_diffCommits_info_45_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_45_vecWen!=rhs_.io_diffCommits_info_45_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_45_vecWen=0x%0h while the rhs_.io_diffCommits_info_45_vecWen=0x%0h",this.io_diffCommits_info_45_vecWen,rhs_.io_diffCommits_info_45_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_45_v0Wen!=rhs_.io_diffCommits_info_45_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_45_v0Wen=0x%0h while the rhs_.io_diffCommits_info_45_v0Wen=0x%0h",this.io_diffCommits_info_45_v0Wen,rhs_.io_diffCommits_info_45_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_45_vlWen!=rhs_.io_diffCommits_info_45_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_45_vlWen=0x%0h while the rhs_.io_diffCommits_info_45_vlWen=0x%0h",this.io_diffCommits_info_45_vlWen,rhs_.io_diffCommits_info_45_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_46_ldest!=rhs_.io_diffCommits_info_46_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_46_ldest=0x%0h while the rhs_.io_diffCommits_info_46_ldest=0x%0h",this.io_diffCommits_info_46_ldest,rhs_.io_diffCommits_info_46_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_46_pdest!=rhs_.io_diffCommits_info_46_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_46_pdest=0x%0h while the rhs_.io_diffCommits_info_46_pdest=0x%0h",this.io_diffCommits_info_46_pdest,rhs_.io_diffCommits_info_46_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_46_rfWen!=rhs_.io_diffCommits_info_46_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_46_rfWen=0x%0h while the rhs_.io_diffCommits_info_46_rfWen=0x%0h",this.io_diffCommits_info_46_rfWen,rhs_.io_diffCommits_info_46_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_46_fpWen!=rhs_.io_diffCommits_info_46_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_46_fpWen=0x%0h while the rhs_.io_diffCommits_info_46_fpWen=0x%0h",this.io_diffCommits_info_46_fpWen,rhs_.io_diffCommits_info_46_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_46_vecWen!=rhs_.io_diffCommits_info_46_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_46_vecWen=0x%0h while the rhs_.io_diffCommits_info_46_vecWen=0x%0h",this.io_diffCommits_info_46_vecWen,rhs_.io_diffCommits_info_46_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_46_v0Wen!=rhs_.io_diffCommits_info_46_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_46_v0Wen=0x%0h while the rhs_.io_diffCommits_info_46_v0Wen=0x%0h",this.io_diffCommits_info_46_v0Wen,rhs_.io_diffCommits_info_46_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_46_vlWen!=rhs_.io_diffCommits_info_46_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_46_vlWen=0x%0h while the rhs_.io_diffCommits_info_46_vlWen=0x%0h",this.io_diffCommits_info_46_vlWen,rhs_.io_diffCommits_info_46_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_47_ldest!=rhs_.io_diffCommits_info_47_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_47_ldest=0x%0h while the rhs_.io_diffCommits_info_47_ldest=0x%0h",this.io_diffCommits_info_47_ldest,rhs_.io_diffCommits_info_47_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_47_pdest!=rhs_.io_diffCommits_info_47_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_47_pdest=0x%0h while the rhs_.io_diffCommits_info_47_pdest=0x%0h",this.io_diffCommits_info_47_pdest,rhs_.io_diffCommits_info_47_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_47_rfWen!=rhs_.io_diffCommits_info_47_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_47_rfWen=0x%0h while the rhs_.io_diffCommits_info_47_rfWen=0x%0h",this.io_diffCommits_info_47_rfWen,rhs_.io_diffCommits_info_47_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_47_fpWen!=rhs_.io_diffCommits_info_47_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_47_fpWen=0x%0h while the rhs_.io_diffCommits_info_47_fpWen=0x%0h",this.io_diffCommits_info_47_fpWen,rhs_.io_diffCommits_info_47_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_47_vecWen!=rhs_.io_diffCommits_info_47_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_47_vecWen=0x%0h while the rhs_.io_diffCommits_info_47_vecWen=0x%0h",this.io_diffCommits_info_47_vecWen,rhs_.io_diffCommits_info_47_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_47_v0Wen!=rhs_.io_diffCommits_info_47_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_47_v0Wen=0x%0h while the rhs_.io_diffCommits_info_47_v0Wen=0x%0h",this.io_diffCommits_info_47_v0Wen,rhs_.io_diffCommits_info_47_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_47_vlWen!=rhs_.io_diffCommits_info_47_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_47_vlWen=0x%0h while the rhs_.io_diffCommits_info_47_vlWen=0x%0h",this.io_diffCommits_info_47_vlWen,rhs_.io_diffCommits_info_47_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_48_ldest!=rhs_.io_diffCommits_info_48_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_48_ldest=0x%0h while the rhs_.io_diffCommits_info_48_ldest=0x%0h",this.io_diffCommits_info_48_ldest,rhs_.io_diffCommits_info_48_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_48_pdest!=rhs_.io_diffCommits_info_48_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_48_pdest=0x%0h while the rhs_.io_diffCommits_info_48_pdest=0x%0h",this.io_diffCommits_info_48_pdest,rhs_.io_diffCommits_info_48_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_48_rfWen!=rhs_.io_diffCommits_info_48_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_48_rfWen=0x%0h while the rhs_.io_diffCommits_info_48_rfWen=0x%0h",this.io_diffCommits_info_48_rfWen,rhs_.io_diffCommits_info_48_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_48_fpWen!=rhs_.io_diffCommits_info_48_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_48_fpWen=0x%0h while the rhs_.io_diffCommits_info_48_fpWen=0x%0h",this.io_diffCommits_info_48_fpWen,rhs_.io_diffCommits_info_48_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_48_vecWen!=rhs_.io_diffCommits_info_48_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_48_vecWen=0x%0h while the rhs_.io_diffCommits_info_48_vecWen=0x%0h",this.io_diffCommits_info_48_vecWen,rhs_.io_diffCommits_info_48_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_48_v0Wen!=rhs_.io_diffCommits_info_48_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_48_v0Wen=0x%0h while the rhs_.io_diffCommits_info_48_v0Wen=0x%0h",this.io_diffCommits_info_48_v0Wen,rhs_.io_diffCommits_info_48_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_48_vlWen!=rhs_.io_diffCommits_info_48_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_48_vlWen=0x%0h while the rhs_.io_diffCommits_info_48_vlWen=0x%0h",this.io_diffCommits_info_48_vlWen,rhs_.io_diffCommits_info_48_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_49_ldest!=rhs_.io_diffCommits_info_49_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_49_ldest=0x%0h while the rhs_.io_diffCommits_info_49_ldest=0x%0h",this.io_diffCommits_info_49_ldest,rhs_.io_diffCommits_info_49_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_49_pdest!=rhs_.io_diffCommits_info_49_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_49_pdest=0x%0h while the rhs_.io_diffCommits_info_49_pdest=0x%0h",this.io_diffCommits_info_49_pdest,rhs_.io_diffCommits_info_49_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_49_rfWen!=rhs_.io_diffCommits_info_49_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_49_rfWen=0x%0h while the rhs_.io_diffCommits_info_49_rfWen=0x%0h",this.io_diffCommits_info_49_rfWen,rhs_.io_diffCommits_info_49_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_49_fpWen!=rhs_.io_diffCommits_info_49_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_49_fpWen=0x%0h while the rhs_.io_diffCommits_info_49_fpWen=0x%0h",this.io_diffCommits_info_49_fpWen,rhs_.io_diffCommits_info_49_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_49_vecWen!=rhs_.io_diffCommits_info_49_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_49_vecWen=0x%0h while the rhs_.io_diffCommits_info_49_vecWen=0x%0h",this.io_diffCommits_info_49_vecWen,rhs_.io_diffCommits_info_49_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_49_v0Wen!=rhs_.io_diffCommits_info_49_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_49_v0Wen=0x%0h while the rhs_.io_diffCommits_info_49_v0Wen=0x%0h",this.io_diffCommits_info_49_v0Wen,rhs_.io_diffCommits_info_49_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_49_vlWen!=rhs_.io_diffCommits_info_49_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_49_vlWen=0x%0h while the rhs_.io_diffCommits_info_49_vlWen=0x%0h",this.io_diffCommits_info_49_vlWen,rhs_.io_diffCommits_info_49_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_50_ldest!=rhs_.io_diffCommits_info_50_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_50_ldest=0x%0h while the rhs_.io_diffCommits_info_50_ldest=0x%0h",this.io_diffCommits_info_50_ldest,rhs_.io_diffCommits_info_50_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_50_pdest!=rhs_.io_diffCommits_info_50_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_50_pdest=0x%0h while the rhs_.io_diffCommits_info_50_pdest=0x%0h",this.io_diffCommits_info_50_pdest,rhs_.io_diffCommits_info_50_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_50_rfWen!=rhs_.io_diffCommits_info_50_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_50_rfWen=0x%0h while the rhs_.io_diffCommits_info_50_rfWen=0x%0h",this.io_diffCommits_info_50_rfWen,rhs_.io_diffCommits_info_50_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_50_fpWen!=rhs_.io_diffCommits_info_50_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_50_fpWen=0x%0h while the rhs_.io_diffCommits_info_50_fpWen=0x%0h",this.io_diffCommits_info_50_fpWen,rhs_.io_diffCommits_info_50_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_50_vecWen!=rhs_.io_diffCommits_info_50_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_50_vecWen=0x%0h while the rhs_.io_diffCommits_info_50_vecWen=0x%0h",this.io_diffCommits_info_50_vecWen,rhs_.io_diffCommits_info_50_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_50_v0Wen!=rhs_.io_diffCommits_info_50_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_50_v0Wen=0x%0h while the rhs_.io_diffCommits_info_50_v0Wen=0x%0h",this.io_diffCommits_info_50_v0Wen,rhs_.io_diffCommits_info_50_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_50_vlWen!=rhs_.io_diffCommits_info_50_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_50_vlWen=0x%0h while the rhs_.io_diffCommits_info_50_vlWen=0x%0h",this.io_diffCommits_info_50_vlWen,rhs_.io_diffCommits_info_50_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_51_ldest!=rhs_.io_diffCommits_info_51_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_51_ldest=0x%0h while the rhs_.io_diffCommits_info_51_ldest=0x%0h",this.io_diffCommits_info_51_ldest,rhs_.io_diffCommits_info_51_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_51_pdest!=rhs_.io_diffCommits_info_51_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_51_pdest=0x%0h while the rhs_.io_diffCommits_info_51_pdest=0x%0h",this.io_diffCommits_info_51_pdest,rhs_.io_diffCommits_info_51_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_51_rfWen!=rhs_.io_diffCommits_info_51_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_51_rfWen=0x%0h while the rhs_.io_diffCommits_info_51_rfWen=0x%0h",this.io_diffCommits_info_51_rfWen,rhs_.io_diffCommits_info_51_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_51_fpWen!=rhs_.io_diffCommits_info_51_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_51_fpWen=0x%0h while the rhs_.io_diffCommits_info_51_fpWen=0x%0h",this.io_diffCommits_info_51_fpWen,rhs_.io_diffCommits_info_51_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_51_vecWen!=rhs_.io_diffCommits_info_51_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_51_vecWen=0x%0h while the rhs_.io_diffCommits_info_51_vecWen=0x%0h",this.io_diffCommits_info_51_vecWen,rhs_.io_diffCommits_info_51_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_51_v0Wen!=rhs_.io_diffCommits_info_51_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_51_v0Wen=0x%0h while the rhs_.io_diffCommits_info_51_v0Wen=0x%0h",this.io_diffCommits_info_51_v0Wen,rhs_.io_diffCommits_info_51_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_51_vlWen!=rhs_.io_diffCommits_info_51_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_51_vlWen=0x%0h while the rhs_.io_diffCommits_info_51_vlWen=0x%0h",this.io_diffCommits_info_51_vlWen,rhs_.io_diffCommits_info_51_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_52_ldest!=rhs_.io_diffCommits_info_52_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_52_ldest=0x%0h while the rhs_.io_diffCommits_info_52_ldest=0x%0h",this.io_diffCommits_info_52_ldest,rhs_.io_diffCommits_info_52_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_52_pdest!=rhs_.io_diffCommits_info_52_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_52_pdest=0x%0h while the rhs_.io_diffCommits_info_52_pdest=0x%0h",this.io_diffCommits_info_52_pdest,rhs_.io_diffCommits_info_52_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_52_rfWen!=rhs_.io_diffCommits_info_52_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_52_rfWen=0x%0h while the rhs_.io_diffCommits_info_52_rfWen=0x%0h",this.io_diffCommits_info_52_rfWen,rhs_.io_diffCommits_info_52_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_52_fpWen!=rhs_.io_diffCommits_info_52_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_52_fpWen=0x%0h while the rhs_.io_diffCommits_info_52_fpWen=0x%0h",this.io_diffCommits_info_52_fpWen,rhs_.io_diffCommits_info_52_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_52_vecWen!=rhs_.io_diffCommits_info_52_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_52_vecWen=0x%0h while the rhs_.io_diffCommits_info_52_vecWen=0x%0h",this.io_diffCommits_info_52_vecWen,rhs_.io_diffCommits_info_52_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_52_v0Wen!=rhs_.io_diffCommits_info_52_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_52_v0Wen=0x%0h while the rhs_.io_diffCommits_info_52_v0Wen=0x%0h",this.io_diffCommits_info_52_v0Wen,rhs_.io_diffCommits_info_52_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_52_vlWen!=rhs_.io_diffCommits_info_52_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_52_vlWen=0x%0h while the rhs_.io_diffCommits_info_52_vlWen=0x%0h",this.io_diffCommits_info_52_vlWen,rhs_.io_diffCommits_info_52_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_53_ldest!=rhs_.io_diffCommits_info_53_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_53_ldest=0x%0h while the rhs_.io_diffCommits_info_53_ldest=0x%0h",this.io_diffCommits_info_53_ldest,rhs_.io_diffCommits_info_53_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_53_pdest!=rhs_.io_diffCommits_info_53_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_53_pdest=0x%0h while the rhs_.io_diffCommits_info_53_pdest=0x%0h",this.io_diffCommits_info_53_pdest,rhs_.io_diffCommits_info_53_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_53_rfWen!=rhs_.io_diffCommits_info_53_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_53_rfWen=0x%0h while the rhs_.io_diffCommits_info_53_rfWen=0x%0h",this.io_diffCommits_info_53_rfWen,rhs_.io_diffCommits_info_53_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_53_fpWen!=rhs_.io_diffCommits_info_53_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_53_fpWen=0x%0h while the rhs_.io_diffCommits_info_53_fpWen=0x%0h",this.io_diffCommits_info_53_fpWen,rhs_.io_diffCommits_info_53_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_53_vecWen!=rhs_.io_diffCommits_info_53_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_53_vecWen=0x%0h while the rhs_.io_diffCommits_info_53_vecWen=0x%0h",this.io_diffCommits_info_53_vecWen,rhs_.io_diffCommits_info_53_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_53_v0Wen!=rhs_.io_diffCommits_info_53_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_53_v0Wen=0x%0h while the rhs_.io_diffCommits_info_53_v0Wen=0x%0h",this.io_diffCommits_info_53_v0Wen,rhs_.io_diffCommits_info_53_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_53_vlWen!=rhs_.io_diffCommits_info_53_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_53_vlWen=0x%0h while the rhs_.io_diffCommits_info_53_vlWen=0x%0h",this.io_diffCommits_info_53_vlWen,rhs_.io_diffCommits_info_53_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_54_ldest!=rhs_.io_diffCommits_info_54_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_54_ldest=0x%0h while the rhs_.io_diffCommits_info_54_ldest=0x%0h",this.io_diffCommits_info_54_ldest,rhs_.io_diffCommits_info_54_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_54_pdest!=rhs_.io_diffCommits_info_54_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_54_pdest=0x%0h while the rhs_.io_diffCommits_info_54_pdest=0x%0h",this.io_diffCommits_info_54_pdest,rhs_.io_diffCommits_info_54_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_54_rfWen!=rhs_.io_diffCommits_info_54_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_54_rfWen=0x%0h while the rhs_.io_diffCommits_info_54_rfWen=0x%0h",this.io_diffCommits_info_54_rfWen,rhs_.io_diffCommits_info_54_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_54_fpWen!=rhs_.io_diffCommits_info_54_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_54_fpWen=0x%0h while the rhs_.io_diffCommits_info_54_fpWen=0x%0h",this.io_diffCommits_info_54_fpWen,rhs_.io_diffCommits_info_54_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_54_vecWen!=rhs_.io_diffCommits_info_54_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_54_vecWen=0x%0h while the rhs_.io_diffCommits_info_54_vecWen=0x%0h",this.io_diffCommits_info_54_vecWen,rhs_.io_diffCommits_info_54_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_54_v0Wen!=rhs_.io_diffCommits_info_54_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_54_v0Wen=0x%0h while the rhs_.io_diffCommits_info_54_v0Wen=0x%0h",this.io_diffCommits_info_54_v0Wen,rhs_.io_diffCommits_info_54_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_54_vlWen!=rhs_.io_diffCommits_info_54_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_54_vlWen=0x%0h while the rhs_.io_diffCommits_info_54_vlWen=0x%0h",this.io_diffCommits_info_54_vlWen,rhs_.io_diffCommits_info_54_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_55_ldest!=rhs_.io_diffCommits_info_55_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_55_ldest=0x%0h while the rhs_.io_diffCommits_info_55_ldest=0x%0h",this.io_diffCommits_info_55_ldest,rhs_.io_diffCommits_info_55_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_55_pdest!=rhs_.io_diffCommits_info_55_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_55_pdest=0x%0h while the rhs_.io_diffCommits_info_55_pdest=0x%0h",this.io_diffCommits_info_55_pdest,rhs_.io_diffCommits_info_55_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_55_rfWen!=rhs_.io_diffCommits_info_55_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_55_rfWen=0x%0h while the rhs_.io_diffCommits_info_55_rfWen=0x%0h",this.io_diffCommits_info_55_rfWen,rhs_.io_diffCommits_info_55_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_55_fpWen!=rhs_.io_diffCommits_info_55_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_55_fpWen=0x%0h while the rhs_.io_diffCommits_info_55_fpWen=0x%0h",this.io_diffCommits_info_55_fpWen,rhs_.io_diffCommits_info_55_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_55_vecWen!=rhs_.io_diffCommits_info_55_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_55_vecWen=0x%0h while the rhs_.io_diffCommits_info_55_vecWen=0x%0h",this.io_diffCommits_info_55_vecWen,rhs_.io_diffCommits_info_55_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_55_v0Wen!=rhs_.io_diffCommits_info_55_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_55_v0Wen=0x%0h while the rhs_.io_diffCommits_info_55_v0Wen=0x%0h",this.io_diffCommits_info_55_v0Wen,rhs_.io_diffCommits_info_55_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_55_vlWen!=rhs_.io_diffCommits_info_55_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_55_vlWen=0x%0h while the rhs_.io_diffCommits_info_55_vlWen=0x%0h",this.io_diffCommits_info_55_vlWen,rhs_.io_diffCommits_info_55_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_56_ldest!=rhs_.io_diffCommits_info_56_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_56_ldest=0x%0h while the rhs_.io_diffCommits_info_56_ldest=0x%0h",this.io_diffCommits_info_56_ldest,rhs_.io_diffCommits_info_56_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_56_pdest!=rhs_.io_diffCommits_info_56_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_56_pdest=0x%0h while the rhs_.io_diffCommits_info_56_pdest=0x%0h",this.io_diffCommits_info_56_pdest,rhs_.io_diffCommits_info_56_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_56_rfWen!=rhs_.io_diffCommits_info_56_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_56_rfWen=0x%0h while the rhs_.io_diffCommits_info_56_rfWen=0x%0h",this.io_diffCommits_info_56_rfWen,rhs_.io_diffCommits_info_56_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_56_fpWen!=rhs_.io_diffCommits_info_56_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_56_fpWen=0x%0h while the rhs_.io_diffCommits_info_56_fpWen=0x%0h",this.io_diffCommits_info_56_fpWen,rhs_.io_diffCommits_info_56_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_56_vecWen!=rhs_.io_diffCommits_info_56_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_56_vecWen=0x%0h while the rhs_.io_diffCommits_info_56_vecWen=0x%0h",this.io_diffCommits_info_56_vecWen,rhs_.io_diffCommits_info_56_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_56_v0Wen!=rhs_.io_diffCommits_info_56_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_56_v0Wen=0x%0h while the rhs_.io_diffCommits_info_56_v0Wen=0x%0h",this.io_diffCommits_info_56_v0Wen,rhs_.io_diffCommits_info_56_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_56_vlWen!=rhs_.io_diffCommits_info_56_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_56_vlWen=0x%0h while the rhs_.io_diffCommits_info_56_vlWen=0x%0h",this.io_diffCommits_info_56_vlWen,rhs_.io_diffCommits_info_56_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_57_ldest!=rhs_.io_diffCommits_info_57_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_57_ldest=0x%0h while the rhs_.io_diffCommits_info_57_ldest=0x%0h",this.io_diffCommits_info_57_ldest,rhs_.io_diffCommits_info_57_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_57_pdest!=rhs_.io_diffCommits_info_57_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_57_pdest=0x%0h while the rhs_.io_diffCommits_info_57_pdest=0x%0h",this.io_diffCommits_info_57_pdest,rhs_.io_diffCommits_info_57_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_57_rfWen!=rhs_.io_diffCommits_info_57_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_57_rfWen=0x%0h while the rhs_.io_diffCommits_info_57_rfWen=0x%0h",this.io_diffCommits_info_57_rfWen,rhs_.io_diffCommits_info_57_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_57_fpWen!=rhs_.io_diffCommits_info_57_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_57_fpWen=0x%0h while the rhs_.io_diffCommits_info_57_fpWen=0x%0h",this.io_diffCommits_info_57_fpWen,rhs_.io_diffCommits_info_57_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_57_vecWen!=rhs_.io_diffCommits_info_57_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_57_vecWen=0x%0h while the rhs_.io_diffCommits_info_57_vecWen=0x%0h",this.io_diffCommits_info_57_vecWen,rhs_.io_diffCommits_info_57_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_57_v0Wen!=rhs_.io_diffCommits_info_57_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_57_v0Wen=0x%0h while the rhs_.io_diffCommits_info_57_v0Wen=0x%0h",this.io_diffCommits_info_57_v0Wen,rhs_.io_diffCommits_info_57_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_57_vlWen!=rhs_.io_diffCommits_info_57_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_57_vlWen=0x%0h while the rhs_.io_diffCommits_info_57_vlWen=0x%0h",this.io_diffCommits_info_57_vlWen,rhs_.io_diffCommits_info_57_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_58_ldest!=rhs_.io_diffCommits_info_58_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_58_ldest=0x%0h while the rhs_.io_diffCommits_info_58_ldest=0x%0h",this.io_diffCommits_info_58_ldest,rhs_.io_diffCommits_info_58_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_58_pdest!=rhs_.io_diffCommits_info_58_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_58_pdest=0x%0h while the rhs_.io_diffCommits_info_58_pdest=0x%0h",this.io_diffCommits_info_58_pdest,rhs_.io_diffCommits_info_58_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_58_rfWen!=rhs_.io_diffCommits_info_58_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_58_rfWen=0x%0h while the rhs_.io_diffCommits_info_58_rfWen=0x%0h",this.io_diffCommits_info_58_rfWen,rhs_.io_diffCommits_info_58_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_58_fpWen!=rhs_.io_diffCommits_info_58_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_58_fpWen=0x%0h while the rhs_.io_diffCommits_info_58_fpWen=0x%0h",this.io_diffCommits_info_58_fpWen,rhs_.io_diffCommits_info_58_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_58_vecWen!=rhs_.io_diffCommits_info_58_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_58_vecWen=0x%0h while the rhs_.io_diffCommits_info_58_vecWen=0x%0h",this.io_diffCommits_info_58_vecWen,rhs_.io_diffCommits_info_58_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_58_v0Wen!=rhs_.io_diffCommits_info_58_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_58_v0Wen=0x%0h while the rhs_.io_diffCommits_info_58_v0Wen=0x%0h",this.io_diffCommits_info_58_v0Wen,rhs_.io_diffCommits_info_58_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_58_vlWen!=rhs_.io_diffCommits_info_58_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_58_vlWen=0x%0h while the rhs_.io_diffCommits_info_58_vlWen=0x%0h",this.io_diffCommits_info_58_vlWen,rhs_.io_diffCommits_info_58_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_59_ldest!=rhs_.io_diffCommits_info_59_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_59_ldest=0x%0h while the rhs_.io_diffCommits_info_59_ldest=0x%0h",this.io_diffCommits_info_59_ldest,rhs_.io_diffCommits_info_59_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_59_pdest!=rhs_.io_diffCommits_info_59_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_59_pdest=0x%0h while the rhs_.io_diffCommits_info_59_pdest=0x%0h",this.io_diffCommits_info_59_pdest,rhs_.io_diffCommits_info_59_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_59_rfWen!=rhs_.io_diffCommits_info_59_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_59_rfWen=0x%0h while the rhs_.io_diffCommits_info_59_rfWen=0x%0h",this.io_diffCommits_info_59_rfWen,rhs_.io_diffCommits_info_59_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_59_fpWen!=rhs_.io_diffCommits_info_59_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_59_fpWen=0x%0h while the rhs_.io_diffCommits_info_59_fpWen=0x%0h",this.io_diffCommits_info_59_fpWen,rhs_.io_diffCommits_info_59_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_59_vecWen!=rhs_.io_diffCommits_info_59_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_59_vecWen=0x%0h while the rhs_.io_diffCommits_info_59_vecWen=0x%0h",this.io_diffCommits_info_59_vecWen,rhs_.io_diffCommits_info_59_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_59_v0Wen!=rhs_.io_diffCommits_info_59_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_59_v0Wen=0x%0h while the rhs_.io_diffCommits_info_59_v0Wen=0x%0h",this.io_diffCommits_info_59_v0Wen,rhs_.io_diffCommits_info_59_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_59_vlWen!=rhs_.io_diffCommits_info_59_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_59_vlWen=0x%0h while the rhs_.io_diffCommits_info_59_vlWen=0x%0h",this.io_diffCommits_info_59_vlWen,rhs_.io_diffCommits_info_59_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_60_ldest!=rhs_.io_diffCommits_info_60_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_60_ldest=0x%0h while the rhs_.io_diffCommits_info_60_ldest=0x%0h",this.io_diffCommits_info_60_ldest,rhs_.io_diffCommits_info_60_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_60_pdest!=rhs_.io_diffCommits_info_60_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_60_pdest=0x%0h while the rhs_.io_diffCommits_info_60_pdest=0x%0h",this.io_diffCommits_info_60_pdest,rhs_.io_diffCommits_info_60_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_60_rfWen!=rhs_.io_diffCommits_info_60_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_60_rfWen=0x%0h while the rhs_.io_diffCommits_info_60_rfWen=0x%0h",this.io_diffCommits_info_60_rfWen,rhs_.io_diffCommits_info_60_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_60_fpWen!=rhs_.io_diffCommits_info_60_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_60_fpWen=0x%0h while the rhs_.io_diffCommits_info_60_fpWen=0x%0h",this.io_diffCommits_info_60_fpWen,rhs_.io_diffCommits_info_60_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_60_vecWen!=rhs_.io_diffCommits_info_60_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_60_vecWen=0x%0h while the rhs_.io_diffCommits_info_60_vecWen=0x%0h",this.io_diffCommits_info_60_vecWen,rhs_.io_diffCommits_info_60_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_60_v0Wen!=rhs_.io_diffCommits_info_60_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_60_v0Wen=0x%0h while the rhs_.io_diffCommits_info_60_v0Wen=0x%0h",this.io_diffCommits_info_60_v0Wen,rhs_.io_diffCommits_info_60_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_60_vlWen!=rhs_.io_diffCommits_info_60_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_60_vlWen=0x%0h while the rhs_.io_diffCommits_info_60_vlWen=0x%0h",this.io_diffCommits_info_60_vlWen,rhs_.io_diffCommits_info_60_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_61_ldest!=rhs_.io_diffCommits_info_61_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_61_ldest=0x%0h while the rhs_.io_diffCommits_info_61_ldest=0x%0h",this.io_diffCommits_info_61_ldest,rhs_.io_diffCommits_info_61_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_61_pdest!=rhs_.io_diffCommits_info_61_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_61_pdest=0x%0h while the rhs_.io_diffCommits_info_61_pdest=0x%0h",this.io_diffCommits_info_61_pdest,rhs_.io_diffCommits_info_61_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_61_rfWen!=rhs_.io_diffCommits_info_61_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_61_rfWen=0x%0h while the rhs_.io_diffCommits_info_61_rfWen=0x%0h",this.io_diffCommits_info_61_rfWen,rhs_.io_diffCommits_info_61_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_61_fpWen!=rhs_.io_diffCommits_info_61_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_61_fpWen=0x%0h while the rhs_.io_diffCommits_info_61_fpWen=0x%0h",this.io_diffCommits_info_61_fpWen,rhs_.io_diffCommits_info_61_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_61_vecWen!=rhs_.io_diffCommits_info_61_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_61_vecWen=0x%0h while the rhs_.io_diffCommits_info_61_vecWen=0x%0h",this.io_diffCommits_info_61_vecWen,rhs_.io_diffCommits_info_61_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_61_v0Wen!=rhs_.io_diffCommits_info_61_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_61_v0Wen=0x%0h while the rhs_.io_diffCommits_info_61_v0Wen=0x%0h",this.io_diffCommits_info_61_v0Wen,rhs_.io_diffCommits_info_61_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_61_vlWen!=rhs_.io_diffCommits_info_61_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_61_vlWen=0x%0h while the rhs_.io_diffCommits_info_61_vlWen=0x%0h",this.io_diffCommits_info_61_vlWen,rhs_.io_diffCommits_info_61_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_62_ldest!=rhs_.io_diffCommits_info_62_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_62_ldest=0x%0h while the rhs_.io_diffCommits_info_62_ldest=0x%0h",this.io_diffCommits_info_62_ldest,rhs_.io_diffCommits_info_62_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_62_pdest!=rhs_.io_diffCommits_info_62_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_62_pdest=0x%0h while the rhs_.io_diffCommits_info_62_pdest=0x%0h",this.io_diffCommits_info_62_pdest,rhs_.io_diffCommits_info_62_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_62_rfWen!=rhs_.io_diffCommits_info_62_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_62_rfWen=0x%0h while the rhs_.io_diffCommits_info_62_rfWen=0x%0h",this.io_diffCommits_info_62_rfWen,rhs_.io_diffCommits_info_62_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_62_fpWen!=rhs_.io_diffCommits_info_62_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_62_fpWen=0x%0h while the rhs_.io_diffCommits_info_62_fpWen=0x%0h",this.io_diffCommits_info_62_fpWen,rhs_.io_diffCommits_info_62_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_62_vecWen!=rhs_.io_diffCommits_info_62_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_62_vecWen=0x%0h while the rhs_.io_diffCommits_info_62_vecWen=0x%0h",this.io_diffCommits_info_62_vecWen,rhs_.io_diffCommits_info_62_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_62_v0Wen!=rhs_.io_diffCommits_info_62_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_62_v0Wen=0x%0h while the rhs_.io_diffCommits_info_62_v0Wen=0x%0h",this.io_diffCommits_info_62_v0Wen,rhs_.io_diffCommits_info_62_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_62_vlWen!=rhs_.io_diffCommits_info_62_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_62_vlWen=0x%0h while the rhs_.io_diffCommits_info_62_vlWen=0x%0h",this.io_diffCommits_info_62_vlWen,rhs_.io_diffCommits_info_62_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_63_ldest!=rhs_.io_diffCommits_info_63_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_63_ldest=0x%0h while the rhs_.io_diffCommits_info_63_ldest=0x%0h",this.io_diffCommits_info_63_ldest,rhs_.io_diffCommits_info_63_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_63_pdest!=rhs_.io_diffCommits_info_63_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_63_pdest=0x%0h while the rhs_.io_diffCommits_info_63_pdest=0x%0h",this.io_diffCommits_info_63_pdest,rhs_.io_diffCommits_info_63_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_63_rfWen!=rhs_.io_diffCommits_info_63_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_63_rfWen=0x%0h while the rhs_.io_diffCommits_info_63_rfWen=0x%0h",this.io_diffCommits_info_63_rfWen,rhs_.io_diffCommits_info_63_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_63_fpWen!=rhs_.io_diffCommits_info_63_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_63_fpWen=0x%0h while the rhs_.io_diffCommits_info_63_fpWen=0x%0h",this.io_diffCommits_info_63_fpWen,rhs_.io_diffCommits_info_63_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_63_vecWen!=rhs_.io_diffCommits_info_63_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_63_vecWen=0x%0h while the rhs_.io_diffCommits_info_63_vecWen=0x%0h",this.io_diffCommits_info_63_vecWen,rhs_.io_diffCommits_info_63_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_63_v0Wen!=rhs_.io_diffCommits_info_63_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_63_v0Wen=0x%0h while the rhs_.io_diffCommits_info_63_v0Wen=0x%0h",this.io_diffCommits_info_63_v0Wen,rhs_.io_diffCommits_info_63_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_63_vlWen!=rhs_.io_diffCommits_info_63_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_63_vlWen=0x%0h while the rhs_.io_diffCommits_info_63_vlWen=0x%0h",this.io_diffCommits_info_63_vlWen,rhs_.io_diffCommits_info_63_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_64_ldest!=rhs_.io_diffCommits_info_64_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_64_ldest=0x%0h while the rhs_.io_diffCommits_info_64_ldest=0x%0h",this.io_diffCommits_info_64_ldest,rhs_.io_diffCommits_info_64_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_64_pdest!=rhs_.io_diffCommits_info_64_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_64_pdest=0x%0h while the rhs_.io_diffCommits_info_64_pdest=0x%0h",this.io_diffCommits_info_64_pdest,rhs_.io_diffCommits_info_64_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_64_rfWen!=rhs_.io_diffCommits_info_64_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_64_rfWen=0x%0h while the rhs_.io_diffCommits_info_64_rfWen=0x%0h",this.io_diffCommits_info_64_rfWen,rhs_.io_diffCommits_info_64_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_64_fpWen!=rhs_.io_diffCommits_info_64_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_64_fpWen=0x%0h while the rhs_.io_diffCommits_info_64_fpWen=0x%0h",this.io_diffCommits_info_64_fpWen,rhs_.io_diffCommits_info_64_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_64_vecWen!=rhs_.io_diffCommits_info_64_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_64_vecWen=0x%0h while the rhs_.io_diffCommits_info_64_vecWen=0x%0h",this.io_diffCommits_info_64_vecWen,rhs_.io_diffCommits_info_64_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_64_v0Wen!=rhs_.io_diffCommits_info_64_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_64_v0Wen=0x%0h while the rhs_.io_diffCommits_info_64_v0Wen=0x%0h",this.io_diffCommits_info_64_v0Wen,rhs_.io_diffCommits_info_64_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_64_vlWen!=rhs_.io_diffCommits_info_64_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_64_vlWen=0x%0h while the rhs_.io_diffCommits_info_64_vlWen=0x%0h",this.io_diffCommits_info_64_vlWen,rhs_.io_diffCommits_info_64_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_65_ldest!=rhs_.io_diffCommits_info_65_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_65_ldest=0x%0h while the rhs_.io_diffCommits_info_65_ldest=0x%0h",this.io_diffCommits_info_65_ldest,rhs_.io_diffCommits_info_65_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_65_pdest!=rhs_.io_diffCommits_info_65_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_65_pdest=0x%0h while the rhs_.io_diffCommits_info_65_pdest=0x%0h",this.io_diffCommits_info_65_pdest,rhs_.io_diffCommits_info_65_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_65_rfWen!=rhs_.io_diffCommits_info_65_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_65_rfWen=0x%0h while the rhs_.io_diffCommits_info_65_rfWen=0x%0h",this.io_diffCommits_info_65_rfWen,rhs_.io_diffCommits_info_65_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_65_fpWen!=rhs_.io_diffCommits_info_65_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_65_fpWen=0x%0h while the rhs_.io_diffCommits_info_65_fpWen=0x%0h",this.io_diffCommits_info_65_fpWen,rhs_.io_diffCommits_info_65_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_65_vecWen!=rhs_.io_diffCommits_info_65_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_65_vecWen=0x%0h while the rhs_.io_diffCommits_info_65_vecWen=0x%0h",this.io_diffCommits_info_65_vecWen,rhs_.io_diffCommits_info_65_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_65_v0Wen!=rhs_.io_diffCommits_info_65_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_65_v0Wen=0x%0h while the rhs_.io_diffCommits_info_65_v0Wen=0x%0h",this.io_diffCommits_info_65_v0Wen,rhs_.io_diffCommits_info_65_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_65_vlWen!=rhs_.io_diffCommits_info_65_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_65_vlWen=0x%0h while the rhs_.io_diffCommits_info_65_vlWen=0x%0h",this.io_diffCommits_info_65_vlWen,rhs_.io_diffCommits_info_65_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_66_ldest!=rhs_.io_diffCommits_info_66_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_66_ldest=0x%0h while the rhs_.io_diffCommits_info_66_ldest=0x%0h",this.io_diffCommits_info_66_ldest,rhs_.io_diffCommits_info_66_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_66_pdest!=rhs_.io_diffCommits_info_66_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_66_pdest=0x%0h while the rhs_.io_diffCommits_info_66_pdest=0x%0h",this.io_diffCommits_info_66_pdest,rhs_.io_diffCommits_info_66_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_66_rfWen!=rhs_.io_diffCommits_info_66_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_66_rfWen=0x%0h while the rhs_.io_diffCommits_info_66_rfWen=0x%0h",this.io_diffCommits_info_66_rfWen,rhs_.io_diffCommits_info_66_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_66_fpWen!=rhs_.io_diffCommits_info_66_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_66_fpWen=0x%0h while the rhs_.io_diffCommits_info_66_fpWen=0x%0h",this.io_diffCommits_info_66_fpWen,rhs_.io_diffCommits_info_66_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_66_vecWen!=rhs_.io_diffCommits_info_66_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_66_vecWen=0x%0h while the rhs_.io_diffCommits_info_66_vecWen=0x%0h",this.io_diffCommits_info_66_vecWen,rhs_.io_diffCommits_info_66_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_66_v0Wen!=rhs_.io_diffCommits_info_66_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_66_v0Wen=0x%0h while the rhs_.io_diffCommits_info_66_v0Wen=0x%0h",this.io_diffCommits_info_66_v0Wen,rhs_.io_diffCommits_info_66_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_66_vlWen!=rhs_.io_diffCommits_info_66_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_66_vlWen=0x%0h while the rhs_.io_diffCommits_info_66_vlWen=0x%0h",this.io_diffCommits_info_66_vlWen,rhs_.io_diffCommits_info_66_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_67_ldest!=rhs_.io_diffCommits_info_67_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_67_ldest=0x%0h while the rhs_.io_diffCommits_info_67_ldest=0x%0h",this.io_diffCommits_info_67_ldest,rhs_.io_diffCommits_info_67_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_67_pdest!=rhs_.io_diffCommits_info_67_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_67_pdest=0x%0h while the rhs_.io_diffCommits_info_67_pdest=0x%0h",this.io_diffCommits_info_67_pdest,rhs_.io_diffCommits_info_67_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_67_rfWen!=rhs_.io_diffCommits_info_67_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_67_rfWen=0x%0h while the rhs_.io_diffCommits_info_67_rfWen=0x%0h",this.io_diffCommits_info_67_rfWen,rhs_.io_diffCommits_info_67_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_67_fpWen!=rhs_.io_diffCommits_info_67_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_67_fpWen=0x%0h while the rhs_.io_diffCommits_info_67_fpWen=0x%0h",this.io_diffCommits_info_67_fpWen,rhs_.io_diffCommits_info_67_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_67_vecWen!=rhs_.io_diffCommits_info_67_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_67_vecWen=0x%0h while the rhs_.io_diffCommits_info_67_vecWen=0x%0h",this.io_diffCommits_info_67_vecWen,rhs_.io_diffCommits_info_67_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_67_v0Wen!=rhs_.io_diffCommits_info_67_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_67_v0Wen=0x%0h while the rhs_.io_diffCommits_info_67_v0Wen=0x%0h",this.io_diffCommits_info_67_v0Wen,rhs_.io_diffCommits_info_67_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_67_vlWen!=rhs_.io_diffCommits_info_67_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_67_vlWen=0x%0h while the rhs_.io_diffCommits_info_67_vlWen=0x%0h",this.io_diffCommits_info_67_vlWen,rhs_.io_diffCommits_info_67_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_68_ldest!=rhs_.io_diffCommits_info_68_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_68_ldest=0x%0h while the rhs_.io_diffCommits_info_68_ldest=0x%0h",this.io_diffCommits_info_68_ldest,rhs_.io_diffCommits_info_68_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_68_pdest!=rhs_.io_diffCommits_info_68_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_68_pdest=0x%0h while the rhs_.io_diffCommits_info_68_pdest=0x%0h",this.io_diffCommits_info_68_pdest,rhs_.io_diffCommits_info_68_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_68_rfWen!=rhs_.io_diffCommits_info_68_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_68_rfWen=0x%0h while the rhs_.io_diffCommits_info_68_rfWen=0x%0h",this.io_diffCommits_info_68_rfWen,rhs_.io_diffCommits_info_68_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_68_fpWen!=rhs_.io_diffCommits_info_68_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_68_fpWen=0x%0h while the rhs_.io_diffCommits_info_68_fpWen=0x%0h",this.io_diffCommits_info_68_fpWen,rhs_.io_diffCommits_info_68_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_68_vecWen!=rhs_.io_diffCommits_info_68_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_68_vecWen=0x%0h while the rhs_.io_diffCommits_info_68_vecWen=0x%0h",this.io_diffCommits_info_68_vecWen,rhs_.io_diffCommits_info_68_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_68_v0Wen!=rhs_.io_diffCommits_info_68_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_68_v0Wen=0x%0h while the rhs_.io_diffCommits_info_68_v0Wen=0x%0h",this.io_diffCommits_info_68_v0Wen,rhs_.io_diffCommits_info_68_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_68_vlWen!=rhs_.io_diffCommits_info_68_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_68_vlWen=0x%0h while the rhs_.io_diffCommits_info_68_vlWen=0x%0h",this.io_diffCommits_info_68_vlWen,rhs_.io_diffCommits_info_68_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_69_ldest!=rhs_.io_diffCommits_info_69_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_69_ldest=0x%0h while the rhs_.io_diffCommits_info_69_ldest=0x%0h",this.io_diffCommits_info_69_ldest,rhs_.io_diffCommits_info_69_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_69_pdest!=rhs_.io_diffCommits_info_69_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_69_pdest=0x%0h while the rhs_.io_diffCommits_info_69_pdest=0x%0h",this.io_diffCommits_info_69_pdest,rhs_.io_diffCommits_info_69_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_69_rfWen!=rhs_.io_diffCommits_info_69_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_69_rfWen=0x%0h while the rhs_.io_diffCommits_info_69_rfWen=0x%0h",this.io_diffCommits_info_69_rfWen,rhs_.io_diffCommits_info_69_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_69_fpWen!=rhs_.io_diffCommits_info_69_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_69_fpWen=0x%0h while the rhs_.io_diffCommits_info_69_fpWen=0x%0h",this.io_diffCommits_info_69_fpWen,rhs_.io_diffCommits_info_69_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_69_vecWen!=rhs_.io_diffCommits_info_69_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_69_vecWen=0x%0h while the rhs_.io_diffCommits_info_69_vecWen=0x%0h",this.io_diffCommits_info_69_vecWen,rhs_.io_diffCommits_info_69_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_69_v0Wen!=rhs_.io_diffCommits_info_69_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_69_v0Wen=0x%0h while the rhs_.io_diffCommits_info_69_v0Wen=0x%0h",this.io_diffCommits_info_69_v0Wen,rhs_.io_diffCommits_info_69_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_69_vlWen!=rhs_.io_diffCommits_info_69_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_69_vlWen=0x%0h while the rhs_.io_diffCommits_info_69_vlWen=0x%0h",this.io_diffCommits_info_69_vlWen,rhs_.io_diffCommits_info_69_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_70_ldest!=rhs_.io_diffCommits_info_70_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_70_ldest=0x%0h while the rhs_.io_diffCommits_info_70_ldest=0x%0h",this.io_diffCommits_info_70_ldest,rhs_.io_diffCommits_info_70_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_70_pdest!=rhs_.io_diffCommits_info_70_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_70_pdest=0x%0h while the rhs_.io_diffCommits_info_70_pdest=0x%0h",this.io_diffCommits_info_70_pdest,rhs_.io_diffCommits_info_70_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_70_rfWen!=rhs_.io_diffCommits_info_70_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_70_rfWen=0x%0h while the rhs_.io_diffCommits_info_70_rfWen=0x%0h",this.io_diffCommits_info_70_rfWen,rhs_.io_diffCommits_info_70_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_70_fpWen!=rhs_.io_diffCommits_info_70_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_70_fpWen=0x%0h while the rhs_.io_diffCommits_info_70_fpWen=0x%0h",this.io_diffCommits_info_70_fpWen,rhs_.io_diffCommits_info_70_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_70_vecWen!=rhs_.io_diffCommits_info_70_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_70_vecWen=0x%0h while the rhs_.io_diffCommits_info_70_vecWen=0x%0h",this.io_diffCommits_info_70_vecWen,rhs_.io_diffCommits_info_70_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_70_v0Wen!=rhs_.io_diffCommits_info_70_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_70_v0Wen=0x%0h while the rhs_.io_diffCommits_info_70_v0Wen=0x%0h",this.io_diffCommits_info_70_v0Wen,rhs_.io_diffCommits_info_70_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_70_vlWen!=rhs_.io_diffCommits_info_70_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_70_vlWen=0x%0h while the rhs_.io_diffCommits_info_70_vlWen=0x%0h",this.io_diffCommits_info_70_vlWen,rhs_.io_diffCommits_info_70_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_71_ldest!=rhs_.io_diffCommits_info_71_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_71_ldest=0x%0h while the rhs_.io_diffCommits_info_71_ldest=0x%0h",this.io_diffCommits_info_71_ldest,rhs_.io_diffCommits_info_71_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_71_pdest!=rhs_.io_diffCommits_info_71_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_71_pdest=0x%0h while the rhs_.io_diffCommits_info_71_pdest=0x%0h",this.io_diffCommits_info_71_pdest,rhs_.io_diffCommits_info_71_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_71_rfWen!=rhs_.io_diffCommits_info_71_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_71_rfWen=0x%0h while the rhs_.io_diffCommits_info_71_rfWen=0x%0h",this.io_diffCommits_info_71_rfWen,rhs_.io_diffCommits_info_71_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_71_fpWen!=rhs_.io_diffCommits_info_71_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_71_fpWen=0x%0h while the rhs_.io_diffCommits_info_71_fpWen=0x%0h",this.io_diffCommits_info_71_fpWen,rhs_.io_diffCommits_info_71_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_71_vecWen!=rhs_.io_diffCommits_info_71_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_71_vecWen=0x%0h while the rhs_.io_diffCommits_info_71_vecWen=0x%0h",this.io_diffCommits_info_71_vecWen,rhs_.io_diffCommits_info_71_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_71_v0Wen!=rhs_.io_diffCommits_info_71_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_71_v0Wen=0x%0h while the rhs_.io_diffCommits_info_71_v0Wen=0x%0h",this.io_diffCommits_info_71_v0Wen,rhs_.io_diffCommits_info_71_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_71_vlWen!=rhs_.io_diffCommits_info_71_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_71_vlWen=0x%0h while the rhs_.io_diffCommits_info_71_vlWen=0x%0h",this.io_diffCommits_info_71_vlWen,rhs_.io_diffCommits_info_71_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_72_ldest!=rhs_.io_diffCommits_info_72_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_72_ldest=0x%0h while the rhs_.io_diffCommits_info_72_ldest=0x%0h",this.io_diffCommits_info_72_ldest,rhs_.io_diffCommits_info_72_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_72_pdest!=rhs_.io_diffCommits_info_72_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_72_pdest=0x%0h while the rhs_.io_diffCommits_info_72_pdest=0x%0h",this.io_diffCommits_info_72_pdest,rhs_.io_diffCommits_info_72_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_72_rfWen!=rhs_.io_diffCommits_info_72_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_72_rfWen=0x%0h while the rhs_.io_diffCommits_info_72_rfWen=0x%0h",this.io_diffCommits_info_72_rfWen,rhs_.io_diffCommits_info_72_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_72_fpWen!=rhs_.io_diffCommits_info_72_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_72_fpWen=0x%0h while the rhs_.io_diffCommits_info_72_fpWen=0x%0h",this.io_diffCommits_info_72_fpWen,rhs_.io_diffCommits_info_72_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_72_vecWen!=rhs_.io_diffCommits_info_72_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_72_vecWen=0x%0h while the rhs_.io_diffCommits_info_72_vecWen=0x%0h",this.io_diffCommits_info_72_vecWen,rhs_.io_diffCommits_info_72_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_72_v0Wen!=rhs_.io_diffCommits_info_72_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_72_v0Wen=0x%0h while the rhs_.io_diffCommits_info_72_v0Wen=0x%0h",this.io_diffCommits_info_72_v0Wen,rhs_.io_diffCommits_info_72_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_72_vlWen!=rhs_.io_diffCommits_info_72_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_72_vlWen=0x%0h while the rhs_.io_diffCommits_info_72_vlWen=0x%0h",this.io_diffCommits_info_72_vlWen,rhs_.io_diffCommits_info_72_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_73_ldest!=rhs_.io_diffCommits_info_73_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_73_ldest=0x%0h while the rhs_.io_diffCommits_info_73_ldest=0x%0h",this.io_diffCommits_info_73_ldest,rhs_.io_diffCommits_info_73_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_73_pdest!=rhs_.io_diffCommits_info_73_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_73_pdest=0x%0h while the rhs_.io_diffCommits_info_73_pdest=0x%0h",this.io_diffCommits_info_73_pdest,rhs_.io_diffCommits_info_73_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_73_rfWen!=rhs_.io_diffCommits_info_73_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_73_rfWen=0x%0h while the rhs_.io_diffCommits_info_73_rfWen=0x%0h",this.io_diffCommits_info_73_rfWen,rhs_.io_diffCommits_info_73_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_73_fpWen!=rhs_.io_diffCommits_info_73_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_73_fpWen=0x%0h while the rhs_.io_diffCommits_info_73_fpWen=0x%0h",this.io_diffCommits_info_73_fpWen,rhs_.io_diffCommits_info_73_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_73_vecWen!=rhs_.io_diffCommits_info_73_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_73_vecWen=0x%0h while the rhs_.io_diffCommits_info_73_vecWen=0x%0h",this.io_diffCommits_info_73_vecWen,rhs_.io_diffCommits_info_73_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_73_v0Wen!=rhs_.io_diffCommits_info_73_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_73_v0Wen=0x%0h while the rhs_.io_diffCommits_info_73_v0Wen=0x%0h",this.io_diffCommits_info_73_v0Wen,rhs_.io_diffCommits_info_73_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_73_vlWen!=rhs_.io_diffCommits_info_73_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_73_vlWen=0x%0h while the rhs_.io_diffCommits_info_73_vlWen=0x%0h",this.io_diffCommits_info_73_vlWen,rhs_.io_diffCommits_info_73_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_74_ldest!=rhs_.io_diffCommits_info_74_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_74_ldest=0x%0h while the rhs_.io_diffCommits_info_74_ldest=0x%0h",this.io_diffCommits_info_74_ldest,rhs_.io_diffCommits_info_74_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_74_pdest!=rhs_.io_diffCommits_info_74_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_74_pdest=0x%0h while the rhs_.io_diffCommits_info_74_pdest=0x%0h",this.io_diffCommits_info_74_pdest,rhs_.io_diffCommits_info_74_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_74_rfWen!=rhs_.io_diffCommits_info_74_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_74_rfWen=0x%0h while the rhs_.io_diffCommits_info_74_rfWen=0x%0h",this.io_diffCommits_info_74_rfWen,rhs_.io_diffCommits_info_74_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_74_fpWen!=rhs_.io_diffCommits_info_74_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_74_fpWen=0x%0h while the rhs_.io_diffCommits_info_74_fpWen=0x%0h",this.io_diffCommits_info_74_fpWen,rhs_.io_diffCommits_info_74_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_74_vecWen!=rhs_.io_diffCommits_info_74_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_74_vecWen=0x%0h while the rhs_.io_diffCommits_info_74_vecWen=0x%0h",this.io_diffCommits_info_74_vecWen,rhs_.io_diffCommits_info_74_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_74_v0Wen!=rhs_.io_diffCommits_info_74_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_74_v0Wen=0x%0h while the rhs_.io_diffCommits_info_74_v0Wen=0x%0h",this.io_diffCommits_info_74_v0Wen,rhs_.io_diffCommits_info_74_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_74_vlWen!=rhs_.io_diffCommits_info_74_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_74_vlWen=0x%0h while the rhs_.io_diffCommits_info_74_vlWen=0x%0h",this.io_diffCommits_info_74_vlWen,rhs_.io_diffCommits_info_74_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_75_ldest!=rhs_.io_diffCommits_info_75_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_75_ldest=0x%0h while the rhs_.io_diffCommits_info_75_ldest=0x%0h",this.io_diffCommits_info_75_ldest,rhs_.io_diffCommits_info_75_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_75_pdest!=rhs_.io_diffCommits_info_75_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_75_pdest=0x%0h while the rhs_.io_diffCommits_info_75_pdest=0x%0h",this.io_diffCommits_info_75_pdest,rhs_.io_diffCommits_info_75_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_75_rfWen!=rhs_.io_diffCommits_info_75_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_75_rfWen=0x%0h while the rhs_.io_diffCommits_info_75_rfWen=0x%0h",this.io_diffCommits_info_75_rfWen,rhs_.io_diffCommits_info_75_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_75_fpWen!=rhs_.io_diffCommits_info_75_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_75_fpWen=0x%0h while the rhs_.io_diffCommits_info_75_fpWen=0x%0h",this.io_diffCommits_info_75_fpWen,rhs_.io_diffCommits_info_75_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_75_vecWen!=rhs_.io_diffCommits_info_75_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_75_vecWen=0x%0h while the rhs_.io_diffCommits_info_75_vecWen=0x%0h",this.io_diffCommits_info_75_vecWen,rhs_.io_diffCommits_info_75_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_75_v0Wen!=rhs_.io_diffCommits_info_75_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_75_v0Wen=0x%0h while the rhs_.io_diffCommits_info_75_v0Wen=0x%0h",this.io_diffCommits_info_75_v0Wen,rhs_.io_diffCommits_info_75_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_75_vlWen!=rhs_.io_diffCommits_info_75_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_75_vlWen=0x%0h while the rhs_.io_diffCommits_info_75_vlWen=0x%0h",this.io_diffCommits_info_75_vlWen,rhs_.io_diffCommits_info_75_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_76_ldest!=rhs_.io_diffCommits_info_76_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_76_ldest=0x%0h while the rhs_.io_diffCommits_info_76_ldest=0x%0h",this.io_diffCommits_info_76_ldest,rhs_.io_diffCommits_info_76_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_76_pdest!=rhs_.io_diffCommits_info_76_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_76_pdest=0x%0h while the rhs_.io_diffCommits_info_76_pdest=0x%0h",this.io_diffCommits_info_76_pdest,rhs_.io_diffCommits_info_76_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_76_rfWen!=rhs_.io_diffCommits_info_76_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_76_rfWen=0x%0h while the rhs_.io_diffCommits_info_76_rfWen=0x%0h",this.io_diffCommits_info_76_rfWen,rhs_.io_diffCommits_info_76_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_76_fpWen!=rhs_.io_diffCommits_info_76_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_76_fpWen=0x%0h while the rhs_.io_diffCommits_info_76_fpWen=0x%0h",this.io_diffCommits_info_76_fpWen,rhs_.io_diffCommits_info_76_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_76_vecWen!=rhs_.io_diffCommits_info_76_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_76_vecWen=0x%0h while the rhs_.io_diffCommits_info_76_vecWen=0x%0h",this.io_diffCommits_info_76_vecWen,rhs_.io_diffCommits_info_76_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_76_v0Wen!=rhs_.io_diffCommits_info_76_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_76_v0Wen=0x%0h while the rhs_.io_diffCommits_info_76_v0Wen=0x%0h",this.io_diffCommits_info_76_v0Wen,rhs_.io_diffCommits_info_76_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_76_vlWen!=rhs_.io_diffCommits_info_76_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_76_vlWen=0x%0h while the rhs_.io_diffCommits_info_76_vlWen=0x%0h",this.io_diffCommits_info_76_vlWen,rhs_.io_diffCommits_info_76_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_77_ldest!=rhs_.io_diffCommits_info_77_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_77_ldest=0x%0h while the rhs_.io_diffCommits_info_77_ldest=0x%0h",this.io_diffCommits_info_77_ldest,rhs_.io_diffCommits_info_77_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_77_pdest!=rhs_.io_diffCommits_info_77_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_77_pdest=0x%0h while the rhs_.io_diffCommits_info_77_pdest=0x%0h",this.io_diffCommits_info_77_pdest,rhs_.io_diffCommits_info_77_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_77_rfWen!=rhs_.io_diffCommits_info_77_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_77_rfWen=0x%0h while the rhs_.io_diffCommits_info_77_rfWen=0x%0h",this.io_diffCommits_info_77_rfWen,rhs_.io_diffCommits_info_77_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_77_fpWen!=rhs_.io_diffCommits_info_77_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_77_fpWen=0x%0h while the rhs_.io_diffCommits_info_77_fpWen=0x%0h",this.io_diffCommits_info_77_fpWen,rhs_.io_diffCommits_info_77_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_77_vecWen!=rhs_.io_diffCommits_info_77_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_77_vecWen=0x%0h while the rhs_.io_diffCommits_info_77_vecWen=0x%0h",this.io_diffCommits_info_77_vecWen,rhs_.io_diffCommits_info_77_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_77_v0Wen!=rhs_.io_diffCommits_info_77_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_77_v0Wen=0x%0h while the rhs_.io_diffCommits_info_77_v0Wen=0x%0h",this.io_diffCommits_info_77_v0Wen,rhs_.io_diffCommits_info_77_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_77_vlWen!=rhs_.io_diffCommits_info_77_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_77_vlWen=0x%0h while the rhs_.io_diffCommits_info_77_vlWen=0x%0h",this.io_diffCommits_info_77_vlWen,rhs_.io_diffCommits_info_77_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_78_ldest!=rhs_.io_diffCommits_info_78_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_78_ldest=0x%0h while the rhs_.io_diffCommits_info_78_ldest=0x%0h",this.io_diffCommits_info_78_ldest,rhs_.io_diffCommits_info_78_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_78_pdest!=rhs_.io_diffCommits_info_78_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_78_pdest=0x%0h while the rhs_.io_diffCommits_info_78_pdest=0x%0h",this.io_diffCommits_info_78_pdest,rhs_.io_diffCommits_info_78_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_78_rfWen!=rhs_.io_diffCommits_info_78_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_78_rfWen=0x%0h while the rhs_.io_diffCommits_info_78_rfWen=0x%0h",this.io_diffCommits_info_78_rfWen,rhs_.io_diffCommits_info_78_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_78_fpWen!=rhs_.io_diffCommits_info_78_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_78_fpWen=0x%0h while the rhs_.io_diffCommits_info_78_fpWen=0x%0h",this.io_diffCommits_info_78_fpWen,rhs_.io_diffCommits_info_78_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_78_vecWen!=rhs_.io_diffCommits_info_78_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_78_vecWen=0x%0h while the rhs_.io_diffCommits_info_78_vecWen=0x%0h",this.io_diffCommits_info_78_vecWen,rhs_.io_diffCommits_info_78_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_78_v0Wen!=rhs_.io_diffCommits_info_78_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_78_v0Wen=0x%0h while the rhs_.io_diffCommits_info_78_v0Wen=0x%0h",this.io_diffCommits_info_78_v0Wen,rhs_.io_diffCommits_info_78_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_78_vlWen!=rhs_.io_diffCommits_info_78_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_78_vlWen=0x%0h while the rhs_.io_diffCommits_info_78_vlWen=0x%0h",this.io_diffCommits_info_78_vlWen,rhs_.io_diffCommits_info_78_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_79_ldest!=rhs_.io_diffCommits_info_79_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_79_ldest=0x%0h while the rhs_.io_diffCommits_info_79_ldest=0x%0h",this.io_diffCommits_info_79_ldest,rhs_.io_diffCommits_info_79_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_79_pdest!=rhs_.io_diffCommits_info_79_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_79_pdest=0x%0h while the rhs_.io_diffCommits_info_79_pdest=0x%0h",this.io_diffCommits_info_79_pdest,rhs_.io_diffCommits_info_79_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_79_rfWen!=rhs_.io_diffCommits_info_79_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_79_rfWen=0x%0h while the rhs_.io_diffCommits_info_79_rfWen=0x%0h",this.io_diffCommits_info_79_rfWen,rhs_.io_diffCommits_info_79_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_79_fpWen!=rhs_.io_diffCommits_info_79_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_79_fpWen=0x%0h while the rhs_.io_diffCommits_info_79_fpWen=0x%0h",this.io_diffCommits_info_79_fpWen,rhs_.io_diffCommits_info_79_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_79_vecWen!=rhs_.io_diffCommits_info_79_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_79_vecWen=0x%0h while the rhs_.io_diffCommits_info_79_vecWen=0x%0h",this.io_diffCommits_info_79_vecWen,rhs_.io_diffCommits_info_79_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_79_v0Wen!=rhs_.io_diffCommits_info_79_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_79_v0Wen=0x%0h while the rhs_.io_diffCommits_info_79_v0Wen=0x%0h",this.io_diffCommits_info_79_v0Wen,rhs_.io_diffCommits_info_79_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_79_vlWen!=rhs_.io_diffCommits_info_79_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_79_vlWen=0x%0h while the rhs_.io_diffCommits_info_79_vlWen=0x%0h",this.io_diffCommits_info_79_vlWen,rhs_.io_diffCommits_info_79_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_80_ldest!=rhs_.io_diffCommits_info_80_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_80_ldest=0x%0h while the rhs_.io_diffCommits_info_80_ldest=0x%0h",this.io_diffCommits_info_80_ldest,rhs_.io_diffCommits_info_80_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_80_pdest!=rhs_.io_diffCommits_info_80_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_80_pdest=0x%0h while the rhs_.io_diffCommits_info_80_pdest=0x%0h",this.io_diffCommits_info_80_pdest,rhs_.io_diffCommits_info_80_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_80_rfWen!=rhs_.io_diffCommits_info_80_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_80_rfWen=0x%0h while the rhs_.io_diffCommits_info_80_rfWen=0x%0h",this.io_diffCommits_info_80_rfWen,rhs_.io_diffCommits_info_80_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_80_fpWen!=rhs_.io_diffCommits_info_80_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_80_fpWen=0x%0h while the rhs_.io_diffCommits_info_80_fpWen=0x%0h",this.io_diffCommits_info_80_fpWen,rhs_.io_diffCommits_info_80_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_80_vecWen!=rhs_.io_diffCommits_info_80_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_80_vecWen=0x%0h while the rhs_.io_diffCommits_info_80_vecWen=0x%0h",this.io_diffCommits_info_80_vecWen,rhs_.io_diffCommits_info_80_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_80_v0Wen!=rhs_.io_diffCommits_info_80_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_80_v0Wen=0x%0h while the rhs_.io_diffCommits_info_80_v0Wen=0x%0h",this.io_diffCommits_info_80_v0Wen,rhs_.io_diffCommits_info_80_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_80_vlWen!=rhs_.io_diffCommits_info_80_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_80_vlWen=0x%0h while the rhs_.io_diffCommits_info_80_vlWen=0x%0h",this.io_diffCommits_info_80_vlWen,rhs_.io_diffCommits_info_80_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_81_ldest!=rhs_.io_diffCommits_info_81_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_81_ldest=0x%0h while the rhs_.io_diffCommits_info_81_ldest=0x%0h",this.io_diffCommits_info_81_ldest,rhs_.io_diffCommits_info_81_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_81_pdest!=rhs_.io_diffCommits_info_81_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_81_pdest=0x%0h while the rhs_.io_diffCommits_info_81_pdest=0x%0h",this.io_diffCommits_info_81_pdest,rhs_.io_diffCommits_info_81_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_81_rfWen!=rhs_.io_diffCommits_info_81_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_81_rfWen=0x%0h while the rhs_.io_diffCommits_info_81_rfWen=0x%0h",this.io_diffCommits_info_81_rfWen,rhs_.io_diffCommits_info_81_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_81_fpWen!=rhs_.io_diffCommits_info_81_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_81_fpWen=0x%0h while the rhs_.io_diffCommits_info_81_fpWen=0x%0h",this.io_diffCommits_info_81_fpWen,rhs_.io_diffCommits_info_81_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_81_vecWen!=rhs_.io_diffCommits_info_81_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_81_vecWen=0x%0h while the rhs_.io_diffCommits_info_81_vecWen=0x%0h",this.io_diffCommits_info_81_vecWen,rhs_.io_diffCommits_info_81_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_81_v0Wen!=rhs_.io_diffCommits_info_81_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_81_v0Wen=0x%0h while the rhs_.io_diffCommits_info_81_v0Wen=0x%0h",this.io_diffCommits_info_81_v0Wen,rhs_.io_diffCommits_info_81_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_81_vlWen!=rhs_.io_diffCommits_info_81_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_81_vlWen=0x%0h while the rhs_.io_diffCommits_info_81_vlWen=0x%0h",this.io_diffCommits_info_81_vlWen,rhs_.io_diffCommits_info_81_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_82_ldest!=rhs_.io_diffCommits_info_82_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_82_ldest=0x%0h while the rhs_.io_diffCommits_info_82_ldest=0x%0h",this.io_diffCommits_info_82_ldest,rhs_.io_diffCommits_info_82_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_82_pdest!=rhs_.io_diffCommits_info_82_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_82_pdest=0x%0h while the rhs_.io_diffCommits_info_82_pdest=0x%0h",this.io_diffCommits_info_82_pdest,rhs_.io_diffCommits_info_82_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_82_rfWen!=rhs_.io_diffCommits_info_82_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_82_rfWen=0x%0h while the rhs_.io_diffCommits_info_82_rfWen=0x%0h",this.io_diffCommits_info_82_rfWen,rhs_.io_diffCommits_info_82_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_82_fpWen!=rhs_.io_diffCommits_info_82_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_82_fpWen=0x%0h while the rhs_.io_diffCommits_info_82_fpWen=0x%0h",this.io_diffCommits_info_82_fpWen,rhs_.io_diffCommits_info_82_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_82_vecWen!=rhs_.io_diffCommits_info_82_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_82_vecWen=0x%0h while the rhs_.io_diffCommits_info_82_vecWen=0x%0h",this.io_diffCommits_info_82_vecWen,rhs_.io_diffCommits_info_82_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_82_v0Wen!=rhs_.io_diffCommits_info_82_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_82_v0Wen=0x%0h while the rhs_.io_diffCommits_info_82_v0Wen=0x%0h",this.io_diffCommits_info_82_v0Wen,rhs_.io_diffCommits_info_82_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_82_vlWen!=rhs_.io_diffCommits_info_82_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_82_vlWen=0x%0h while the rhs_.io_diffCommits_info_82_vlWen=0x%0h",this.io_diffCommits_info_82_vlWen,rhs_.io_diffCommits_info_82_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_83_ldest!=rhs_.io_diffCommits_info_83_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_83_ldest=0x%0h while the rhs_.io_diffCommits_info_83_ldest=0x%0h",this.io_diffCommits_info_83_ldest,rhs_.io_diffCommits_info_83_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_83_pdest!=rhs_.io_diffCommits_info_83_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_83_pdest=0x%0h while the rhs_.io_diffCommits_info_83_pdest=0x%0h",this.io_diffCommits_info_83_pdest,rhs_.io_diffCommits_info_83_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_83_rfWen!=rhs_.io_diffCommits_info_83_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_83_rfWen=0x%0h while the rhs_.io_diffCommits_info_83_rfWen=0x%0h",this.io_diffCommits_info_83_rfWen,rhs_.io_diffCommits_info_83_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_83_fpWen!=rhs_.io_diffCommits_info_83_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_83_fpWen=0x%0h while the rhs_.io_diffCommits_info_83_fpWen=0x%0h",this.io_diffCommits_info_83_fpWen,rhs_.io_diffCommits_info_83_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_83_vecWen!=rhs_.io_diffCommits_info_83_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_83_vecWen=0x%0h while the rhs_.io_diffCommits_info_83_vecWen=0x%0h",this.io_diffCommits_info_83_vecWen,rhs_.io_diffCommits_info_83_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_83_v0Wen!=rhs_.io_diffCommits_info_83_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_83_v0Wen=0x%0h while the rhs_.io_diffCommits_info_83_v0Wen=0x%0h",this.io_diffCommits_info_83_v0Wen,rhs_.io_diffCommits_info_83_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_83_vlWen!=rhs_.io_diffCommits_info_83_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_83_vlWen=0x%0h while the rhs_.io_diffCommits_info_83_vlWen=0x%0h",this.io_diffCommits_info_83_vlWen,rhs_.io_diffCommits_info_83_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_84_ldest!=rhs_.io_diffCommits_info_84_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_84_ldest=0x%0h while the rhs_.io_diffCommits_info_84_ldest=0x%0h",this.io_diffCommits_info_84_ldest,rhs_.io_diffCommits_info_84_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_84_pdest!=rhs_.io_diffCommits_info_84_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_84_pdest=0x%0h while the rhs_.io_diffCommits_info_84_pdest=0x%0h",this.io_diffCommits_info_84_pdest,rhs_.io_diffCommits_info_84_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_84_rfWen!=rhs_.io_diffCommits_info_84_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_84_rfWen=0x%0h while the rhs_.io_diffCommits_info_84_rfWen=0x%0h",this.io_diffCommits_info_84_rfWen,rhs_.io_diffCommits_info_84_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_84_fpWen!=rhs_.io_diffCommits_info_84_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_84_fpWen=0x%0h while the rhs_.io_diffCommits_info_84_fpWen=0x%0h",this.io_diffCommits_info_84_fpWen,rhs_.io_diffCommits_info_84_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_84_vecWen!=rhs_.io_diffCommits_info_84_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_84_vecWen=0x%0h while the rhs_.io_diffCommits_info_84_vecWen=0x%0h",this.io_diffCommits_info_84_vecWen,rhs_.io_diffCommits_info_84_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_84_v0Wen!=rhs_.io_diffCommits_info_84_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_84_v0Wen=0x%0h while the rhs_.io_diffCommits_info_84_v0Wen=0x%0h",this.io_diffCommits_info_84_v0Wen,rhs_.io_diffCommits_info_84_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_84_vlWen!=rhs_.io_diffCommits_info_84_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_84_vlWen=0x%0h while the rhs_.io_diffCommits_info_84_vlWen=0x%0h",this.io_diffCommits_info_84_vlWen,rhs_.io_diffCommits_info_84_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_85_ldest!=rhs_.io_diffCommits_info_85_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_85_ldest=0x%0h while the rhs_.io_diffCommits_info_85_ldest=0x%0h",this.io_diffCommits_info_85_ldest,rhs_.io_diffCommits_info_85_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_85_pdest!=rhs_.io_diffCommits_info_85_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_85_pdest=0x%0h while the rhs_.io_diffCommits_info_85_pdest=0x%0h",this.io_diffCommits_info_85_pdest,rhs_.io_diffCommits_info_85_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_85_rfWen!=rhs_.io_diffCommits_info_85_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_85_rfWen=0x%0h while the rhs_.io_diffCommits_info_85_rfWen=0x%0h",this.io_diffCommits_info_85_rfWen,rhs_.io_diffCommits_info_85_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_85_fpWen!=rhs_.io_diffCommits_info_85_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_85_fpWen=0x%0h while the rhs_.io_diffCommits_info_85_fpWen=0x%0h",this.io_diffCommits_info_85_fpWen,rhs_.io_diffCommits_info_85_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_85_vecWen!=rhs_.io_diffCommits_info_85_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_85_vecWen=0x%0h while the rhs_.io_diffCommits_info_85_vecWen=0x%0h",this.io_diffCommits_info_85_vecWen,rhs_.io_diffCommits_info_85_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_85_v0Wen!=rhs_.io_diffCommits_info_85_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_85_v0Wen=0x%0h while the rhs_.io_diffCommits_info_85_v0Wen=0x%0h",this.io_diffCommits_info_85_v0Wen,rhs_.io_diffCommits_info_85_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_85_vlWen!=rhs_.io_diffCommits_info_85_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_85_vlWen=0x%0h while the rhs_.io_diffCommits_info_85_vlWen=0x%0h",this.io_diffCommits_info_85_vlWen,rhs_.io_diffCommits_info_85_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_86_ldest!=rhs_.io_diffCommits_info_86_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_86_ldest=0x%0h while the rhs_.io_diffCommits_info_86_ldest=0x%0h",this.io_diffCommits_info_86_ldest,rhs_.io_diffCommits_info_86_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_86_pdest!=rhs_.io_diffCommits_info_86_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_86_pdest=0x%0h while the rhs_.io_diffCommits_info_86_pdest=0x%0h",this.io_diffCommits_info_86_pdest,rhs_.io_diffCommits_info_86_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_86_rfWen!=rhs_.io_diffCommits_info_86_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_86_rfWen=0x%0h while the rhs_.io_diffCommits_info_86_rfWen=0x%0h",this.io_diffCommits_info_86_rfWen,rhs_.io_diffCommits_info_86_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_86_fpWen!=rhs_.io_diffCommits_info_86_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_86_fpWen=0x%0h while the rhs_.io_diffCommits_info_86_fpWen=0x%0h",this.io_diffCommits_info_86_fpWen,rhs_.io_diffCommits_info_86_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_86_vecWen!=rhs_.io_diffCommits_info_86_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_86_vecWen=0x%0h while the rhs_.io_diffCommits_info_86_vecWen=0x%0h",this.io_diffCommits_info_86_vecWen,rhs_.io_diffCommits_info_86_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_86_v0Wen!=rhs_.io_diffCommits_info_86_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_86_v0Wen=0x%0h while the rhs_.io_diffCommits_info_86_v0Wen=0x%0h",this.io_diffCommits_info_86_v0Wen,rhs_.io_diffCommits_info_86_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_86_vlWen!=rhs_.io_diffCommits_info_86_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_86_vlWen=0x%0h while the rhs_.io_diffCommits_info_86_vlWen=0x%0h",this.io_diffCommits_info_86_vlWen,rhs_.io_diffCommits_info_86_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_87_ldest!=rhs_.io_diffCommits_info_87_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_87_ldest=0x%0h while the rhs_.io_diffCommits_info_87_ldest=0x%0h",this.io_diffCommits_info_87_ldest,rhs_.io_diffCommits_info_87_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_87_pdest!=rhs_.io_diffCommits_info_87_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_87_pdest=0x%0h while the rhs_.io_diffCommits_info_87_pdest=0x%0h",this.io_diffCommits_info_87_pdest,rhs_.io_diffCommits_info_87_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_87_rfWen!=rhs_.io_diffCommits_info_87_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_87_rfWen=0x%0h while the rhs_.io_diffCommits_info_87_rfWen=0x%0h",this.io_diffCommits_info_87_rfWen,rhs_.io_diffCommits_info_87_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_87_fpWen!=rhs_.io_diffCommits_info_87_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_87_fpWen=0x%0h while the rhs_.io_diffCommits_info_87_fpWen=0x%0h",this.io_diffCommits_info_87_fpWen,rhs_.io_diffCommits_info_87_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_87_vecWen!=rhs_.io_diffCommits_info_87_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_87_vecWen=0x%0h while the rhs_.io_diffCommits_info_87_vecWen=0x%0h",this.io_diffCommits_info_87_vecWen,rhs_.io_diffCommits_info_87_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_87_v0Wen!=rhs_.io_diffCommits_info_87_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_87_v0Wen=0x%0h while the rhs_.io_diffCommits_info_87_v0Wen=0x%0h",this.io_diffCommits_info_87_v0Wen,rhs_.io_diffCommits_info_87_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_87_vlWen!=rhs_.io_diffCommits_info_87_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_87_vlWen=0x%0h while the rhs_.io_diffCommits_info_87_vlWen=0x%0h",this.io_diffCommits_info_87_vlWen,rhs_.io_diffCommits_info_87_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_88_ldest!=rhs_.io_diffCommits_info_88_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_88_ldest=0x%0h while the rhs_.io_diffCommits_info_88_ldest=0x%0h",this.io_diffCommits_info_88_ldest,rhs_.io_diffCommits_info_88_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_88_pdest!=rhs_.io_diffCommits_info_88_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_88_pdest=0x%0h while the rhs_.io_diffCommits_info_88_pdest=0x%0h",this.io_diffCommits_info_88_pdest,rhs_.io_diffCommits_info_88_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_88_rfWen!=rhs_.io_diffCommits_info_88_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_88_rfWen=0x%0h while the rhs_.io_diffCommits_info_88_rfWen=0x%0h",this.io_diffCommits_info_88_rfWen,rhs_.io_diffCommits_info_88_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_88_fpWen!=rhs_.io_diffCommits_info_88_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_88_fpWen=0x%0h while the rhs_.io_diffCommits_info_88_fpWen=0x%0h",this.io_diffCommits_info_88_fpWen,rhs_.io_diffCommits_info_88_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_88_vecWen!=rhs_.io_diffCommits_info_88_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_88_vecWen=0x%0h while the rhs_.io_diffCommits_info_88_vecWen=0x%0h",this.io_diffCommits_info_88_vecWen,rhs_.io_diffCommits_info_88_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_88_v0Wen!=rhs_.io_diffCommits_info_88_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_88_v0Wen=0x%0h while the rhs_.io_diffCommits_info_88_v0Wen=0x%0h",this.io_diffCommits_info_88_v0Wen,rhs_.io_diffCommits_info_88_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_88_vlWen!=rhs_.io_diffCommits_info_88_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_88_vlWen=0x%0h while the rhs_.io_diffCommits_info_88_vlWen=0x%0h",this.io_diffCommits_info_88_vlWen,rhs_.io_diffCommits_info_88_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_89_ldest!=rhs_.io_diffCommits_info_89_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_89_ldest=0x%0h while the rhs_.io_diffCommits_info_89_ldest=0x%0h",this.io_diffCommits_info_89_ldest,rhs_.io_diffCommits_info_89_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_89_pdest!=rhs_.io_diffCommits_info_89_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_89_pdest=0x%0h while the rhs_.io_diffCommits_info_89_pdest=0x%0h",this.io_diffCommits_info_89_pdest,rhs_.io_diffCommits_info_89_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_89_rfWen!=rhs_.io_diffCommits_info_89_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_89_rfWen=0x%0h while the rhs_.io_diffCommits_info_89_rfWen=0x%0h",this.io_diffCommits_info_89_rfWen,rhs_.io_diffCommits_info_89_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_89_fpWen!=rhs_.io_diffCommits_info_89_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_89_fpWen=0x%0h while the rhs_.io_diffCommits_info_89_fpWen=0x%0h",this.io_diffCommits_info_89_fpWen,rhs_.io_diffCommits_info_89_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_89_vecWen!=rhs_.io_diffCommits_info_89_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_89_vecWen=0x%0h while the rhs_.io_diffCommits_info_89_vecWen=0x%0h",this.io_diffCommits_info_89_vecWen,rhs_.io_diffCommits_info_89_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_89_v0Wen!=rhs_.io_diffCommits_info_89_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_89_v0Wen=0x%0h while the rhs_.io_diffCommits_info_89_v0Wen=0x%0h",this.io_diffCommits_info_89_v0Wen,rhs_.io_diffCommits_info_89_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_89_vlWen!=rhs_.io_diffCommits_info_89_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_89_vlWen=0x%0h while the rhs_.io_diffCommits_info_89_vlWen=0x%0h",this.io_diffCommits_info_89_vlWen,rhs_.io_diffCommits_info_89_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_90_ldest!=rhs_.io_diffCommits_info_90_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_90_ldest=0x%0h while the rhs_.io_diffCommits_info_90_ldest=0x%0h",this.io_diffCommits_info_90_ldest,rhs_.io_diffCommits_info_90_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_90_pdest!=rhs_.io_diffCommits_info_90_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_90_pdest=0x%0h while the rhs_.io_diffCommits_info_90_pdest=0x%0h",this.io_diffCommits_info_90_pdest,rhs_.io_diffCommits_info_90_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_90_rfWen!=rhs_.io_diffCommits_info_90_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_90_rfWen=0x%0h while the rhs_.io_diffCommits_info_90_rfWen=0x%0h",this.io_diffCommits_info_90_rfWen,rhs_.io_diffCommits_info_90_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_90_fpWen!=rhs_.io_diffCommits_info_90_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_90_fpWen=0x%0h while the rhs_.io_diffCommits_info_90_fpWen=0x%0h",this.io_diffCommits_info_90_fpWen,rhs_.io_diffCommits_info_90_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_90_vecWen!=rhs_.io_diffCommits_info_90_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_90_vecWen=0x%0h while the rhs_.io_diffCommits_info_90_vecWen=0x%0h",this.io_diffCommits_info_90_vecWen,rhs_.io_diffCommits_info_90_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_90_v0Wen!=rhs_.io_diffCommits_info_90_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_90_v0Wen=0x%0h while the rhs_.io_diffCommits_info_90_v0Wen=0x%0h",this.io_diffCommits_info_90_v0Wen,rhs_.io_diffCommits_info_90_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_90_vlWen!=rhs_.io_diffCommits_info_90_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_90_vlWen=0x%0h while the rhs_.io_diffCommits_info_90_vlWen=0x%0h",this.io_diffCommits_info_90_vlWen,rhs_.io_diffCommits_info_90_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_91_ldest!=rhs_.io_diffCommits_info_91_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_91_ldest=0x%0h while the rhs_.io_diffCommits_info_91_ldest=0x%0h",this.io_diffCommits_info_91_ldest,rhs_.io_diffCommits_info_91_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_91_pdest!=rhs_.io_diffCommits_info_91_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_91_pdest=0x%0h while the rhs_.io_diffCommits_info_91_pdest=0x%0h",this.io_diffCommits_info_91_pdest,rhs_.io_diffCommits_info_91_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_91_rfWen!=rhs_.io_diffCommits_info_91_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_91_rfWen=0x%0h while the rhs_.io_diffCommits_info_91_rfWen=0x%0h",this.io_diffCommits_info_91_rfWen,rhs_.io_diffCommits_info_91_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_91_fpWen!=rhs_.io_diffCommits_info_91_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_91_fpWen=0x%0h while the rhs_.io_diffCommits_info_91_fpWen=0x%0h",this.io_diffCommits_info_91_fpWen,rhs_.io_diffCommits_info_91_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_91_vecWen!=rhs_.io_diffCommits_info_91_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_91_vecWen=0x%0h while the rhs_.io_diffCommits_info_91_vecWen=0x%0h",this.io_diffCommits_info_91_vecWen,rhs_.io_diffCommits_info_91_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_91_v0Wen!=rhs_.io_diffCommits_info_91_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_91_v0Wen=0x%0h while the rhs_.io_diffCommits_info_91_v0Wen=0x%0h",this.io_diffCommits_info_91_v0Wen,rhs_.io_diffCommits_info_91_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_91_vlWen!=rhs_.io_diffCommits_info_91_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_91_vlWen=0x%0h while the rhs_.io_diffCommits_info_91_vlWen=0x%0h",this.io_diffCommits_info_91_vlWen,rhs_.io_diffCommits_info_91_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_92_ldest!=rhs_.io_diffCommits_info_92_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_92_ldest=0x%0h while the rhs_.io_diffCommits_info_92_ldest=0x%0h",this.io_diffCommits_info_92_ldest,rhs_.io_diffCommits_info_92_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_92_pdest!=rhs_.io_diffCommits_info_92_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_92_pdest=0x%0h while the rhs_.io_diffCommits_info_92_pdest=0x%0h",this.io_diffCommits_info_92_pdest,rhs_.io_diffCommits_info_92_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_92_rfWen!=rhs_.io_diffCommits_info_92_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_92_rfWen=0x%0h while the rhs_.io_diffCommits_info_92_rfWen=0x%0h",this.io_diffCommits_info_92_rfWen,rhs_.io_diffCommits_info_92_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_92_fpWen!=rhs_.io_diffCommits_info_92_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_92_fpWen=0x%0h while the rhs_.io_diffCommits_info_92_fpWen=0x%0h",this.io_diffCommits_info_92_fpWen,rhs_.io_diffCommits_info_92_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_92_vecWen!=rhs_.io_diffCommits_info_92_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_92_vecWen=0x%0h while the rhs_.io_diffCommits_info_92_vecWen=0x%0h",this.io_diffCommits_info_92_vecWen,rhs_.io_diffCommits_info_92_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_92_v0Wen!=rhs_.io_diffCommits_info_92_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_92_v0Wen=0x%0h while the rhs_.io_diffCommits_info_92_v0Wen=0x%0h",this.io_diffCommits_info_92_v0Wen,rhs_.io_diffCommits_info_92_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_92_vlWen!=rhs_.io_diffCommits_info_92_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_92_vlWen=0x%0h while the rhs_.io_diffCommits_info_92_vlWen=0x%0h",this.io_diffCommits_info_92_vlWen,rhs_.io_diffCommits_info_92_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_93_ldest!=rhs_.io_diffCommits_info_93_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_93_ldest=0x%0h while the rhs_.io_diffCommits_info_93_ldest=0x%0h",this.io_diffCommits_info_93_ldest,rhs_.io_diffCommits_info_93_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_93_pdest!=rhs_.io_diffCommits_info_93_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_93_pdest=0x%0h while the rhs_.io_diffCommits_info_93_pdest=0x%0h",this.io_diffCommits_info_93_pdest,rhs_.io_diffCommits_info_93_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_93_rfWen!=rhs_.io_diffCommits_info_93_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_93_rfWen=0x%0h while the rhs_.io_diffCommits_info_93_rfWen=0x%0h",this.io_diffCommits_info_93_rfWen,rhs_.io_diffCommits_info_93_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_93_fpWen!=rhs_.io_diffCommits_info_93_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_93_fpWen=0x%0h while the rhs_.io_diffCommits_info_93_fpWen=0x%0h",this.io_diffCommits_info_93_fpWen,rhs_.io_diffCommits_info_93_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_93_vecWen!=rhs_.io_diffCommits_info_93_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_93_vecWen=0x%0h while the rhs_.io_diffCommits_info_93_vecWen=0x%0h",this.io_diffCommits_info_93_vecWen,rhs_.io_diffCommits_info_93_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_93_v0Wen!=rhs_.io_diffCommits_info_93_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_93_v0Wen=0x%0h while the rhs_.io_diffCommits_info_93_v0Wen=0x%0h",this.io_diffCommits_info_93_v0Wen,rhs_.io_diffCommits_info_93_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_93_vlWen!=rhs_.io_diffCommits_info_93_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_93_vlWen=0x%0h while the rhs_.io_diffCommits_info_93_vlWen=0x%0h",this.io_diffCommits_info_93_vlWen,rhs_.io_diffCommits_info_93_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_94_ldest!=rhs_.io_diffCommits_info_94_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_94_ldest=0x%0h while the rhs_.io_diffCommits_info_94_ldest=0x%0h",this.io_diffCommits_info_94_ldest,rhs_.io_diffCommits_info_94_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_94_pdest!=rhs_.io_diffCommits_info_94_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_94_pdest=0x%0h while the rhs_.io_diffCommits_info_94_pdest=0x%0h",this.io_diffCommits_info_94_pdest,rhs_.io_diffCommits_info_94_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_94_rfWen!=rhs_.io_diffCommits_info_94_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_94_rfWen=0x%0h while the rhs_.io_diffCommits_info_94_rfWen=0x%0h",this.io_diffCommits_info_94_rfWen,rhs_.io_diffCommits_info_94_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_94_fpWen!=rhs_.io_diffCommits_info_94_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_94_fpWen=0x%0h while the rhs_.io_diffCommits_info_94_fpWen=0x%0h",this.io_diffCommits_info_94_fpWen,rhs_.io_diffCommits_info_94_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_94_vecWen!=rhs_.io_diffCommits_info_94_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_94_vecWen=0x%0h while the rhs_.io_diffCommits_info_94_vecWen=0x%0h",this.io_diffCommits_info_94_vecWen,rhs_.io_diffCommits_info_94_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_94_v0Wen!=rhs_.io_diffCommits_info_94_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_94_v0Wen=0x%0h while the rhs_.io_diffCommits_info_94_v0Wen=0x%0h",this.io_diffCommits_info_94_v0Wen,rhs_.io_diffCommits_info_94_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_94_vlWen!=rhs_.io_diffCommits_info_94_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_94_vlWen=0x%0h while the rhs_.io_diffCommits_info_94_vlWen=0x%0h",this.io_diffCommits_info_94_vlWen,rhs_.io_diffCommits_info_94_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_95_ldest!=rhs_.io_diffCommits_info_95_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_95_ldest=0x%0h while the rhs_.io_diffCommits_info_95_ldest=0x%0h",this.io_diffCommits_info_95_ldest,rhs_.io_diffCommits_info_95_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_95_pdest!=rhs_.io_diffCommits_info_95_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_95_pdest=0x%0h while the rhs_.io_diffCommits_info_95_pdest=0x%0h",this.io_diffCommits_info_95_pdest,rhs_.io_diffCommits_info_95_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_95_rfWen!=rhs_.io_diffCommits_info_95_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_95_rfWen=0x%0h while the rhs_.io_diffCommits_info_95_rfWen=0x%0h",this.io_diffCommits_info_95_rfWen,rhs_.io_diffCommits_info_95_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_95_fpWen!=rhs_.io_diffCommits_info_95_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_95_fpWen=0x%0h while the rhs_.io_diffCommits_info_95_fpWen=0x%0h",this.io_diffCommits_info_95_fpWen,rhs_.io_diffCommits_info_95_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_95_vecWen!=rhs_.io_diffCommits_info_95_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_95_vecWen=0x%0h while the rhs_.io_diffCommits_info_95_vecWen=0x%0h",this.io_diffCommits_info_95_vecWen,rhs_.io_diffCommits_info_95_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_95_v0Wen!=rhs_.io_diffCommits_info_95_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_95_v0Wen=0x%0h while the rhs_.io_diffCommits_info_95_v0Wen=0x%0h",this.io_diffCommits_info_95_v0Wen,rhs_.io_diffCommits_info_95_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_95_vlWen!=rhs_.io_diffCommits_info_95_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_95_vlWen=0x%0h while the rhs_.io_diffCommits_info_95_vlWen=0x%0h",this.io_diffCommits_info_95_vlWen,rhs_.io_diffCommits_info_95_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_96_ldest!=rhs_.io_diffCommits_info_96_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_96_ldest=0x%0h while the rhs_.io_diffCommits_info_96_ldest=0x%0h",this.io_diffCommits_info_96_ldest,rhs_.io_diffCommits_info_96_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_96_pdest!=rhs_.io_diffCommits_info_96_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_96_pdest=0x%0h while the rhs_.io_diffCommits_info_96_pdest=0x%0h",this.io_diffCommits_info_96_pdest,rhs_.io_diffCommits_info_96_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_96_rfWen!=rhs_.io_diffCommits_info_96_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_96_rfWen=0x%0h while the rhs_.io_diffCommits_info_96_rfWen=0x%0h",this.io_diffCommits_info_96_rfWen,rhs_.io_diffCommits_info_96_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_96_fpWen!=rhs_.io_diffCommits_info_96_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_96_fpWen=0x%0h while the rhs_.io_diffCommits_info_96_fpWen=0x%0h",this.io_diffCommits_info_96_fpWen,rhs_.io_diffCommits_info_96_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_96_vecWen!=rhs_.io_diffCommits_info_96_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_96_vecWen=0x%0h while the rhs_.io_diffCommits_info_96_vecWen=0x%0h",this.io_diffCommits_info_96_vecWen,rhs_.io_diffCommits_info_96_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_96_v0Wen!=rhs_.io_diffCommits_info_96_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_96_v0Wen=0x%0h while the rhs_.io_diffCommits_info_96_v0Wen=0x%0h",this.io_diffCommits_info_96_v0Wen,rhs_.io_diffCommits_info_96_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_96_vlWen!=rhs_.io_diffCommits_info_96_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_96_vlWen=0x%0h while the rhs_.io_diffCommits_info_96_vlWen=0x%0h",this.io_diffCommits_info_96_vlWen,rhs_.io_diffCommits_info_96_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_97_ldest!=rhs_.io_diffCommits_info_97_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_97_ldest=0x%0h while the rhs_.io_diffCommits_info_97_ldest=0x%0h",this.io_diffCommits_info_97_ldest,rhs_.io_diffCommits_info_97_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_97_pdest!=rhs_.io_diffCommits_info_97_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_97_pdest=0x%0h while the rhs_.io_diffCommits_info_97_pdest=0x%0h",this.io_diffCommits_info_97_pdest,rhs_.io_diffCommits_info_97_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_97_rfWen!=rhs_.io_diffCommits_info_97_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_97_rfWen=0x%0h while the rhs_.io_diffCommits_info_97_rfWen=0x%0h",this.io_diffCommits_info_97_rfWen,rhs_.io_diffCommits_info_97_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_97_fpWen!=rhs_.io_diffCommits_info_97_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_97_fpWen=0x%0h while the rhs_.io_diffCommits_info_97_fpWen=0x%0h",this.io_diffCommits_info_97_fpWen,rhs_.io_diffCommits_info_97_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_97_vecWen!=rhs_.io_diffCommits_info_97_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_97_vecWen=0x%0h while the rhs_.io_diffCommits_info_97_vecWen=0x%0h",this.io_diffCommits_info_97_vecWen,rhs_.io_diffCommits_info_97_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_97_v0Wen!=rhs_.io_diffCommits_info_97_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_97_v0Wen=0x%0h while the rhs_.io_diffCommits_info_97_v0Wen=0x%0h",this.io_diffCommits_info_97_v0Wen,rhs_.io_diffCommits_info_97_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_97_vlWen!=rhs_.io_diffCommits_info_97_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_97_vlWen=0x%0h while the rhs_.io_diffCommits_info_97_vlWen=0x%0h",this.io_diffCommits_info_97_vlWen,rhs_.io_diffCommits_info_97_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_98_ldest!=rhs_.io_diffCommits_info_98_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_98_ldest=0x%0h while the rhs_.io_diffCommits_info_98_ldest=0x%0h",this.io_diffCommits_info_98_ldest,rhs_.io_diffCommits_info_98_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_98_pdest!=rhs_.io_diffCommits_info_98_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_98_pdest=0x%0h while the rhs_.io_diffCommits_info_98_pdest=0x%0h",this.io_diffCommits_info_98_pdest,rhs_.io_diffCommits_info_98_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_98_rfWen!=rhs_.io_diffCommits_info_98_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_98_rfWen=0x%0h while the rhs_.io_diffCommits_info_98_rfWen=0x%0h",this.io_diffCommits_info_98_rfWen,rhs_.io_diffCommits_info_98_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_98_fpWen!=rhs_.io_diffCommits_info_98_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_98_fpWen=0x%0h while the rhs_.io_diffCommits_info_98_fpWen=0x%0h",this.io_diffCommits_info_98_fpWen,rhs_.io_diffCommits_info_98_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_98_vecWen!=rhs_.io_diffCommits_info_98_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_98_vecWen=0x%0h while the rhs_.io_diffCommits_info_98_vecWen=0x%0h",this.io_diffCommits_info_98_vecWen,rhs_.io_diffCommits_info_98_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_98_v0Wen!=rhs_.io_diffCommits_info_98_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_98_v0Wen=0x%0h while the rhs_.io_diffCommits_info_98_v0Wen=0x%0h",this.io_diffCommits_info_98_v0Wen,rhs_.io_diffCommits_info_98_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_98_vlWen!=rhs_.io_diffCommits_info_98_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_98_vlWen=0x%0h while the rhs_.io_diffCommits_info_98_vlWen=0x%0h",this.io_diffCommits_info_98_vlWen,rhs_.io_diffCommits_info_98_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_99_ldest!=rhs_.io_diffCommits_info_99_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_99_ldest=0x%0h while the rhs_.io_diffCommits_info_99_ldest=0x%0h",this.io_diffCommits_info_99_ldest,rhs_.io_diffCommits_info_99_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_99_pdest!=rhs_.io_diffCommits_info_99_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_99_pdest=0x%0h while the rhs_.io_diffCommits_info_99_pdest=0x%0h",this.io_diffCommits_info_99_pdest,rhs_.io_diffCommits_info_99_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_99_rfWen!=rhs_.io_diffCommits_info_99_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_99_rfWen=0x%0h while the rhs_.io_diffCommits_info_99_rfWen=0x%0h",this.io_diffCommits_info_99_rfWen,rhs_.io_diffCommits_info_99_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_99_fpWen!=rhs_.io_diffCommits_info_99_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_99_fpWen=0x%0h while the rhs_.io_diffCommits_info_99_fpWen=0x%0h",this.io_diffCommits_info_99_fpWen,rhs_.io_diffCommits_info_99_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_99_vecWen!=rhs_.io_diffCommits_info_99_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_99_vecWen=0x%0h while the rhs_.io_diffCommits_info_99_vecWen=0x%0h",this.io_diffCommits_info_99_vecWen,rhs_.io_diffCommits_info_99_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_99_v0Wen!=rhs_.io_diffCommits_info_99_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_99_v0Wen=0x%0h while the rhs_.io_diffCommits_info_99_v0Wen=0x%0h",this.io_diffCommits_info_99_v0Wen,rhs_.io_diffCommits_info_99_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_99_vlWen!=rhs_.io_diffCommits_info_99_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_99_vlWen=0x%0h while the rhs_.io_diffCommits_info_99_vlWen=0x%0h",this.io_diffCommits_info_99_vlWen,rhs_.io_diffCommits_info_99_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_100_ldest!=rhs_.io_diffCommits_info_100_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_100_ldest=0x%0h while the rhs_.io_diffCommits_info_100_ldest=0x%0h",this.io_diffCommits_info_100_ldest,rhs_.io_diffCommits_info_100_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_100_pdest!=rhs_.io_diffCommits_info_100_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_100_pdest=0x%0h while the rhs_.io_diffCommits_info_100_pdest=0x%0h",this.io_diffCommits_info_100_pdest,rhs_.io_diffCommits_info_100_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_100_rfWen!=rhs_.io_diffCommits_info_100_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_100_rfWen=0x%0h while the rhs_.io_diffCommits_info_100_rfWen=0x%0h",this.io_diffCommits_info_100_rfWen,rhs_.io_diffCommits_info_100_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_100_fpWen!=rhs_.io_diffCommits_info_100_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_100_fpWen=0x%0h while the rhs_.io_diffCommits_info_100_fpWen=0x%0h",this.io_diffCommits_info_100_fpWen,rhs_.io_diffCommits_info_100_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_100_vecWen!=rhs_.io_diffCommits_info_100_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_100_vecWen=0x%0h while the rhs_.io_diffCommits_info_100_vecWen=0x%0h",this.io_diffCommits_info_100_vecWen,rhs_.io_diffCommits_info_100_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_100_v0Wen!=rhs_.io_diffCommits_info_100_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_100_v0Wen=0x%0h while the rhs_.io_diffCommits_info_100_v0Wen=0x%0h",this.io_diffCommits_info_100_v0Wen,rhs_.io_diffCommits_info_100_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_100_vlWen!=rhs_.io_diffCommits_info_100_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_100_vlWen=0x%0h while the rhs_.io_diffCommits_info_100_vlWen=0x%0h",this.io_diffCommits_info_100_vlWen,rhs_.io_diffCommits_info_100_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_101_ldest!=rhs_.io_diffCommits_info_101_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_101_ldest=0x%0h while the rhs_.io_diffCommits_info_101_ldest=0x%0h",this.io_diffCommits_info_101_ldest,rhs_.io_diffCommits_info_101_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_101_pdest!=rhs_.io_diffCommits_info_101_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_101_pdest=0x%0h while the rhs_.io_diffCommits_info_101_pdest=0x%0h",this.io_diffCommits_info_101_pdest,rhs_.io_diffCommits_info_101_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_101_rfWen!=rhs_.io_diffCommits_info_101_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_101_rfWen=0x%0h while the rhs_.io_diffCommits_info_101_rfWen=0x%0h",this.io_diffCommits_info_101_rfWen,rhs_.io_diffCommits_info_101_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_101_fpWen!=rhs_.io_diffCommits_info_101_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_101_fpWen=0x%0h while the rhs_.io_diffCommits_info_101_fpWen=0x%0h",this.io_diffCommits_info_101_fpWen,rhs_.io_diffCommits_info_101_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_101_vecWen!=rhs_.io_diffCommits_info_101_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_101_vecWen=0x%0h while the rhs_.io_diffCommits_info_101_vecWen=0x%0h",this.io_diffCommits_info_101_vecWen,rhs_.io_diffCommits_info_101_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_101_v0Wen!=rhs_.io_diffCommits_info_101_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_101_v0Wen=0x%0h while the rhs_.io_diffCommits_info_101_v0Wen=0x%0h",this.io_diffCommits_info_101_v0Wen,rhs_.io_diffCommits_info_101_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_101_vlWen!=rhs_.io_diffCommits_info_101_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_101_vlWen=0x%0h while the rhs_.io_diffCommits_info_101_vlWen=0x%0h",this.io_diffCommits_info_101_vlWen,rhs_.io_diffCommits_info_101_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_102_ldest!=rhs_.io_diffCommits_info_102_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_102_ldest=0x%0h while the rhs_.io_diffCommits_info_102_ldest=0x%0h",this.io_diffCommits_info_102_ldest,rhs_.io_diffCommits_info_102_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_102_pdest!=rhs_.io_diffCommits_info_102_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_102_pdest=0x%0h while the rhs_.io_diffCommits_info_102_pdest=0x%0h",this.io_diffCommits_info_102_pdest,rhs_.io_diffCommits_info_102_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_102_rfWen!=rhs_.io_diffCommits_info_102_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_102_rfWen=0x%0h while the rhs_.io_diffCommits_info_102_rfWen=0x%0h",this.io_diffCommits_info_102_rfWen,rhs_.io_diffCommits_info_102_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_102_fpWen!=rhs_.io_diffCommits_info_102_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_102_fpWen=0x%0h while the rhs_.io_diffCommits_info_102_fpWen=0x%0h",this.io_diffCommits_info_102_fpWen,rhs_.io_diffCommits_info_102_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_102_vecWen!=rhs_.io_diffCommits_info_102_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_102_vecWen=0x%0h while the rhs_.io_diffCommits_info_102_vecWen=0x%0h",this.io_diffCommits_info_102_vecWen,rhs_.io_diffCommits_info_102_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_102_v0Wen!=rhs_.io_diffCommits_info_102_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_102_v0Wen=0x%0h while the rhs_.io_diffCommits_info_102_v0Wen=0x%0h",this.io_diffCommits_info_102_v0Wen,rhs_.io_diffCommits_info_102_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_102_vlWen!=rhs_.io_diffCommits_info_102_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_102_vlWen=0x%0h while the rhs_.io_diffCommits_info_102_vlWen=0x%0h",this.io_diffCommits_info_102_vlWen,rhs_.io_diffCommits_info_102_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_103_ldest!=rhs_.io_diffCommits_info_103_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_103_ldest=0x%0h while the rhs_.io_diffCommits_info_103_ldest=0x%0h",this.io_diffCommits_info_103_ldest,rhs_.io_diffCommits_info_103_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_103_pdest!=rhs_.io_diffCommits_info_103_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_103_pdest=0x%0h while the rhs_.io_diffCommits_info_103_pdest=0x%0h",this.io_diffCommits_info_103_pdest,rhs_.io_diffCommits_info_103_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_103_rfWen!=rhs_.io_diffCommits_info_103_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_103_rfWen=0x%0h while the rhs_.io_diffCommits_info_103_rfWen=0x%0h",this.io_diffCommits_info_103_rfWen,rhs_.io_diffCommits_info_103_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_103_fpWen!=rhs_.io_diffCommits_info_103_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_103_fpWen=0x%0h while the rhs_.io_diffCommits_info_103_fpWen=0x%0h",this.io_diffCommits_info_103_fpWen,rhs_.io_diffCommits_info_103_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_103_vecWen!=rhs_.io_diffCommits_info_103_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_103_vecWen=0x%0h while the rhs_.io_diffCommits_info_103_vecWen=0x%0h",this.io_diffCommits_info_103_vecWen,rhs_.io_diffCommits_info_103_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_103_v0Wen!=rhs_.io_diffCommits_info_103_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_103_v0Wen=0x%0h while the rhs_.io_diffCommits_info_103_v0Wen=0x%0h",this.io_diffCommits_info_103_v0Wen,rhs_.io_diffCommits_info_103_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_103_vlWen!=rhs_.io_diffCommits_info_103_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_103_vlWen=0x%0h while the rhs_.io_diffCommits_info_103_vlWen=0x%0h",this.io_diffCommits_info_103_vlWen,rhs_.io_diffCommits_info_103_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_104_ldest!=rhs_.io_diffCommits_info_104_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_104_ldest=0x%0h while the rhs_.io_diffCommits_info_104_ldest=0x%0h",this.io_diffCommits_info_104_ldest,rhs_.io_diffCommits_info_104_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_104_pdest!=rhs_.io_diffCommits_info_104_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_104_pdest=0x%0h while the rhs_.io_diffCommits_info_104_pdest=0x%0h",this.io_diffCommits_info_104_pdest,rhs_.io_diffCommits_info_104_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_104_rfWen!=rhs_.io_diffCommits_info_104_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_104_rfWen=0x%0h while the rhs_.io_diffCommits_info_104_rfWen=0x%0h",this.io_diffCommits_info_104_rfWen,rhs_.io_diffCommits_info_104_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_104_fpWen!=rhs_.io_diffCommits_info_104_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_104_fpWen=0x%0h while the rhs_.io_diffCommits_info_104_fpWen=0x%0h",this.io_diffCommits_info_104_fpWen,rhs_.io_diffCommits_info_104_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_104_vecWen!=rhs_.io_diffCommits_info_104_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_104_vecWen=0x%0h while the rhs_.io_diffCommits_info_104_vecWen=0x%0h",this.io_diffCommits_info_104_vecWen,rhs_.io_diffCommits_info_104_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_104_v0Wen!=rhs_.io_diffCommits_info_104_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_104_v0Wen=0x%0h while the rhs_.io_diffCommits_info_104_v0Wen=0x%0h",this.io_diffCommits_info_104_v0Wen,rhs_.io_diffCommits_info_104_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_104_vlWen!=rhs_.io_diffCommits_info_104_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_104_vlWen=0x%0h while the rhs_.io_diffCommits_info_104_vlWen=0x%0h",this.io_diffCommits_info_104_vlWen,rhs_.io_diffCommits_info_104_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_105_ldest!=rhs_.io_diffCommits_info_105_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_105_ldest=0x%0h while the rhs_.io_diffCommits_info_105_ldest=0x%0h",this.io_diffCommits_info_105_ldest,rhs_.io_diffCommits_info_105_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_105_pdest!=rhs_.io_diffCommits_info_105_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_105_pdest=0x%0h while the rhs_.io_diffCommits_info_105_pdest=0x%0h",this.io_diffCommits_info_105_pdest,rhs_.io_diffCommits_info_105_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_105_rfWen!=rhs_.io_diffCommits_info_105_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_105_rfWen=0x%0h while the rhs_.io_diffCommits_info_105_rfWen=0x%0h",this.io_diffCommits_info_105_rfWen,rhs_.io_diffCommits_info_105_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_105_fpWen!=rhs_.io_diffCommits_info_105_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_105_fpWen=0x%0h while the rhs_.io_diffCommits_info_105_fpWen=0x%0h",this.io_diffCommits_info_105_fpWen,rhs_.io_diffCommits_info_105_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_105_vecWen!=rhs_.io_diffCommits_info_105_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_105_vecWen=0x%0h while the rhs_.io_diffCommits_info_105_vecWen=0x%0h",this.io_diffCommits_info_105_vecWen,rhs_.io_diffCommits_info_105_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_105_v0Wen!=rhs_.io_diffCommits_info_105_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_105_v0Wen=0x%0h while the rhs_.io_diffCommits_info_105_v0Wen=0x%0h",this.io_diffCommits_info_105_v0Wen,rhs_.io_diffCommits_info_105_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_105_vlWen!=rhs_.io_diffCommits_info_105_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_105_vlWen=0x%0h while the rhs_.io_diffCommits_info_105_vlWen=0x%0h",this.io_diffCommits_info_105_vlWen,rhs_.io_diffCommits_info_105_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_106_ldest!=rhs_.io_diffCommits_info_106_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_106_ldest=0x%0h while the rhs_.io_diffCommits_info_106_ldest=0x%0h",this.io_diffCommits_info_106_ldest,rhs_.io_diffCommits_info_106_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_106_pdest!=rhs_.io_diffCommits_info_106_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_106_pdest=0x%0h while the rhs_.io_diffCommits_info_106_pdest=0x%0h",this.io_diffCommits_info_106_pdest,rhs_.io_diffCommits_info_106_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_106_rfWen!=rhs_.io_diffCommits_info_106_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_106_rfWen=0x%0h while the rhs_.io_diffCommits_info_106_rfWen=0x%0h",this.io_diffCommits_info_106_rfWen,rhs_.io_diffCommits_info_106_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_106_fpWen!=rhs_.io_diffCommits_info_106_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_106_fpWen=0x%0h while the rhs_.io_diffCommits_info_106_fpWen=0x%0h",this.io_diffCommits_info_106_fpWen,rhs_.io_diffCommits_info_106_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_106_vecWen!=rhs_.io_diffCommits_info_106_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_106_vecWen=0x%0h while the rhs_.io_diffCommits_info_106_vecWen=0x%0h",this.io_diffCommits_info_106_vecWen,rhs_.io_diffCommits_info_106_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_106_v0Wen!=rhs_.io_diffCommits_info_106_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_106_v0Wen=0x%0h while the rhs_.io_diffCommits_info_106_v0Wen=0x%0h",this.io_diffCommits_info_106_v0Wen,rhs_.io_diffCommits_info_106_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_106_vlWen!=rhs_.io_diffCommits_info_106_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_106_vlWen=0x%0h while the rhs_.io_diffCommits_info_106_vlWen=0x%0h",this.io_diffCommits_info_106_vlWen,rhs_.io_diffCommits_info_106_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_107_ldest!=rhs_.io_diffCommits_info_107_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_107_ldest=0x%0h while the rhs_.io_diffCommits_info_107_ldest=0x%0h",this.io_diffCommits_info_107_ldest,rhs_.io_diffCommits_info_107_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_107_pdest!=rhs_.io_diffCommits_info_107_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_107_pdest=0x%0h while the rhs_.io_diffCommits_info_107_pdest=0x%0h",this.io_diffCommits_info_107_pdest,rhs_.io_diffCommits_info_107_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_107_rfWen!=rhs_.io_diffCommits_info_107_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_107_rfWen=0x%0h while the rhs_.io_diffCommits_info_107_rfWen=0x%0h",this.io_diffCommits_info_107_rfWen,rhs_.io_diffCommits_info_107_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_107_fpWen!=rhs_.io_diffCommits_info_107_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_107_fpWen=0x%0h while the rhs_.io_diffCommits_info_107_fpWen=0x%0h",this.io_diffCommits_info_107_fpWen,rhs_.io_diffCommits_info_107_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_107_vecWen!=rhs_.io_diffCommits_info_107_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_107_vecWen=0x%0h while the rhs_.io_diffCommits_info_107_vecWen=0x%0h",this.io_diffCommits_info_107_vecWen,rhs_.io_diffCommits_info_107_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_107_v0Wen!=rhs_.io_diffCommits_info_107_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_107_v0Wen=0x%0h while the rhs_.io_diffCommits_info_107_v0Wen=0x%0h",this.io_diffCommits_info_107_v0Wen,rhs_.io_diffCommits_info_107_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_107_vlWen!=rhs_.io_diffCommits_info_107_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_107_vlWen=0x%0h while the rhs_.io_diffCommits_info_107_vlWen=0x%0h",this.io_diffCommits_info_107_vlWen,rhs_.io_diffCommits_info_107_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_108_ldest!=rhs_.io_diffCommits_info_108_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_108_ldest=0x%0h while the rhs_.io_diffCommits_info_108_ldest=0x%0h",this.io_diffCommits_info_108_ldest,rhs_.io_diffCommits_info_108_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_108_pdest!=rhs_.io_diffCommits_info_108_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_108_pdest=0x%0h while the rhs_.io_diffCommits_info_108_pdest=0x%0h",this.io_diffCommits_info_108_pdest,rhs_.io_diffCommits_info_108_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_108_rfWen!=rhs_.io_diffCommits_info_108_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_108_rfWen=0x%0h while the rhs_.io_diffCommits_info_108_rfWen=0x%0h",this.io_diffCommits_info_108_rfWen,rhs_.io_diffCommits_info_108_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_108_fpWen!=rhs_.io_diffCommits_info_108_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_108_fpWen=0x%0h while the rhs_.io_diffCommits_info_108_fpWen=0x%0h",this.io_diffCommits_info_108_fpWen,rhs_.io_diffCommits_info_108_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_108_vecWen!=rhs_.io_diffCommits_info_108_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_108_vecWen=0x%0h while the rhs_.io_diffCommits_info_108_vecWen=0x%0h",this.io_diffCommits_info_108_vecWen,rhs_.io_diffCommits_info_108_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_108_v0Wen!=rhs_.io_diffCommits_info_108_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_108_v0Wen=0x%0h while the rhs_.io_diffCommits_info_108_v0Wen=0x%0h",this.io_diffCommits_info_108_v0Wen,rhs_.io_diffCommits_info_108_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_108_vlWen!=rhs_.io_diffCommits_info_108_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_108_vlWen=0x%0h while the rhs_.io_diffCommits_info_108_vlWen=0x%0h",this.io_diffCommits_info_108_vlWen,rhs_.io_diffCommits_info_108_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_109_ldest!=rhs_.io_diffCommits_info_109_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_109_ldest=0x%0h while the rhs_.io_diffCommits_info_109_ldest=0x%0h",this.io_diffCommits_info_109_ldest,rhs_.io_diffCommits_info_109_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_109_pdest!=rhs_.io_diffCommits_info_109_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_109_pdest=0x%0h while the rhs_.io_diffCommits_info_109_pdest=0x%0h",this.io_diffCommits_info_109_pdest,rhs_.io_diffCommits_info_109_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_109_rfWen!=rhs_.io_diffCommits_info_109_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_109_rfWen=0x%0h while the rhs_.io_diffCommits_info_109_rfWen=0x%0h",this.io_diffCommits_info_109_rfWen,rhs_.io_diffCommits_info_109_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_109_fpWen!=rhs_.io_diffCommits_info_109_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_109_fpWen=0x%0h while the rhs_.io_diffCommits_info_109_fpWen=0x%0h",this.io_diffCommits_info_109_fpWen,rhs_.io_diffCommits_info_109_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_109_vecWen!=rhs_.io_diffCommits_info_109_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_109_vecWen=0x%0h while the rhs_.io_diffCommits_info_109_vecWen=0x%0h",this.io_diffCommits_info_109_vecWen,rhs_.io_diffCommits_info_109_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_109_v0Wen!=rhs_.io_diffCommits_info_109_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_109_v0Wen=0x%0h while the rhs_.io_diffCommits_info_109_v0Wen=0x%0h",this.io_diffCommits_info_109_v0Wen,rhs_.io_diffCommits_info_109_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_109_vlWen!=rhs_.io_diffCommits_info_109_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_109_vlWen=0x%0h while the rhs_.io_diffCommits_info_109_vlWen=0x%0h",this.io_diffCommits_info_109_vlWen,rhs_.io_diffCommits_info_109_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_110_ldest!=rhs_.io_diffCommits_info_110_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_110_ldest=0x%0h while the rhs_.io_diffCommits_info_110_ldest=0x%0h",this.io_diffCommits_info_110_ldest,rhs_.io_diffCommits_info_110_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_110_pdest!=rhs_.io_diffCommits_info_110_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_110_pdest=0x%0h while the rhs_.io_diffCommits_info_110_pdest=0x%0h",this.io_diffCommits_info_110_pdest,rhs_.io_diffCommits_info_110_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_110_rfWen!=rhs_.io_diffCommits_info_110_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_110_rfWen=0x%0h while the rhs_.io_diffCommits_info_110_rfWen=0x%0h",this.io_diffCommits_info_110_rfWen,rhs_.io_diffCommits_info_110_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_110_fpWen!=rhs_.io_diffCommits_info_110_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_110_fpWen=0x%0h while the rhs_.io_diffCommits_info_110_fpWen=0x%0h",this.io_diffCommits_info_110_fpWen,rhs_.io_diffCommits_info_110_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_110_vecWen!=rhs_.io_diffCommits_info_110_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_110_vecWen=0x%0h while the rhs_.io_diffCommits_info_110_vecWen=0x%0h",this.io_diffCommits_info_110_vecWen,rhs_.io_diffCommits_info_110_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_110_v0Wen!=rhs_.io_diffCommits_info_110_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_110_v0Wen=0x%0h while the rhs_.io_diffCommits_info_110_v0Wen=0x%0h",this.io_diffCommits_info_110_v0Wen,rhs_.io_diffCommits_info_110_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_110_vlWen!=rhs_.io_diffCommits_info_110_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_110_vlWen=0x%0h while the rhs_.io_diffCommits_info_110_vlWen=0x%0h",this.io_diffCommits_info_110_vlWen,rhs_.io_diffCommits_info_110_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_111_ldest!=rhs_.io_diffCommits_info_111_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_111_ldest=0x%0h while the rhs_.io_diffCommits_info_111_ldest=0x%0h",this.io_diffCommits_info_111_ldest,rhs_.io_diffCommits_info_111_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_111_pdest!=rhs_.io_diffCommits_info_111_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_111_pdest=0x%0h while the rhs_.io_diffCommits_info_111_pdest=0x%0h",this.io_diffCommits_info_111_pdest,rhs_.io_diffCommits_info_111_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_111_rfWen!=rhs_.io_diffCommits_info_111_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_111_rfWen=0x%0h while the rhs_.io_diffCommits_info_111_rfWen=0x%0h",this.io_diffCommits_info_111_rfWen,rhs_.io_diffCommits_info_111_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_111_fpWen!=rhs_.io_diffCommits_info_111_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_111_fpWen=0x%0h while the rhs_.io_diffCommits_info_111_fpWen=0x%0h",this.io_diffCommits_info_111_fpWen,rhs_.io_diffCommits_info_111_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_111_vecWen!=rhs_.io_diffCommits_info_111_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_111_vecWen=0x%0h while the rhs_.io_diffCommits_info_111_vecWen=0x%0h",this.io_diffCommits_info_111_vecWen,rhs_.io_diffCommits_info_111_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_111_v0Wen!=rhs_.io_diffCommits_info_111_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_111_v0Wen=0x%0h while the rhs_.io_diffCommits_info_111_v0Wen=0x%0h",this.io_diffCommits_info_111_v0Wen,rhs_.io_diffCommits_info_111_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_111_vlWen!=rhs_.io_diffCommits_info_111_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_111_vlWen=0x%0h while the rhs_.io_diffCommits_info_111_vlWen=0x%0h",this.io_diffCommits_info_111_vlWen,rhs_.io_diffCommits_info_111_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_112_ldest!=rhs_.io_diffCommits_info_112_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_112_ldest=0x%0h while the rhs_.io_diffCommits_info_112_ldest=0x%0h",this.io_diffCommits_info_112_ldest,rhs_.io_diffCommits_info_112_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_112_pdest!=rhs_.io_diffCommits_info_112_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_112_pdest=0x%0h while the rhs_.io_diffCommits_info_112_pdest=0x%0h",this.io_diffCommits_info_112_pdest,rhs_.io_diffCommits_info_112_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_112_rfWen!=rhs_.io_diffCommits_info_112_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_112_rfWen=0x%0h while the rhs_.io_diffCommits_info_112_rfWen=0x%0h",this.io_diffCommits_info_112_rfWen,rhs_.io_diffCommits_info_112_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_112_fpWen!=rhs_.io_diffCommits_info_112_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_112_fpWen=0x%0h while the rhs_.io_diffCommits_info_112_fpWen=0x%0h",this.io_diffCommits_info_112_fpWen,rhs_.io_diffCommits_info_112_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_112_vecWen!=rhs_.io_diffCommits_info_112_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_112_vecWen=0x%0h while the rhs_.io_diffCommits_info_112_vecWen=0x%0h",this.io_diffCommits_info_112_vecWen,rhs_.io_diffCommits_info_112_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_112_v0Wen!=rhs_.io_diffCommits_info_112_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_112_v0Wen=0x%0h while the rhs_.io_diffCommits_info_112_v0Wen=0x%0h",this.io_diffCommits_info_112_v0Wen,rhs_.io_diffCommits_info_112_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_112_vlWen!=rhs_.io_diffCommits_info_112_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_112_vlWen=0x%0h while the rhs_.io_diffCommits_info_112_vlWen=0x%0h",this.io_diffCommits_info_112_vlWen,rhs_.io_diffCommits_info_112_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_113_ldest!=rhs_.io_diffCommits_info_113_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_113_ldest=0x%0h while the rhs_.io_diffCommits_info_113_ldest=0x%0h",this.io_diffCommits_info_113_ldest,rhs_.io_diffCommits_info_113_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_113_pdest!=rhs_.io_diffCommits_info_113_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_113_pdest=0x%0h while the rhs_.io_diffCommits_info_113_pdest=0x%0h",this.io_diffCommits_info_113_pdest,rhs_.io_diffCommits_info_113_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_113_rfWen!=rhs_.io_diffCommits_info_113_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_113_rfWen=0x%0h while the rhs_.io_diffCommits_info_113_rfWen=0x%0h",this.io_diffCommits_info_113_rfWen,rhs_.io_diffCommits_info_113_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_113_fpWen!=rhs_.io_diffCommits_info_113_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_113_fpWen=0x%0h while the rhs_.io_diffCommits_info_113_fpWen=0x%0h",this.io_diffCommits_info_113_fpWen,rhs_.io_diffCommits_info_113_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_113_vecWen!=rhs_.io_diffCommits_info_113_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_113_vecWen=0x%0h while the rhs_.io_diffCommits_info_113_vecWen=0x%0h",this.io_diffCommits_info_113_vecWen,rhs_.io_diffCommits_info_113_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_113_v0Wen!=rhs_.io_diffCommits_info_113_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_113_v0Wen=0x%0h while the rhs_.io_diffCommits_info_113_v0Wen=0x%0h",this.io_diffCommits_info_113_v0Wen,rhs_.io_diffCommits_info_113_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_113_vlWen!=rhs_.io_diffCommits_info_113_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_113_vlWen=0x%0h while the rhs_.io_diffCommits_info_113_vlWen=0x%0h",this.io_diffCommits_info_113_vlWen,rhs_.io_diffCommits_info_113_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_114_ldest!=rhs_.io_diffCommits_info_114_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_114_ldest=0x%0h while the rhs_.io_diffCommits_info_114_ldest=0x%0h",this.io_diffCommits_info_114_ldest,rhs_.io_diffCommits_info_114_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_114_pdest!=rhs_.io_diffCommits_info_114_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_114_pdest=0x%0h while the rhs_.io_diffCommits_info_114_pdest=0x%0h",this.io_diffCommits_info_114_pdest,rhs_.io_diffCommits_info_114_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_114_rfWen!=rhs_.io_diffCommits_info_114_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_114_rfWen=0x%0h while the rhs_.io_diffCommits_info_114_rfWen=0x%0h",this.io_diffCommits_info_114_rfWen,rhs_.io_diffCommits_info_114_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_114_fpWen!=rhs_.io_diffCommits_info_114_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_114_fpWen=0x%0h while the rhs_.io_diffCommits_info_114_fpWen=0x%0h",this.io_diffCommits_info_114_fpWen,rhs_.io_diffCommits_info_114_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_114_vecWen!=rhs_.io_diffCommits_info_114_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_114_vecWen=0x%0h while the rhs_.io_diffCommits_info_114_vecWen=0x%0h",this.io_diffCommits_info_114_vecWen,rhs_.io_diffCommits_info_114_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_114_v0Wen!=rhs_.io_diffCommits_info_114_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_114_v0Wen=0x%0h while the rhs_.io_diffCommits_info_114_v0Wen=0x%0h",this.io_diffCommits_info_114_v0Wen,rhs_.io_diffCommits_info_114_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_114_vlWen!=rhs_.io_diffCommits_info_114_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_114_vlWen=0x%0h while the rhs_.io_diffCommits_info_114_vlWen=0x%0h",this.io_diffCommits_info_114_vlWen,rhs_.io_diffCommits_info_114_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_115_ldest!=rhs_.io_diffCommits_info_115_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_115_ldest=0x%0h while the rhs_.io_diffCommits_info_115_ldest=0x%0h",this.io_diffCommits_info_115_ldest,rhs_.io_diffCommits_info_115_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_115_pdest!=rhs_.io_diffCommits_info_115_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_115_pdest=0x%0h while the rhs_.io_diffCommits_info_115_pdest=0x%0h",this.io_diffCommits_info_115_pdest,rhs_.io_diffCommits_info_115_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_115_rfWen!=rhs_.io_diffCommits_info_115_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_115_rfWen=0x%0h while the rhs_.io_diffCommits_info_115_rfWen=0x%0h",this.io_diffCommits_info_115_rfWen,rhs_.io_diffCommits_info_115_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_115_fpWen!=rhs_.io_diffCommits_info_115_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_115_fpWen=0x%0h while the rhs_.io_diffCommits_info_115_fpWen=0x%0h",this.io_diffCommits_info_115_fpWen,rhs_.io_diffCommits_info_115_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_115_vecWen!=rhs_.io_diffCommits_info_115_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_115_vecWen=0x%0h while the rhs_.io_diffCommits_info_115_vecWen=0x%0h",this.io_diffCommits_info_115_vecWen,rhs_.io_diffCommits_info_115_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_115_v0Wen!=rhs_.io_diffCommits_info_115_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_115_v0Wen=0x%0h while the rhs_.io_diffCommits_info_115_v0Wen=0x%0h",this.io_diffCommits_info_115_v0Wen,rhs_.io_diffCommits_info_115_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_115_vlWen!=rhs_.io_diffCommits_info_115_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_115_vlWen=0x%0h while the rhs_.io_diffCommits_info_115_vlWen=0x%0h",this.io_diffCommits_info_115_vlWen,rhs_.io_diffCommits_info_115_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_116_ldest!=rhs_.io_diffCommits_info_116_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_116_ldest=0x%0h while the rhs_.io_diffCommits_info_116_ldest=0x%0h",this.io_diffCommits_info_116_ldest,rhs_.io_diffCommits_info_116_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_116_pdest!=rhs_.io_diffCommits_info_116_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_116_pdest=0x%0h while the rhs_.io_diffCommits_info_116_pdest=0x%0h",this.io_diffCommits_info_116_pdest,rhs_.io_diffCommits_info_116_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_116_rfWen!=rhs_.io_diffCommits_info_116_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_116_rfWen=0x%0h while the rhs_.io_diffCommits_info_116_rfWen=0x%0h",this.io_diffCommits_info_116_rfWen,rhs_.io_diffCommits_info_116_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_116_fpWen!=rhs_.io_diffCommits_info_116_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_116_fpWen=0x%0h while the rhs_.io_diffCommits_info_116_fpWen=0x%0h",this.io_diffCommits_info_116_fpWen,rhs_.io_diffCommits_info_116_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_116_vecWen!=rhs_.io_diffCommits_info_116_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_116_vecWen=0x%0h while the rhs_.io_diffCommits_info_116_vecWen=0x%0h",this.io_diffCommits_info_116_vecWen,rhs_.io_diffCommits_info_116_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_116_v0Wen!=rhs_.io_diffCommits_info_116_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_116_v0Wen=0x%0h while the rhs_.io_diffCommits_info_116_v0Wen=0x%0h",this.io_diffCommits_info_116_v0Wen,rhs_.io_diffCommits_info_116_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_116_vlWen!=rhs_.io_diffCommits_info_116_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_116_vlWen=0x%0h while the rhs_.io_diffCommits_info_116_vlWen=0x%0h",this.io_diffCommits_info_116_vlWen,rhs_.io_diffCommits_info_116_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_117_ldest!=rhs_.io_diffCommits_info_117_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_117_ldest=0x%0h while the rhs_.io_diffCommits_info_117_ldest=0x%0h",this.io_diffCommits_info_117_ldest,rhs_.io_diffCommits_info_117_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_117_pdest!=rhs_.io_diffCommits_info_117_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_117_pdest=0x%0h while the rhs_.io_diffCommits_info_117_pdest=0x%0h",this.io_diffCommits_info_117_pdest,rhs_.io_diffCommits_info_117_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_117_rfWen!=rhs_.io_diffCommits_info_117_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_117_rfWen=0x%0h while the rhs_.io_diffCommits_info_117_rfWen=0x%0h",this.io_diffCommits_info_117_rfWen,rhs_.io_diffCommits_info_117_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_117_fpWen!=rhs_.io_diffCommits_info_117_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_117_fpWen=0x%0h while the rhs_.io_diffCommits_info_117_fpWen=0x%0h",this.io_diffCommits_info_117_fpWen,rhs_.io_diffCommits_info_117_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_117_vecWen!=rhs_.io_diffCommits_info_117_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_117_vecWen=0x%0h while the rhs_.io_diffCommits_info_117_vecWen=0x%0h",this.io_diffCommits_info_117_vecWen,rhs_.io_diffCommits_info_117_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_117_v0Wen!=rhs_.io_diffCommits_info_117_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_117_v0Wen=0x%0h while the rhs_.io_diffCommits_info_117_v0Wen=0x%0h",this.io_diffCommits_info_117_v0Wen,rhs_.io_diffCommits_info_117_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_117_vlWen!=rhs_.io_diffCommits_info_117_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_117_vlWen=0x%0h while the rhs_.io_diffCommits_info_117_vlWen=0x%0h",this.io_diffCommits_info_117_vlWen,rhs_.io_diffCommits_info_117_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_118_ldest!=rhs_.io_diffCommits_info_118_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_118_ldest=0x%0h while the rhs_.io_diffCommits_info_118_ldest=0x%0h",this.io_diffCommits_info_118_ldest,rhs_.io_diffCommits_info_118_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_118_pdest!=rhs_.io_diffCommits_info_118_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_118_pdest=0x%0h while the rhs_.io_diffCommits_info_118_pdest=0x%0h",this.io_diffCommits_info_118_pdest,rhs_.io_diffCommits_info_118_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_118_rfWen!=rhs_.io_diffCommits_info_118_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_118_rfWen=0x%0h while the rhs_.io_diffCommits_info_118_rfWen=0x%0h",this.io_diffCommits_info_118_rfWen,rhs_.io_diffCommits_info_118_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_118_fpWen!=rhs_.io_diffCommits_info_118_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_118_fpWen=0x%0h while the rhs_.io_diffCommits_info_118_fpWen=0x%0h",this.io_diffCommits_info_118_fpWen,rhs_.io_diffCommits_info_118_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_118_vecWen!=rhs_.io_diffCommits_info_118_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_118_vecWen=0x%0h while the rhs_.io_diffCommits_info_118_vecWen=0x%0h",this.io_diffCommits_info_118_vecWen,rhs_.io_diffCommits_info_118_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_118_v0Wen!=rhs_.io_diffCommits_info_118_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_118_v0Wen=0x%0h while the rhs_.io_diffCommits_info_118_v0Wen=0x%0h",this.io_diffCommits_info_118_v0Wen,rhs_.io_diffCommits_info_118_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_118_vlWen!=rhs_.io_diffCommits_info_118_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_118_vlWen=0x%0h while the rhs_.io_diffCommits_info_118_vlWen=0x%0h",this.io_diffCommits_info_118_vlWen,rhs_.io_diffCommits_info_118_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_119_ldest!=rhs_.io_diffCommits_info_119_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_119_ldest=0x%0h while the rhs_.io_diffCommits_info_119_ldest=0x%0h",this.io_diffCommits_info_119_ldest,rhs_.io_diffCommits_info_119_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_119_pdest!=rhs_.io_diffCommits_info_119_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_119_pdest=0x%0h while the rhs_.io_diffCommits_info_119_pdest=0x%0h",this.io_diffCommits_info_119_pdest,rhs_.io_diffCommits_info_119_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_119_rfWen!=rhs_.io_diffCommits_info_119_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_119_rfWen=0x%0h while the rhs_.io_diffCommits_info_119_rfWen=0x%0h",this.io_diffCommits_info_119_rfWen,rhs_.io_diffCommits_info_119_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_119_fpWen!=rhs_.io_diffCommits_info_119_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_119_fpWen=0x%0h while the rhs_.io_diffCommits_info_119_fpWen=0x%0h",this.io_diffCommits_info_119_fpWen,rhs_.io_diffCommits_info_119_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_119_vecWen!=rhs_.io_diffCommits_info_119_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_119_vecWen=0x%0h while the rhs_.io_diffCommits_info_119_vecWen=0x%0h",this.io_diffCommits_info_119_vecWen,rhs_.io_diffCommits_info_119_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_119_v0Wen!=rhs_.io_diffCommits_info_119_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_119_v0Wen=0x%0h while the rhs_.io_diffCommits_info_119_v0Wen=0x%0h",this.io_diffCommits_info_119_v0Wen,rhs_.io_diffCommits_info_119_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_119_vlWen!=rhs_.io_diffCommits_info_119_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_119_vlWen=0x%0h while the rhs_.io_diffCommits_info_119_vlWen=0x%0h",this.io_diffCommits_info_119_vlWen,rhs_.io_diffCommits_info_119_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_120_ldest!=rhs_.io_diffCommits_info_120_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_120_ldest=0x%0h while the rhs_.io_diffCommits_info_120_ldest=0x%0h",this.io_diffCommits_info_120_ldest,rhs_.io_diffCommits_info_120_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_120_pdest!=rhs_.io_diffCommits_info_120_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_120_pdest=0x%0h while the rhs_.io_diffCommits_info_120_pdest=0x%0h",this.io_diffCommits_info_120_pdest,rhs_.io_diffCommits_info_120_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_120_rfWen!=rhs_.io_diffCommits_info_120_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_120_rfWen=0x%0h while the rhs_.io_diffCommits_info_120_rfWen=0x%0h",this.io_diffCommits_info_120_rfWen,rhs_.io_diffCommits_info_120_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_120_fpWen!=rhs_.io_diffCommits_info_120_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_120_fpWen=0x%0h while the rhs_.io_diffCommits_info_120_fpWen=0x%0h",this.io_diffCommits_info_120_fpWen,rhs_.io_diffCommits_info_120_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_120_vecWen!=rhs_.io_diffCommits_info_120_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_120_vecWen=0x%0h while the rhs_.io_diffCommits_info_120_vecWen=0x%0h",this.io_diffCommits_info_120_vecWen,rhs_.io_diffCommits_info_120_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_120_v0Wen!=rhs_.io_diffCommits_info_120_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_120_v0Wen=0x%0h while the rhs_.io_diffCommits_info_120_v0Wen=0x%0h",this.io_diffCommits_info_120_v0Wen,rhs_.io_diffCommits_info_120_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_120_vlWen!=rhs_.io_diffCommits_info_120_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_120_vlWen=0x%0h while the rhs_.io_diffCommits_info_120_vlWen=0x%0h",this.io_diffCommits_info_120_vlWen,rhs_.io_diffCommits_info_120_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_121_ldest!=rhs_.io_diffCommits_info_121_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_121_ldest=0x%0h while the rhs_.io_diffCommits_info_121_ldest=0x%0h",this.io_diffCommits_info_121_ldest,rhs_.io_diffCommits_info_121_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_121_pdest!=rhs_.io_diffCommits_info_121_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_121_pdest=0x%0h while the rhs_.io_diffCommits_info_121_pdest=0x%0h",this.io_diffCommits_info_121_pdest,rhs_.io_diffCommits_info_121_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_121_rfWen!=rhs_.io_diffCommits_info_121_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_121_rfWen=0x%0h while the rhs_.io_diffCommits_info_121_rfWen=0x%0h",this.io_diffCommits_info_121_rfWen,rhs_.io_diffCommits_info_121_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_121_fpWen!=rhs_.io_diffCommits_info_121_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_121_fpWen=0x%0h while the rhs_.io_diffCommits_info_121_fpWen=0x%0h",this.io_diffCommits_info_121_fpWen,rhs_.io_diffCommits_info_121_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_121_vecWen!=rhs_.io_diffCommits_info_121_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_121_vecWen=0x%0h while the rhs_.io_diffCommits_info_121_vecWen=0x%0h",this.io_diffCommits_info_121_vecWen,rhs_.io_diffCommits_info_121_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_121_v0Wen!=rhs_.io_diffCommits_info_121_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_121_v0Wen=0x%0h while the rhs_.io_diffCommits_info_121_v0Wen=0x%0h",this.io_diffCommits_info_121_v0Wen,rhs_.io_diffCommits_info_121_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_121_vlWen!=rhs_.io_diffCommits_info_121_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_121_vlWen=0x%0h while the rhs_.io_diffCommits_info_121_vlWen=0x%0h",this.io_diffCommits_info_121_vlWen,rhs_.io_diffCommits_info_121_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_122_ldest!=rhs_.io_diffCommits_info_122_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_122_ldest=0x%0h while the rhs_.io_diffCommits_info_122_ldest=0x%0h",this.io_diffCommits_info_122_ldest,rhs_.io_diffCommits_info_122_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_122_pdest!=rhs_.io_diffCommits_info_122_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_122_pdest=0x%0h while the rhs_.io_diffCommits_info_122_pdest=0x%0h",this.io_diffCommits_info_122_pdest,rhs_.io_diffCommits_info_122_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_122_rfWen!=rhs_.io_diffCommits_info_122_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_122_rfWen=0x%0h while the rhs_.io_diffCommits_info_122_rfWen=0x%0h",this.io_diffCommits_info_122_rfWen,rhs_.io_diffCommits_info_122_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_122_fpWen!=rhs_.io_diffCommits_info_122_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_122_fpWen=0x%0h while the rhs_.io_diffCommits_info_122_fpWen=0x%0h",this.io_diffCommits_info_122_fpWen,rhs_.io_diffCommits_info_122_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_122_vecWen!=rhs_.io_diffCommits_info_122_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_122_vecWen=0x%0h while the rhs_.io_diffCommits_info_122_vecWen=0x%0h",this.io_diffCommits_info_122_vecWen,rhs_.io_diffCommits_info_122_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_122_v0Wen!=rhs_.io_diffCommits_info_122_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_122_v0Wen=0x%0h while the rhs_.io_diffCommits_info_122_v0Wen=0x%0h",this.io_diffCommits_info_122_v0Wen,rhs_.io_diffCommits_info_122_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_122_vlWen!=rhs_.io_diffCommits_info_122_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_122_vlWen=0x%0h while the rhs_.io_diffCommits_info_122_vlWen=0x%0h",this.io_diffCommits_info_122_vlWen,rhs_.io_diffCommits_info_122_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_123_ldest!=rhs_.io_diffCommits_info_123_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_123_ldest=0x%0h while the rhs_.io_diffCommits_info_123_ldest=0x%0h",this.io_diffCommits_info_123_ldest,rhs_.io_diffCommits_info_123_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_123_pdest!=rhs_.io_diffCommits_info_123_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_123_pdest=0x%0h while the rhs_.io_diffCommits_info_123_pdest=0x%0h",this.io_diffCommits_info_123_pdest,rhs_.io_diffCommits_info_123_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_123_rfWen!=rhs_.io_diffCommits_info_123_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_123_rfWen=0x%0h while the rhs_.io_diffCommits_info_123_rfWen=0x%0h",this.io_diffCommits_info_123_rfWen,rhs_.io_diffCommits_info_123_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_123_fpWen!=rhs_.io_diffCommits_info_123_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_123_fpWen=0x%0h while the rhs_.io_diffCommits_info_123_fpWen=0x%0h",this.io_diffCommits_info_123_fpWen,rhs_.io_diffCommits_info_123_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_123_vecWen!=rhs_.io_diffCommits_info_123_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_123_vecWen=0x%0h while the rhs_.io_diffCommits_info_123_vecWen=0x%0h",this.io_diffCommits_info_123_vecWen,rhs_.io_diffCommits_info_123_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_123_v0Wen!=rhs_.io_diffCommits_info_123_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_123_v0Wen=0x%0h while the rhs_.io_diffCommits_info_123_v0Wen=0x%0h",this.io_diffCommits_info_123_v0Wen,rhs_.io_diffCommits_info_123_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_123_vlWen!=rhs_.io_diffCommits_info_123_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_123_vlWen=0x%0h while the rhs_.io_diffCommits_info_123_vlWen=0x%0h",this.io_diffCommits_info_123_vlWen,rhs_.io_diffCommits_info_123_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_124_ldest!=rhs_.io_diffCommits_info_124_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_124_ldest=0x%0h while the rhs_.io_diffCommits_info_124_ldest=0x%0h",this.io_diffCommits_info_124_ldest,rhs_.io_diffCommits_info_124_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_124_pdest!=rhs_.io_diffCommits_info_124_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_124_pdest=0x%0h while the rhs_.io_diffCommits_info_124_pdest=0x%0h",this.io_diffCommits_info_124_pdest,rhs_.io_diffCommits_info_124_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_124_rfWen!=rhs_.io_diffCommits_info_124_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_124_rfWen=0x%0h while the rhs_.io_diffCommits_info_124_rfWen=0x%0h",this.io_diffCommits_info_124_rfWen,rhs_.io_diffCommits_info_124_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_124_fpWen!=rhs_.io_diffCommits_info_124_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_124_fpWen=0x%0h while the rhs_.io_diffCommits_info_124_fpWen=0x%0h",this.io_diffCommits_info_124_fpWen,rhs_.io_diffCommits_info_124_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_124_vecWen!=rhs_.io_diffCommits_info_124_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_124_vecWen=0x%0h while the rhs_.io_diffCommits_info_124_vecWen=0x%0h",this.io_diffCommits_info_124_vecWen,rhs_.io_diffCommits_info_124_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_124_v0Wen!=rhs_.io_diffCommits_info_124_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_124_v0Wen=0x%0h while the rhs_.io_diffCommits_info_124_v0Wen=0x%0h",this.io_diffCommits_info_124_v0Wen,rhs_.io_diffCommits_info_124_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_124_vlWen!=rhs_.io_diffCommits_info_124_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_124_vlWen=0x%0h while the rhs_.io_diffCommits_info_124_vlWen=0x%0h",this.io_diffCommits_info_124_vlWen,rhs_.io_diffCommits_info_124_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_125_ldest!=rhs_.io_diffCommits_info_125_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_125_ldest=0x%0h while the rhs_.io_diffCommits_info_125_ldest=0x%0h",this.io_diffCommits_info_125_ldest,rhs_.io_diffCommits_info_125_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_125_pdest!=rhs_.io_diffCommits_info_125_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_125_pdest=0x%0h while the rhs_.io_diffCommits_info_125_pdest=0x%0h",this.io_diffCommits_info_125_pdest,rhs_.io_diffCommits_info_125_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_125_rfWen!=rhs_.io_diffCommits_info_125_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_125_rfWen=0x%0h while the rhs_.io_diffCommits_info_125_rfWen=0x%0h",this.io_diffCommits_info_125_rfWen,rhs_.io_diffCommits_info_125_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_125_fpWen!=rhs_.io_diffCommits_info_125_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_125_fpWen=0x%0h while the rhs_.io_diffCommits_info_125_fpWen=0x%0h",this.io_diffCommits_info_125_fpWen,rhs_.io_diffCommits_info_125_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_125_vecWen!=rhs_.io_diffCommits_info_125_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_125_vecWen=0x%0h while the rhs_.io_diffCommits_info_125_vecWen=0x%0h",this.io_diffCommits_info_125_vecWen,rhs_.io_diffCommits_info_125_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_125_v0Wen!=rhs_.io_diffCommits_info_125_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_125_v0Wen=0x%0h while the rhs_.io_diffCommits_info_125_v0Wen=0x%0h",this.io_diffCommits_info_125_v0Wen,rhs_.io_diffCommits_info_125_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_125_vlWen!=rhs_.io_diffCommits_info_125_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_125_vlWen=0x%0h while the rhs_.io_diffCommits_info_125_vlWen=0x%0h",this.io_diffCommits_info_125_vlWen,rhs_.io_diffCommits_info_125_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_126_ldest!=rhs_.io_diffCommits_info_126_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_126_ldest=0x%0h while the rhs_.io_diffCommits_info_126_ldest=0x%0h",this.io_diffCommits_info_126_ldest,rhs_.io_diffCommits_info_126_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_126_pdest!=rhs_.io_diffCommits_info_126_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_126_pdest=0x%0h while the rhs_.io_diffCommits_info_126_pdest=0x%0h",this.io_diffCommits_info_126_pdest,rhs_.io_diffCommits_info_126_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_126_rfWen!=rhs_.io_diffCommits_info_126_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_126_rfWen=0x%0h while the rhs_.io_diffCommits_info_126_rfWen=0x%0h",this.io_diffCommits_info_126_rfWen,rhs_.io_diffCommits_info_126_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_126_fpWen!=rhs_.io_diffCommits_info_126_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_126_fpWen=0x%0h while the rhs_.io_diffCommits_info_126_fpWen=0x%0h",this.io_diffCommits_info_126_fpWen,rhs_.io_diffCommits_info_126_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_126_vecWen!=rhs_.io_diffCommits_info_126_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_126_vecWen=0x%0h while the rhs_.io_diffCommits_info_126_vecWen=0x%0h",this.io_diffCommits_info_126_vecWen,rhs_.io_diffCommits_info_126_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_126_v0Wen!=rhs_.io_diffCommits_info_126_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_126_v0Wen=0x%0h while the rhs_.io_diffCommits_info_126_v0Wen=0x%0h",this.io_diffCommits_info_126_v0Wen,rhs_.io_diffCommits_info_126_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_126_vlWen!=rhs_.io_diffCommits_info_126_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_126_vlWen=0x%0h while the rhs_.io_diffCommits_info_126_vlWen=0x%0h",this.io_diffCommits_info_126_vlWen,rhs_.io_diffCommits_info_126_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_127_ldest!=rhs_.io_diffCommits_info_127_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_127_ldest=0x%0h while the rhs_.io_diffCommits_info_127_ldest=0x%0h",this.io_diffCommits_info_127_ldest,rhs_.io_diffCommits_info_127_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_127_pdest!=rhs_.io_diffCommits_info_127_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_127_pdest=0x%0h while the rhs_.io_diffCommits_info_127_pdest=0x%0h",this.io_diffCommits_info_127_pdest,rhs_.io_diffCommits_info_127_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_127_rfWen!=rhs_.io_diffCommits_info_127_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_127_rfWen=0x%0h while the rhs_.io_diffCommits_info_127_rfWen=0x%0h",this.io_diffCommits_info_127_rfWen,rhs_.io_diffCommits_info_127_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_127_fpWen!=rhs_.io_diffCommits_info_127_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_127_fpWen=0x%0h while the rhs_.io_diffCommits_info_127_fpWen=0x%0h",this.io_diffCommits_info_127_fpWen,rhs_.io_diffCommits_info_127_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_127_vecWen!=rhs_.io_diffCommits_info_127_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_127_vecWen=0x%0h while the rhs_.io_diffCommits_info_127_vecWen=0x%0h",this.io_diffCommits_info_127_vecWen,rhs_.io_diffCommits_info_127_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_127_v0Wen!=rhs_.io_diffCommits_info_127_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_127_v0Wen=0x%0h while the rhs_.io_diffCommits_info_127_v0Wen=0x%0h",this.io_diffCommits_info_127_v0Wen,rhs_.io_diffCommits_info_127_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_127_vlWen!=rhs_.io_diffCommits_info_127_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_127_vlWen=0x%0h while the rhs_.io_diffCommits_info_127_vlWen=0x%0h",this.io_diffCommits_info_127_vlWen,rhs_.io_diffCommits_info_127_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_128_ldest!=rhs_.io_diffCommits_info_128_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_128_ldest=0x%0h while the rhs_.io_diffCommits_info_128_ldest=0x%0h",this.io_diffCommits_info_128_ldest,rhs_.io_diffCommits_info_128_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_128_pdest!=rhs_.io_diffCommits_info_128_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_128_pdest=0x%0h while the rhs_.io_diffCommits_info_128_pdest=0x%0h",this.io_diffCommits_info_128_pdest,rhs_.io_diffCommits_info_128_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_128_rfWen!=rhs_.io_diffCommits_info_128_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_128_rfWen=0x%0h while the rhs_.io_diffCommits_info_128_rfWen=0x%0h",this.io_diffCommits_info_128_rfWen,rhs_.io_diffCommits_info_128_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_128_fpWen!=rhs_.io_diffCommits_info_128_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_128_fpWen=0x%0h while the rhs_.io_diffCommits_info_128_fpWen=0x%0h",this.io_diffCommits_info_128_fpWen,rhs_.io_diffCommits_info_128_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_128_vecWen!=rhs_.io_diffCommits_info_128_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_128_vecWen=0x%0h while the rhs_.io_diffCommits_info_128_vecWen=0x%0h",this.io_diffCommits_info_128_vecWen,rhs_.io_diffCommits_info_128_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_128_v0Wen!=rhs_.io_diffCommits_info_128_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_128_v0Wen=0x%0h while the rhs_.io_diffCommits_info_128_v0Wen=0x%0h",this.io_diffCommits_info_128_v0Wen,rhs_.io_diffCommits_info_128_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_128_vlWen!=rhs_.io_diffCommits_info_128_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_128_vlWen=0x%0h while the rhs_.io_diffCommits_info_128_vlWen=0x%0h",this.io_diffCommits_info_128_vlWen,rhs_.io_diffCommits_info_128_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_129_ldest!=rhs_.io_diffCommits_info_129_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_129_ldest=0x%0h while the rhs_.io_diffCommits_info_129_ldest=0x%0h",this.io_diffCommits_info_129_ldest,rhs_.io_diffCommits_info_129_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_129_pdest!=rhs_.io_diffCommits_info_129_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_129_pdest=0x%0h while the rhs_.io_diffCommits_info_129_pdest=0x%0h",this.io_diffCommits_info_129_pdest,rhs_.io_diffCommits_info_129_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_129_rfWen!=rhs_.io_diffCommits_info_129_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_129_rfWen=0x%0h while the rhs_.io_diffCommits_info_129_rfWen=0x%0h",this.io_diffCommits_info_129_rfWen,rhs_.io_diffCommits_info_129_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_129_fpWen!=rhs_.io_diffCommits_info_129_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_129_fpWen=0x%0h while the rhs_.io_diffCommits_info_129_fpWen=0x%0h",this.io_diffCommits_info_129_fpWen,rhs_.io_diffCommits_info_129_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_129_vecWen!=rhs_.io_diffCommits_info_129_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_129_vecWen=0x%0h while the rhs_.io_diffCommits_info_129_vecWen=0x%0h",this.io_diffCommits_info_129_vecWen,rhs_.io_diffCommits_info_129_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_129_v0Wen!=rhs_.io_diffCommits_info_129_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_129_v0Wen=0x%0h while the rhs_.io_diffCommits_info_129_v0Wen=0x%0h",this.io_diffCommits_info_129_v0Wen,rhs_.io_diffCommits_info_129_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_129_vlWen!=rhs_.io_diffCommits_info_129_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_129_vlWen=0x%0h while the rhs_.io_diffCommits_info_129_vlWen=0x%0h",this.io_diffCommits_info_129_vlWen,rhs_.io_diffCommits_info_129_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_130_ldest!=rhs_.io_diffCommits_info_130_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_130_ldest=0x%0h while the rhs_.io_diffCommits_info_130_ldest=0x%0h",this.io_diffCommits_info_130_ldest,rhs_.io_diffCommits_info_130_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_130_pdest!=rhs_.io_diffCommits_info_130_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_130_pdest=0x%0h while the rhs_.io_diffCommits_info_130_pdest=0x%0h",this.io_diffCommits_info_130_pdest,rhs_.io_diffCommits_info_130_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_130_rfWen!=rhs_.io_diffCommits_info_130_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_130_rfWen=0x%0h while the rhs_.io_diffCommits_info_130_rfWen=0x%0h",this.io_diffCommits_info_130_rfWen,rhs_.io_diffCommits_info_130_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_130_fpWen!=rhs_.io_diffCommits_info_130_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_130_fpWen=0x%0h while the rhs_.io_diffCommits_info_130_fpWen=0x%0h",this.io_diffCommits_info_130_fpWen,rhs_.io_diffCommits_info_130_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_130_vecWen!=rhs_.io_diffCommits_info_130_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_130_vecWen=0x%0h while the rhs_.io_diffCommits_info_130_vecWen=0x%0h",this.io_diffCommits_info_130_vecWen,rhs_.io_diffCommits_info_130_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_130_v0Wen!=rhs_.io_diffCommits_info_130_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_130_v0Wen=0x%0h while the rhs_.io_diffCommits_info_130_v0Wen=0x%0h",this.io_diffCommits_info_130_v0Wen,rhs_.io_diffCommits_info_130_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_130_vlWen!=rhs_.io_diffCommits_info_130_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_130_vlWen=0x%0h while the rhs_.io_diffCommits_info_130_vlWen=0x%0h",this.io_diffCommits_info_130_vlWen,rhs_.io_diffCommits_info_130_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_131_ldest!=rhs_.io_diffCommits_info_131_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_131_ldest=0x%0h while the rhs_.io_diffCommits_info_131_ldest=0x%0h",this.io_diffCommits_info_131_ldest,rhs_.io_diffCommits_info_131_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_131_pdest!=rhs_.io_diffCommits_info_131_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_131_pdest=0x%0h while the rhs_.io_diffCommits_info_131_pdest=0x%0h",this.io_diffCommits_info_131_pdest,rhs_.io_diffCommits_info_131_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_131_rfWen!=rhs_.io_diffCommits_info_131_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_131_rfWen=0x%0h while the rhs_.io_diffCommits_info_131_rfWen=0x%0h",this.io_diffCommits_info_131_rfWen,rhs_.io_diffCommits_info_131_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_131_fpWen!=rhs_.io_diffCommits_info_131_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_131_fpWen=0x%0h while the rhs_.io_diffCommits_info_131_fpWen=0x%0h",this.io_diffCommits_info_131_fpWen,rhs_.io_diffCommits_info_131_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_131_vecWen!=rhs_.io_diffCommits_info_131_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_131_vecWen=0x%0h while the rhs_.io_diffCommits_info_131_vecWen=0x%0h",this.io_diffCommits_info_131_vecWen,rhs_.io_diffCommits_info_131_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_131_v0Wen!=rhs_.io_diffCommits_info_131_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_131_v0Wen=0x%0h while the rhs_.io_diffCommits_info_131_v0Wen=0x%0h",this.io_diffCommits_info_131_v0Wen,rhs_.io_diffCommits_info_131_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_131_vlWen!=rhs_.io_diffCommits_info_131_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_131_vlWen=0x%0h while the rhs_.io_diffCommits_info_131_vlWen=0x%0h",this.io_diffCommits_info_131_vlWen,rhs_.io_diffCommits_info_131_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_132_ldest!=rhs_.io_diffCommits_info_132_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_132_ldest=0x%0h while the rhs_.io_diffCommits_info_132_ldest=0x%0h",this.io_diffCommits_info_132_ldest,rhs_.io_diffCommits_info_132_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_132_pdest!=rhs_.io_diffCommits_info_132_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_132_pdest=0x%0h while the rhs_.io_diffCommits_info_132_pdest=0x%0h",this.io_diffCommits_info_132_pdest,rhs_.io_diffCommits_info_132_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_132_rfWen!=rhs_.io_diffCommits_info_132_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_132_rfWen=0x%0h while the rhs_.io_diffCommits_info_132_rfWen=0x%0h",this.io_diffCommits_info_132_rfWen,rhs_.io_diffCommits_info_132_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_132_fpWen!=rhs_.io_diffCommits_info_132_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_132_fpWen=0x%0h while the rhs_.io_diffCommits_info_132_fpWen=0x%0h",this.io_diffCommits_info_132_fpWen,rhs_.io_diffCommits_info_132_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_132_vecWen!=rhs_.io_diffCommits_info_132_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_132_vecWen=0x%0h while the rhs_.io_diffCommits_info_132_vecWen=0x%0h",this.io_diffCommits_info_132_vecWen,rhs_.io_diffCommits_info_132_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_132_v0Wen!=rhs_.io_diffCommits_info_132_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_132_v0Wen=0x%0h while the rhs_.io_diffCommits_info_132_v0Wen=0x%0h",this.io_diffCommits_info_132_v0Wen,rhs_.io_diffCommits_info_132_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_132_vlWen!=rhs_.io_diffCommits_info_132_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_132_vlWen=0x%0h while the rhs_.io_diffCommits_info_132_vlWen=0x%0h",this.io_diffCommits_info_132_vlWen,rhs_.io_diffCommits_info_132_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_133_ldest!=rhs_.io_diffCommits_info_133_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_133_ldest=0x%0h while the rhs_.io_diffCommits_info_133_ldest=0x%0h",this.io_diffCommits_info_133_ldest,rhs_.io_diffCommits_info_133_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_133_pdest!=rhs_.io_diffCommits_info_133_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_133_pdest=0x%0h while the rhs_.io_diffCommits_info_133_pdest=0x%0h",this.io_diffCommits_info_133_pdest,rhs_.io_diffCommits_info_133_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_133_rfWen!=rhs_.io_diffCommits_info_133_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_133_rfWen=0x%0h while the rhs_.io_diffCommits_info_133_rfWen=0x%0h",this.io_diffCommits_info_133_rfWen,rhs_.io_diffCommits_info_133_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_133_fpWen!=rhs_.io_diffCommits_info_133_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_133_fpWen=0x%0h while the rhs_.io_diffCommits_info_133_fpWen=0x%0h",this.io_diffCommits_info_133_fpWen,rhs_.io_diffCommits_info_133_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_133_vecWen!=rhs_.io_diffCommits_info_133_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_133_vecWen=0x%0h while the rhs_.io_diffCommits_info_133_vecWen=0x%0h",this.io_diffCommits_info_133_vecWen,rhs_.io_diffCommits_info_133_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_133_v0Wen!=rhs_.io_diffCommits_info_133_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_133_v0Wen=0x%0h while the rhs_.io_diffCommits_info_133_v0Wen=0x%0h",this.io_diffCommits_info_133_v0Wen,rhs_.io_diffCommits_info_133_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_133_vlWen!=rhs_.io_diffCommits_info_133_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_133_vlWen=0x%0h while the rhs_.io_diffCommits_info_133_vlWen=0x%0h",this.io_diffCommits_info_133_vlWen,rhs_.io_diffCommits_info_133_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_134_ldest!=rhs_.io_diffCommits_info_134_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_134_ldest=0x%0h while the rhs_.io_diffCommits_info_134_ldest=0x%0h",this.io_diffCommits_info_134_ldest,rhs_.io_diffCommits_info_134_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_134_pdest!=rhs_.io_diffCommits_info_134_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_134_pdest=0x%0h while the rhs_.io_diffCommits_info_134_pdest=0x%0h",this.io_diffCommits_info_134_pdest,rhs_.io_diffCommits_info_134_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_134_rfWen!=rhs_.io_diffCommits_info_134_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_134_rfWen=0x%0h while the rhs_.io_diffCommits_info_134_rfWen=0x%0h",this.io_diffCommits_info_134_rfWen,rhs_.io_diffCommits_info_134_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_134_fpWen!=rhs_.io_diffCommits_info_134_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_134_fpWen=0x%0h while the rhs_.io_diffCommits_info_134_fpWen=0x%0h",this.io_diffCommits_info_134_fpWen,rhs_.io_diffCommits_info_134_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_134_vecWen!=rhs_.io_diffCommits_info_134_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_134_vecWen=0x%0h while the rhs_.io_diffCommits_info_134_vecWen=0x%0h",this.io_diffCommits_info_134_vecWen,rhs_.io_diffCommits_info_134_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_134_v0Wen!=rhs_.io_diffCommits_info_134_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_134_v0Wen=0x%0h while the rhs_.io_diffCommits_info_134_v0Wen=0x%0h",this.io_diffCommits_info_134_v0Wen,rhs_.io_diffCommits_info_134_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_134_vlWen!=rhs_.io_diffCommits_info_134_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_134_vlWen=0x%0h while the rhs_.io_diffCommits_info_134_vlWen=0x%0h",this.io_diffCommits_info_134_vlWen,rhs_.io_diffCommits_info_134_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_135_ldest!=rhs_.io_diffCommits_info_135_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_135_ldest=0x%0h while the rhs_.io_diffCommits_info_135_ldest=0x%0h",this.io_diffCommits_info_135_ldest,rhs_.io_diffCommits_info_135_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_135_pdest!=rhs_.io_diffCommits_info_135_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_135_pdest=0x%0h while the rhs_.io_diffCommits_info_135_pdest=0x%0h",this.io_diffCommits_info_135_pdest,rhs_.io_diffCommits_info_135_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_135_rfWen!=rhs_.io_diffCommits_info_135_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_135_rfWen=0x%0h while the rhs_.io_diffCommits_info_135_rfWen=0x%0h",this.io_diffCommits_info_135_rfWen,rhs_.io_diffCommits_info_135_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_135_fpWen!=rhs_.io_diffCommits_info_135_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_135_fpWen=0x%0h while the rhs_.io_diffCommits_info_135_fpWen=0x%0h",this.io_diffCommits_info_135_fpWen,rhs_.io_diffCommits_info_135_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_135_vecWen!=rhs_.io_diffCommits_info_135_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_135_vecWen=0x%0h while the rhs_.io_diffCommits_info_135_vecWen=0x%0h",this.io_diffCommits_info_135_vecWen,rhs_.io_diffCommits_info_135_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_135_v0Wen!=rhs_.io_diffCommits_info_135_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_135_v0Wen=0x%0h while the rhs_.io_diffCommits_info_135_v0Wen=0x%0h",this.io_diffCommits_info_135_v0Wen,rhs_.io_diffCommits_info_135_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_135_vlWen!=rhs_.io_diffCommits_info_135_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_135_vlWen=0x%0h while the rhs_.io_diffCommits_info_135_vlWen=0x%0h",this.io_diffCommits_info_135_vlWen,rhs_.io_diffCommits_info_135_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_136_ldest!=rhs_.io_diffCommits_info_136_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_136_ldest=0x%0h while the rhs_.io_diffCommits_info_136_ldest=0x%0h",this.io_diffCommits_info_136_ldest,rhs_.io_diffCommits_info_136_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_136_pdest!=rhs_.io_diffCommits_info_136_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_136_pdest=0x%0h while the rhs_.io_diffCommits_info_136_pdest=0x%0h",this.io_diffCommits_info_136_pdest,rhs_.io_diffCommits_info_136_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_136_rfWen!=rhs_.io_diffCommits_info_136_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_136_rfWen=0x%0h while the rhs_.io_diffCommits_info_136_rfWen=0x%0h",this.io_diffCommits_info_136_rfWen,rhs_.io_diffCommits_info_136_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_136_fpWen!=rhs_.io_diffCommits_info_136_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_136_fpWen=0x%0h while the rhs_.io_diffCommits_info_136_fpWen=0x%0h",this.io_diffCommits_info_136_fpWen,rhs_.io_diffCommits_info_136_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_136_vecWen!=rhs_.io_diffCommits_info_136_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_136_vecWen=0x%0h while the rhs_.io_diffCommits_info_136_vecWen=0x%0h",this.io_diffCommits_info_136_vecWen,rhs_.io_diffCommits_info_136_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_136_v0Wen!=rhs_.io_diffCommits_info_136_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_136_v0Wen=0x%0h while the rhs_.io_diffCommits_info_136_v0Wen=0x%0h",this.io_diffCommits_info_136_v0Wen,rhs_.io_diffCommits_info_136_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_136_vlWen!=rhs_.io_diffCommits_info_136_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_136_vlWen=0x%0h while the rhs_.io_diffCommits_info_136_vlWen=0x%0h",this.io_diffCommits_info_136_vlWen,rhs_.io_diffCommits_info_136_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_137_ldest!=rhs_.io_diffCommits_info_137_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_137_ldest=0x%0h while the rhs_.io_diffCommits_info_137_ldest=0x%0h",this.io_diffCommits_info_137_ldest,rhs_.io_diffCommits_info_137_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_137_pdest!=rhs_.io_diffCommits_info_137_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_137_pdest=0x%0h while the rhs_.io_diffCommits_info_137_pdest=0x%0h",this.io_diffCommits_info_137_pdest,rhs_.io_diffCommits_info_137_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_137_rfWen!=rhs_.io_diffCommits_info_137_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_137_rfWen=0x%0h while the rhs_.io_diffCommits_info_137_rfWen=0x%0h",this.io_diffCommits_info_137_rfWen,rhs_.io_diffCommits_info_137_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_137_fpWen!=rhs_.io_diffCommits_info_137_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_137_fpWen=0x%0h while the rhs_.io_diffCommits_info_137_fpWen=0x%0h",this.io_diffCommits_info_137_fpWen,rhs_.io_diffCommits_info_137_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_137_vecWen!=rhs_.io_diffCommits_info_137_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_137_vecWen=0x%0h while the rhs_.io_diffCommits_info_137_vecWen=0x%0h",this.io_diffCommits_info_137_vecWen,rhs_.io_diffCommits_info_137_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_137_v0Wen!=rhs_.io_diffCommits_info_137_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_137_v0Wen=0x%0h while the rhs_.io_diffCommits_info_137_v0Wen=0x%0h",this.io_diffCommits_info_137_v0Wen,rhs_.io_diffCommits_info_137_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_137_vlWen!=rhs_.io_diffCommits_info_137_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_137_vlWen=0x%0h while the rhs_.io_diffCommits_info_137_vlWen=0x%0h",this.io_diffCommits_info_137_vlWen,rhs_.io_diffCommits_info_137_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_138_ldest!=rhs_.io_diffCommits_info_138_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_138_ldest=0x%0h while the rhs_.io_diffCommits_info_138_ldest=0x%0h",this.io_diffCommits_info_138_ldest,rhs_.io_diffCommits_info_138_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_138_pdest!=rhs_.io_diffCommits_info_138_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_138_pdest=0x%0h while the rhs_.io_diffCommits_info_138_pdest=0x%0h",this.io_diffCommits_info_138_pdest,rhs_.io_diffCommits_info_138_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_138_rfWen!=rhs_.io_diffCommits_info_138_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_138_rfWen=0x%0h while the rhs_.io_diffCommits_info_138_rfWen=0x%0h",this.io_diffCommits_info_138_rfWen,rhs_.io_diffCommits_info_138_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_138_fpWen!=rhs_.io_diffCommits_info_138_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_138_fpWen=0x%0h while the rhs_.io_diffCommits_info_138_fpWen=0x%0h",this.io_diffCommits_info_138_fpWen,rhs_.io_diffCommits_info_138_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_138_vecWen!=rhs_.io_diffCommits_info_138_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_138_vecWen=0x%0h while the rhs_.io_diffCommits_info_138_vecWen=0x%0h",this.io_diffCommits_info_138_vecWen,rhs_.io_diffCommits_info_138_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_138_v0Wen!=rhs_.io_diffCommits_info_138_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_138_v0Wen=0x%0h while the rhs_.io_diffCommits_info_138_v0Wen=0x%0h",this.io_diffCommits_info_138_v0Wen,rhs_.io_diffCommits_info_138_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_138_vlWen!=rhs_.io_diffCommits_info_138_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_138_vlWen=0x%0h while the rhs_.io_diffCommits_info_138_vlWen=0x%0h",this.io_diffCommits_info_138_vlWen,rhs_.io_diffCommits_info_138_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_139_ldest!=rhs_.io_diffCommits_info_139_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_139_ldest=0x%0h while the rhs_.io_diffCommits_info_139_ldest=0x%0h",this.io_diffCommits_info_139_ldest,rhs_.io_diffCommits_info_139_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_139_pdest!=rhs_.io_diffCommits_info_139_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_139_pdest=0x%0h while the rhs_.io_diffCommits_info_139_pdest=0x%0h",this.io_diffCommits_info_139_pdest,rhs_.io_diffCommits_info_139_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_139_rfWen!=rhs_.io_diffCommits_info_139_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_139_rfWen=0x%0h while the rhs_.io_diffCommits_info_139_rfWen=0x%0h",this.io_diffCommits_info_139_rfWen,rhs_.io_diffCommits_info_139_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_139_fpWen!=rhs_.io_diffCommits_info_139_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_139_fpWen=0x%0h while the rhs_.io_diffCommits_info_139_fpWen=0x%0h",this.io_diffCommits_info_139_fpWen,rhs_.io_diffCommits_info_139_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_139_vecWen!=rhs_.io_diffCommits_info_139_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_139_vecWen=0x%0h while the rhs_.io_diffCommits_info_139_vecWen=0x%0h",this.io_diffCommits_info_139_vecWen,rhs_.io_diffCommits_info_139_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_139_v0Wen!=rhs_.io_diffCommits_info_139_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_139_v0Wen=0x%0h while the rhs_.io_diffCommits_info_139_v0Wen=0x%0h",this.io_diffCommits_info_139_v0Wen,rhs_.io_diffCommits_info_139_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_139_vlWen!=rhs_.io_diffCommits_info_139_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_139_vlWen=0x%0h while the rhs_.io_diffCommits_info_139_vlWen=0x%0h",this.io_diffCommits_info_139_vlWen,rhs_.io_diffCommits_info_139_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_140_ldest!=rhs_.io_diffCommits_info_140_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_140_ldest=0x%0h while the rhs_.io_diffCommits_info_140_ldest=0x%0h",this.io_diffCommits_info_140_ldest,rhs_.io_diffCommits_info_140_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_140_pdest!=rhs_.io_diffCommits_info_140_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_140_pdest=0x%0h while the rhs_.io_diffCommits_info_140_pdest=0x%0h",this.io_diffCommits_info_140_pdest,rhs_.io_diffCommits_info_140_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_140_rfWen!=rhs_.io_diffCommits_info_140_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_140_rfWen=0x%0h while the rhs_.io_diffCommits_info_140_rfWen=0x%0h",this.io_diffCommits_info_140_rfWen,rhs_.io_diffCommits_info_140_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_140_fpWen!=rhs_.io_diffCommits_info_140_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_140_fpWen=0x%0h while the rhs_.io_diffCommits_info_140_fpWen=0x%0h",this.io_diffCommits_info_140_fpWen,rhs_.io_diffCommits_info_140_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_140_vecWen!=rhs_.io_diffCommits_info_140_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_140_vecWen=0x%0h while the rhs_.io_diffCommits_info_140_vecWen=0x%0h",this.io_diffCommits_info_140_vecWen,rhs_.io_diffCommits_info_140_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_140_v0Wen!=rhs_.io_diffCommits_info_140_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_140_v0Wen=0x%0h while the rhs_.io_diffCommits_info_140_v0Wen=0x%0h",this.io_diffCommits_info_140_v0Wen,rhs_.io_diffCommits_info_140_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_140_vlWen!=rhs_.io_diffCommits_info_140_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_140_vlWen=0x%0h while the rhs_.io_diffCommits_info_140_vlWen=0x%0h",this.io_diffCommits_info_140_vlWen,rhs_.io_diffCommits_info_140_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_141_ldest!=rhs_.io_diffCommits_info_141_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_141_ldest=0x%0h while the rhs_.io_diffCommits_info_141_ldest=0x%0h",this.io_diffCommits_info_141_ldest,rhs_.io_diffCommits_info_141_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_141_pdest!=rhs_.io_diffCommits_info_141_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_141_pdest=0x%0h while the rhs_.io_diffCommits_info_141_pdest=0x%0h",this.io_diffCommits_info_141_pdest,rhs_.io_diffCommits_info_141_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_141_rfWen!=rhs_.io_diffCommits_info_141_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_141_rfWen=0x%0h while the rhs_.io_diffCommits_info_141_rfWen=0x%0h",this.io_diffCommits_info_141_rfWen,rhs_.io_diffCommits_info_141_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_141_fpWen!=rhs_.io_diffCommits_info_141_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_141_fpWen=0x%0h while the rhs_.io_diffCommits_info_141_fpWen=0x%0h",this.io_diffCommits_info_141_fpWen,rhs_.io_diffCommits_info_141_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_141_vecWen!=rhs_.io_diffCommits_info_141_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_141_vecWen=0x%0h while the rhs_.io_diffCommits_info_141_vecWen=0x%0h",this.io_diffCommits_info_141_vecWen,rhs_.io_diffCommits_info_141_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_141_v0Wen!=rhs_.io_diffCommits_info_141_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_141_v0Wen=0x%0h while the rhs_.io_diffCommits_info_141_v0Wen=0x%0h",this.io_diffCommits_info_141_v0Wen,rhs_.io_diffCommits_info_141_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_141_vlWen!=rhs_.io_diffCommits_info_141_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_141_vlWen=0x%0h while the rhs_.io_diffCommits_info_141_vlWen=0x%0h",this.io_diffCommits_info_141_vlWen,rhs_.io_diffCommits_info_141_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_142_ldest!=rhs_.io_diffCommits_info_142_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_142_ldest=0x%0h while the rhs_.io_diffCommits_info_142_ldest=0x%0h",this.io_diffCommits_info_142_ldest,rhs_.io_diffCommits_info_142_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_142_pdest!=rhs_.io_diffCommits_info_142_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_142_pdest=0x%0h while the rhs_.io_diffCommits_info_142_pdest=0x%0h",this.io_diffCommits_info_142_pdest,rhs_.io_diffCommits_info_142_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_142_rfWen!=rhs_.io_diffCommits_info_142_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_142_rfWen=0x%0h while the rhs_.io_diffCommits_info_142_rfWen=0x%0h",this.io_diffCommits_info_142_rfWen,rhs_.io_diffCommits_info_142_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_142_fpWen!=rhs_.io_diffCommits_info_142_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_142_fpWen=0x%0h while the rhs_.io_diffCommits_info_142_fpWen=0x%0h",this.io_diffCommits_info_142_fpWen,rhs_.io_diffCommits_info_142_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_142_vecWen!=rhs_.io_diffCommits_info_142_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_142_vecWen=0x%0h while the rhs_.io_diffCommits_info_142_vecWen=0x%0h",this.io_diffCommits_info_142_vecWen,rhs_.io_diffCommits_info_142_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_142_v0Wen!=rhs_.io_diffCommits_info_142_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_142_v0Wen=0x%0h while the rhs_.io_diffCommits_info_142_v0Wen=0x%0h",this.io_diffCommits_info_142_v0Wen,rhs_.io_diffCommits_info_142_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_142_vlWen!=rhs_.io_diffCommits_info_142_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_142_vlWen=0x%0h while the rhs_.io_diffCommits_info_142_vlWen=0x%0h",this.io_diffCommits_info_142_vlWen,rhs_.io_diffCommits_info_142_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_143_ldest!=rhs_.io_diffCommits_info_143_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_143_ldest=0x%0h while the rhs_.io_diffCommits_info_143_ldest=0x%0h",this.io_diffCommits_info_143_ldest,rhs_.io_diffCommits_info_143_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_143_pdest!=rhs_.io_diffCommits_info_143_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_143_pdest=0x%0h while the rhs_.io_diffCommits_info_143_pdest=0x%0h",this.io_diffCommits_info_143_pdest,rhs_.io_diffCommits_info_143_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_143_rfWen!=rhs_.io_diffCommits_info_143_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_143_rfWen=0x%0h while the rhs_.io_diffCommits_info_143_rfWen=0x%0h",this.io_diffCommits_info_143_rfWen,rhs_.io_diffCommits_info_143_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_143_fpWen!=rhs_.io_diffCommits_info_143_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_143_fpWen=0x%0h while the rhs_.io_diffCommits_info_143_fpWen=0x%0h",this.io_diffCommits_info_143_fpWen,rhs_.io_diffCommits_info_143_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_143_vecWen!=rhs_.io_diffCommits_info_143_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_143_vecWen=0x%0h while the rhs_.io_diffCommits_info_143_vecWen=0x%0h",this.io_diffCommits_info_143_vecWen,rhs_.io_diffCommits_info_143_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_143_v0Wen!=rhs_.io_diffCommits_info_143_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_143_v0Wen=0x%0h while the rhs_.io_diffCommits_info_143_v0Wen=0x%0h",this.io_diffCommits_info_143_v0Wen,rhs_.io_diffCommits_info_143_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_143_vlWen!=rhs_.io_diffCommits_info_143_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_143_vlWen=0x%0h while the rhs_.io_diffCommits_info_143_vlWen=0x%0h",this.io_diffCommits_info_143_vlWen,rhs_.io_diffCommits_info_143_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_144_ldest!=rhs_.io_diffCommits_info_144_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_144_ldest=0x%0h while the rhs_.io_diffCommits_info_144_ldest=0x%0h",this.io_diffCommits_info_144_ldest,rhs_.io_diffCommits_info_144_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_144_pdest!=rhs_.io_diffCommits_info_144_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_144_pdest=0x%0h while the rhs_.io_diffCommits_info_144_pdest=0x%0h",this.io_diffCommits_info_144_pdest,rhs_.io_diffCommits_info_144_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_144_rfWen!=rhs_.io_diffCommits_info_144_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_144_rfWen=0x%0h while the rhs_.io_diffCommits_info_144_rfWen=0x%0h",this.io_diffCommits_info_144_rfWen,rhs_.io_diffCommits_info_144_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_144_fpWen!=rhs_.io_diffCommits_info_144_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_144_fpWen=0x%0h while the rhs_.io_diffCommits_info_144_fpWen=0x%0h",this.io_diffCommits_info_144_fpWen,rhs_.io_diffCommits_info_144_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_144_vecWen!=rhs_.io_diffCommits_info_144_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_144_vecWen=0x%0h while the rhs_.io_diffCommits_info_144_vecWen=0x%0h",this.io_diffCommits_info_144_vecWen,rhs_.io_diffCommits_info_144_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_144_v0Wen!=rhs_.io_diffCommits_info_144_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_144_v0Wen=0x%0h while the rhs_.io_diffCommits_info_144_v0Wen=0x%0h",this.io_diffCommits_info_144_v0Wen,rhs_.io_diffCommits_info_144_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_144_vlWen!=rhs_.io_diffCommits_info_144_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_144_vlWen=0x%0h while the rhs_.io_diffCommits_info_144_vlWen=0x%0h",this.io_diffCommits_info_144_vlWen,rhs_.io_diffCommits_info_144_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_145_ldest!=rhs_.io_diffCommits_info_145_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_145_ldest=0x%0h while the rhs_.io_diffCommits_info_145_ldest=0x%0h",this.io_diffCommits_info_145_ldest,rhs_.io_diffCommits_info_145_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_145_pdest!=rhs_.io_diffCommits_info_145_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_145_pdest=0x%0h while the rhs_.io_diffCommits_info_145_pdest=0x%0h",this.io_diffCommits_info_145_pdest,rhs_.io_diffCommits_info_145_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_145_rfWen!=rhs_.io_diffCommits_info_145_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_145_rfWen=0x%0h while the rhs_.io_diffCommits_info_145_rfWen=0x%0h",this.io_diffCommits_info_145_rfWen,rhs_.io_diffCommits_info_145_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_145_fpWen!=rhs_.io_diffCommits_info_145_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_145_fpWen=0x%0h while the rhs_.io_diffCommits_info_145_fpWen=0x%0h",this.io_diffCommits_info_145_fpWen,rhs_.io_diffCommits_info_145_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_145_vecWen!=rhs_.io_diffCommits_info_145_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_145_vecWen=0x%0h while the rhs_.io_diffCommits_info_145_vecWen=0x%0h",this.io_diffCommits_info_145_vecWen,rhs_.io_diffCommits_info_145_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_145_v0Wen!=rhs_.io_diffCommits_info_145_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_145_v0Wen=0x%0h while the rhs_.io_diffCommits_info_145_v0Wen=0x%0h",this.io_diffCommits_info_145_v0Wen,rhs_.io_diffCommits_info_145_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_145_vlWen!=rhs_.io_diffCommits_info_145_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_145_vlWen=0x%0h while the rhs_.io_diffCommits_info_145_vlWen=0x%0h",this.io_diffCommits_info_145_vlWen,rhs_.io_diffCommits_info_145_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_146_ldest!=rhs_.io_diffCommits_info_146_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_146_ldest=0x%0h while the rhs_.io_diffCommits_info_146_ldest=0x%0h",this.io_diffCommits_info_146_ldest,rhs_.io_diffCommits_info_146_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_146_pdest!=rhs_.io_diffCommits_info_146_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_146_pdest=0x%0h while the rhs_.io_diffCommits_info_146_pdest=0x%0h",this.io_diffCommits_info_146_pdest,rhs_.io_diffCommits_info_146_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_146_rfWen!=rhs_.io_diffCommits_info_146_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_146_rfWen=0x%0h while the rhs_.io_diffCommits_info_146_rfWen=0x%0h",this.io_diffCommits_info_146_rfWen,rhs_.io_diffCommits_info_146_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_146_fpWen!=rhs_.io_diffCommits_info_146_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_146_fpWen=0x%0h while the rhs_.io_diffCommits_info_146_fpWen=0x%0h",this.io_diffCommits_info_146_fpWen,rhs_.io_diffCommits_info_146_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_146_vecWen!=rhs_.io_diffCommits_info_146_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_146_vecWen=0x%0h while the rhs_.io_diffCommits_info_146_vecWen=0x%0h",this.io_diffCommits_info_146_vecWen,rhs_.io_diffCommits_info_146_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_146_v0Wen!=rhs_.io_diffCommits_info_146_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_146_v0Wen=0x%0h while the rhs_.io_diffCommits_info_146_v0Wen=0x%0h",this.io_diffCommits_info_146_v0Wen,rhs_.io_diffCommits_info_146_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_146_vlWen!=rhs_.io_diffCommits_info_146_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_146_vlWen=0x%0h while the rhs_.io_diffCommits_info_146_vlWen=0x%0h",this.io_diffCommits_info_146_vlWen,rhs_.io_diffCommits_info_146_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_147_ldest!=rhs_.io_diffCommits_info_147_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_147_ldest=0x%0h while the rhs_.io_diffCommits_info_147_ldest=0x%0h",this.io_diffCommits_info_147_ldest,rhs_.io_diffCommits_info_147_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_147_pdest!=rhs_.io_diffCommits_info_147_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_147_pdest=0x%0h while the rhs_.io_diffCommits_info_147_pdest=0x%0h",this.io_diffCommits_info_147_pdest,rhs_.io_diffCommits_info_147_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_147_rfWen!=rhs_.io_diffCommits_info_147_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_147_rfWen=0x%0h while the rhs_.io_diffCommits_info_147_rfWen=0x%0h",this.io_diffCommits_info_147_rfWen,rhs_.io_diffCommits_info_147_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_147_fpWen!=rhs_.io_diffCommits_info_147_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_147_fpWen=0x%0h while the rhs_.io_diffCommits_info_147_fpWen=0x%0h",this.io_diffCommits_info_147_fpWen,rhs_.io_diffCommits_info_147_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_147_vecWen!=rhs_.io_diffCommits_info_147_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_147_vecWen=0x%0h while the rhs_.io_diffCommits_info_147_vecWen=0x%0h",this.io_diffCommits_info_147_vecWen,rhs_.io_diffCommits_info_147_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_147_v0Wen!=rhs_.io_diffCommits_info_147_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_147_v0Wen=0x%0h while the rhs_.io_diffCommits_info_147_v0Wen=0x%0h",this.io_diffCommits_info_147_v0Wen,rhs_.io_diffCommits_info_147_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_147_vlWen!=rhs_.io_diffCommits_info_147_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_147_vlWen=0x%0h while the rhs_.io_diffCommits_info_147_vlWen=0x%0h",this.io_diffCommits_info_147_vlWen,rhs_.io_diffCommits_info_147_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_148_ldest!=rhs_.io_diffCommits_info_148_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_148_ldest=0x%0h while the rhs_.io_diffCommits_info_148_ldest=0x%0h",this.io_diffCommits_info_148_ldest,rhs_.io_diffCommits_info_148_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_148_pdest!=rhs_.io_diffCommits_info_148_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_148_pdest=0x%0h while the rhs_.io_diffCommits_info_148_pdest=0x%0h",this.io_diffCommits_info_148_pdest,rhs_.io_diffCommits_info_148_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_148_rfWen!=rhs_.io_diffCommits_info_148_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_148_rfWen=0x%0h while the rhs_.io_diffCommits_info_148_rfWen=0x%0h",this.io_diffCommits_info_148_rfWen,rhs_.io_diffCommits_info_148_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_148_fpWen!=rhs_.io_diffCommits_info_148_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_148_fpWen=0x%0h while the rhs_.io_diffCommits_info_148_fpWen=0x%0h",this.io_diffCommits_info_148_fpWen,rhs_.io_diffCommits_info_148_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_148_vecWen!=rhs_.io_diffCommits_info_148_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_148_vecWen=0x%0h while the rhs_.io_diffCommits_info_148_vecWen=0x%0h",this.io_diffCommits_info_148_vecWen,rhs_.io_diffCommits_info_148_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_148_v0Wen!=rhs_.io_diffCommits_info_148_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_148_v0Wen=0x%0h while the rhs_.io_diffCommits_info_148_v0Wen=0x%0h",this.io_diffCommits_info_148_v0Wen,rhs_.io_diffCommits_info_148_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_148_vlWen!=rhs_.io_diffCommits_info_148_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_148_vlWen=0x%0h while the rhs_.io_diffCommits_info_148_vlWen=0x%0h",this.io_diffCommits_info_148_vlWen,rhs_.io_diffCommits_info_148_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_149_ldest!=rhs_.io_diffCommits_info_149_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_149_ldest=0x%0h while the rhs_.io_diffCommits_info_149_ldest=0x%0h",this.io_diffCommits_info_149_ldest,rhs_.io_diffCommits_info_149_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_149_pdest!=rhs_.io_diffCommits_info_149_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_149_pdest=0x%0h while the rhs_.io_diffCommits_info_149_pdest=0x%0h",this.io_diffCommits_info_149_pdest,rhs_.io_diffCommits_info_149_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_149_rfWen!=rhs_.io_diffCommits_info_149_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_149_rfWen=0x%0h while the rhs_.io_diffCommits_info_149_rfWen=0x%0h",this.io_diffCommits_info_149_rfWen,rhs_.io_diffCommits_info_149_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_149_fpWen!=rhs_.io_diffCommits_info_149_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_149_fpWen=0x%0h while the rhs_.io_diffCommits_info_149_fpWen=0x%0h",this.io_diffCommits_info_149_fpWen,rhs_.io_diffCommits_info_149_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_149_vecWen!=rhs_.io_diffCommits_info_149_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_149_vecWen=0x%0h while the rhs_.io_diffCommits_info_149_vecWen=0x%0h",this.io_diffCommits_info_149_vecWen,rhs_.io_diffCommits_info_149_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_149_v0Wen!=rhs_.io_diffCommits_info_149_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_149_v0Wen=0x%0h while the rhs_.io_diffCommits_info_149_v0Wen=0x%0h",this.io_diffCommits_info_149_v0Wen,rhs_.io_diffCommits_info_149_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_149_vlWen!=rhs_.io_diffCommits_info_149_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_149_vlWen=0x%0h while the rhs_.io_diffCommits_info_149_vlWen=0x%0h",this.io_diffCommits_info_149_vlWen,rhs_.io_diffCommits_info_149_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_150_ldest!=rhs_.io_diffCommits_info_150_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_150_ldest=0x%0h while the rhs_.io_diffCommits_info_150_ldest=0x%0h",this.io_diffCommits_info_150_ldest,rhs_.io_diffCommits_info_150_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_150_pdest!=rhs_.io_diffCommits_info_150_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_150_pdest=0x%0h while the rhs_.io_diffCommits_info_150_pdest=0x%0h",this.io_diffCommits_info_150_pdest,rhs_.io_diffCommits_info_150_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_150_rfWen!=rhs_.io_diffCommits_info_150_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_150_rfWen=0x%0h while the rhs_.io_diffCommits_info_150_rfWen=0x%0h",this.io_diffCommits_info_150_rfWen,rhs_.io_diffCommits_info_150_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_150_fpWen!=rhs_.io_diffCommits_info_150_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_150_fpWen=0x%0h while the rhs_.io_diffCommits_info_150_fpWen=0x%0h",this.io_diffCommits_info_150_fpWen,rhs_.io_diffCommits_info_150_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_150_vecWen!=rhs_.io_diffCommits_info_150_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_150_vecWen=0x%0h while the rhs_.io_diffCommits_info_150_vecWen=0x%0h",this.io_diffCommits_info_150_vecWen,rhs_.io_diffCommits_info_150_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_150_v0Wen!=rhs_.io_diffCommits_info_150_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_150_v0Wen=0x%0h while the rhs_.io_diffCommits_info_150_v0Wen=0x%0h",this.io_diffCommits_info_150_v0Wen,rhs_.io_diffCommits_info_150_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_150_vlWen!=rhs_.io_diffCommits_info_150_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_150_vlWen=0x%0h while the rhs_.io_diffCommits_info_150_vlWen=0x%0h",this.io_diffCommits_info_150_vlWen,rhs_.io_diffCommits_info_150_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_151_ldest!=rhs_.io_diffCommits_info_151_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_151_ldest=0x%0h while the rhs_.io_diffCommits_info_151_ldest=0x%0h",this.io_diffCommits_info_151_ldest,rhs_.io_diffCommits_info_151_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_151_pdest!=rhs_.io_diffCommits_info_151_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_151_pdest=0x%0h while the rhs_.io_diffCommits_info_151_pdest=0x%0h",this.io_diffCommits_info_151_pdest,rhs_.io_diffCommits_info_151_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_151_rfWen!=rhs_.io_diffCommits_info_151_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_151_rfWen=0x%0h while the rhs_.io_diffCommits_info_151_rfWen=0x%0h",this.io_diffCommits_info_151_rfWen,rhs_.io_diffCommits_info_151_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_151_fpWen!=rhs_.io_diffCommits_info_151_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_151_fpWen=0x%0h while the rhs_.io_diffCommits_info_151_fpWen=0x%0h",this.io_diffCommits_info_151_fpWen,rhs_.io_diffCommits_info_151_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_151_vecWen!=rhs_.io_diffCommits_info_151_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_151_vecWen=0x%0h while the rhs_.io_diffCommits_info_151_vecWen=0x%0h",this.io_diffCommits_info_151_vecWen,rhs_.io_diffCommits_info_151_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_151_v0Wen!=rhs_.io_diffCommits_info_151_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_151_v0Wen=0x%0h while the rhs_.io_diffCommits_info_151_v0Wen=0x%0h",this.io_diffCommits_info_151_v0Wen,rhs_.io_diffCommits_info_151_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_151_vlWen!=rhs_.io_diffCommits_info_151_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_151_vlWen=0x%0h while the rhs_.io_diffCommits_info_151_vlWen=0x%0h",this.io_diffCommits_info_151_vlWen,rhs_.io_diffCommits_info_151_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_152_ldest!=rhs_.io_diffCommits_info_152_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_152_ldest=0x%0h while the rhs_.io_diffCommits_info_152_ldest=0x%0h",this.io_diffCommits_info_152_ldest,rhs_.io_diffCommits_info_152_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_152_pdest!=rhs_.io_diffCommits_info_152_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_152_pdest=0x%0h while the rhs_.io_diffCommits_info_152_pdest=0x%0h",this.io_diffCommits_info_152_pdest,rhs_.io_diffCommits_info_152_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_152_rfWen!=rhs_.io_diffCommits_info_152_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_152_rfWen=0x%0h while the rhs_.io_diffCommits_info_152_rfWen=0x%0h",this.io_diffCommits_info_152_rfWen,rhs_.io_diffCommits_info_152_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_152_fpWen!=rhs_.io_diffCommits_info_152_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_152_fpWen=0x%0h while the rhs_.io_diffCommits_info_152_fpWen=0x%0h",this.io_diffCommits_info_152_fpWen,rhs_.io_diffCommits_info_152_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_152_vecWen!=rhs_.io_diffCommits_info_152_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_152_vecWen=0x%0h while the rhs_.io_diffCommits_info_152_vecWen=0x%0h",this.io_diffCommits_info_152_vecWen,rhs_.io_diffCommits_info_152_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_152_v0Wen!=rhs_.io_diffCommits_info_152_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_152_v0Wen=0x%0h while the rhs_.io_diffCommits_info_152_v0Wen=0x%0h",this.io_diffCommits_info_152_v0Wen,rhs_.io_diffCommits_info_152_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_152_vlWen!=rhs_.io_diffCommits_info_152_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_152_vlWen=0x%0h while the rhs_.io_diffCommits_info_152_vlWen=0x%0h",this.io_diffCommits_info_152_vlWen,rhs_.io_diffCommits_info_152_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_153_ldest!=rhs_.io_diffCommits_info_153_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_153_ldest=0x%0h while the rhs_.io_diffCommits_info_153_ldest=0x%0h",this.io_diffCommits_info_153_ldest,rhs_.io_diffCommits_info_153_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_153_pdest!=rhs_.io_diffCommits_info_153_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_153_pdest=0x%0h while the rhs_.io_diffCommits_info_153_pdest=0x%0h",this.io_diffCommits_info_153_pdest,rhs_.io_diffCommits_info_153_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_153_rfWen!=rhs_.io_diffCommits_info_153_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_153_rfWen=0x%0h while the rhs_.io_diffCommits_info_153_rfWen=0x%0h",this.io_diffCommits_info_153_rfWen,rhs_.io_diffCommits_info_153_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_153_fpWen!=rhs_.io_diffCommits_info_153_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_153_fpWen=0x%0h while the rhs_.io_diffCommits_info_153_fpWen=0x%0h",this.io_diffCommits_info_153_fpWen,rhs_.io_diffCommits_info_153_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_153_vecWen!=rhs_.io_diffCommits_info_153_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_153_vecWen=0x%0h while the rhs_.io_diffCommits_info_153_vecWen=0x%0h",this.io_diffCommits_info_153_vecWen,rhs_.io_diffCommits_info_153_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_153_v0Wen!=rhs_.io_diffCommits_info_153_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_153_v0Wen=0x%0h while the rhs_.io_diffCommits_info_153_v0Wen=0x%0h",this.io_diffCommits_info_153_v0Wen,rhs_.io_diffCommits_info_153_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_153_vlWen!=rhs_.io_diffCommits_info_153_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_153_vlWen=0x%0h while the rhs_.io_diffCommits_info_153_vlWen=0x%0h",this.io_diffCommits_info_153_vlWen,rhs_.io_diffCommits_info_153_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_154_ldest!=rhs_.io_diffCommits_info_154_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_154_ldest=0x%0h while the rhs_.io_diffCommits_info_154_ldest=0x%0h",this.io_diffCommits_info_154_ldest,rhs_.io_diffCommits_info_154_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_154_pdest!=rhs_.io_diffCommits_info_154_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_154_pdest=0x%0h while the rhs_.io_diffCommits_info_154_pdest=0x%0h",this.io_diffCommits_info_154_pdest,rhs_.io_diffCommits_info_154_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_154_rfWen!=rhs_.io_diffCommits_info_154_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_154_rfWen=0x%0h while the rhs_.io_diffCommits_info_154_rfWen=0x%0h",this.io_diffCommits_info_154_rfWen,rhs_.io_diffCommits_info_154_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_154_fpWen!=rhs_.io_diffCommits_info_154_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_154_fpWen=0x%0h while the rhs_.io_diffCommits_info_154_fpWen=0x%0h",this.io_diffCommits_info_154_fpWen,rhs_.io_diffCommits_info_154_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_154_vecWen!=rhs_.io_diffCommits_info_154_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_154_vecWen=0x%0h while the rhs_.io_diffCommits_info_154_vecWen=0x%0h",this.io_diffCommits_info_154_vecWen,rhs_.io_diffCommits_info_154_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_154_v0Wen!=rhs_.io_diffCommits_info_154_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_154_v0Wen=0x%0h while the rhs_.io_diffCommits_info_154_v0Wen=0x%0h",this.io_diffCommits_info_154_v0Wen,rhs_.io_diffCommits_info_154_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_154_vlWen!=rhs_.io_diffCommits_info_154_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_154_vlWen=0x%0h while the rhs_.io_diffCommits_info_154_vlWen=0x%0h",this.io_diffCommits_info_154_vlWen,rhs_.io_diffCommits_info_154_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_155_ldest!=rhs_.io_diffCommits_info_155_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_155_ldest=0x%0h while the rhs_.io_diffCommits_info_155_ldest=0x%0h",this.io_diffCommits_info_155_ldest,rhs_.io_diffCommits_info_155_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_155_pdest!=rhs_.io_diffCommits_info_155_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_155_pdest=0x%0h while the rhs_.io_diffCommits_info_155_pdest=0x%0h",this.io_diffCommits_info_155_pdest,rhs_.io_diffCommits_info_155_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_155_rfWen!=rhs_.io_diffCommits_info_155_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_155_rfWen=0x%0h while the rhs_.io_diffCommits_info_155_rfWen=0x%0h",this.io_diffCommits_info_155_rfWen,rhs_.io_diffCommits_info_155_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_155_fpWen!=rhs_.io_diffCommits_info_155_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_155_fpWen=0x%0h while the rhs_.io_diffCommits_info_155_fpWen=0x%0h",this.io_diffCommits_info_155_fpWen,rhs_.io_diffCommits_info_155_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_155_vecWen!=rhs_.io_diffCommits_info_155_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_155_vecWen=0x%0h while the rhs_.io_diffCommits_info_155_vecWen=0x%0h",this.io_diffCommits_info_155_vecWen,rhs_.io_diffCommits_info_155_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_155_v0Wen!=rhs_.io_diffCommits_info_155_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_155_v0Wen=0x%0h while the rhs_.io_diffCommits_info_155_v0Wen=0x%0h",this.io_diffCommits_info_155_v0Wen,rhs_.io_diffCommits_info_155_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_155_vlWen!=rhs_.io_diffCommits_info_155_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_155_vlWen=0x%0h while the rhs_.io_diffCommits_info_155_vlWen=0x%0h",this.io_diffCommits_info_155_vlWen,rhs_.io_diffCommits_info_155_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_156_ldest!=rhs_.io_diffCommits_info_156_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_156_ldest=0x%0h while the rhs_.io_diffCommits_info_156_ldest=0x%0h",this.io_diffCommits_info_156_ldest,rhs_.io_diffCommits_info_156_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_156_pdest!=rhs_.io_diffCommits_info_156_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_156_pdest=0x%0h while the rhs_.io_diffCommits_info_156_pdest=0x%0h",this.io_diffCommits_info_156_pdest,rhs_.io_diffCommits_info_156_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_156_rfWen!=rhs_.io_diffCommits_info_156_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_156_rfWen=0x%0h while the rhs_.io_diffCommits_info_156_rfWen=0x%0h",this.io_diffCommits_info_156_rfWen,rhs_.io_diffCommits_info_156_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_156_fpWen!=rhs_.io_diffCommits_info_156_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_156_fpWen=0x%0h while the rhs_.io_diffCommits_info_156_fpWen=0x%0h",this.io_diffCommits_info_156_fpWen,rhs_.io_diffCommits_info_156_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_156_vecWen!=rhs_.io_diffCommits_info_156_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_156_vecWen=0x%0h while the rhs_.io_diffCommits_info_156_vecWen=0x%0h",this.io_diffCommits_info_156_vecWen,rhs_.io_diffCommits_info_156_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_156_v0Wen!=rhs_.io_diffCommits_info_156_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_156_v0Wen=0x%0h while the rhs_.io_diffCommits_info_156_v0Wen=0x%0h",this.io_diffCommits_info_156_v0Wen,rhs_.io_diffCommits_info_156_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_156_vlWen!=rhs_.io_diffCommits_info_156_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_156_vlWen=0x%0h while the rhs_.io_diffCommits_info_156_vlWen=0x%0h",this.io_diffCommits_info_156_vlWen,rhs_.io_diffCommits_info_156_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_157_ldest!=rhs_.io_diffCommits_info_157_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_157_ldest=0x%0h while the rhs_.io_diffCommits_info_157_ldest=0x%0h",this.io_diffCommits_info_157_ldest,rhs_.io_diffCommits_info_157_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_157_pdest!=rhs_.io_diffCommits_info_157_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_157_pdest=0x%0h while the rhs_.io_diffCommits_info_157_pdest=0x%0h",this.io_diffCommits_info_157_pdest,rhs_.io_diffCommits_info_157_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_157_rfWen!=rhs_.io_diffCommits_info_157_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_157_rfWen=0x%0h while the rhs_.io_diffCommits_info_157_rfWen=0x%0h",this.io_diffCommits_info_157_rfWen,rhs_.io_diffCommits_info_157_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_157_fpWen!=rhs_.io_diffCommits_info_157_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_157_fpWen=0x%0h while the rhs_.io_diffCommits_info_157_fpWen=0x%0h",this.io_diffCommits_info_157_fpWen,rhs_.io_diffCommits_info_157_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_157_vecWen!=rhs_.io_diffCommits_info_157_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_157_vecWen=0x%0h while the rhs_.io_diffCommits_info_157_vecWen=0x%0h",this.io_diffCommits_info_157_vecWen,rhs_.io_diffCommits_info_157_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_157_v0Wen!=rhs_.io_diffCommits_info_157_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_157_v0Wen=0x%0h while the rhs_.io_diffCommits_info_157_v0Wen=0x%0h",this.io_diffCommits_info_157_v0Wen,rhs_.io_diffCommits_info_157_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_157_vlWen!=rhs_.io_diffCommits_info_157_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_157_vlWen=0x%0h while the rhs_.io_diffCommits_info_157_vlWen=0x%0h",this.io_diffCommits_info_157_vlWen,rhs_.io_diffCommits_info_157_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_158_ldest!=rhs_.io_diffCommits_info_158_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_158_ldest=0x%0h while the rhs_.io_diffCommits_info_158_ldest=0x%0h",this.io_diffCommits_info_158_ldest,rhs_.io_diffCommits_info_158_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_158_pdest!=rhs_.io_diffCommits_info_158_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_158_pdest=0x%0h while the rhs_.io_diffCommits_info_158_pdest=0x%0h",this.io_diffCommits_info_158_pdest,rhs_.io_diffCommits_info_158_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_158_rfWen!=rhs_.io_diffCommits_info_158_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_158_rfWen=0x%0h while the rhs_.io_diffCommits_info_158_rfWen=0x%0h",this.io_diffCommits_info_158_rfWen,rhs_.io_diffCommits_info_158_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_158_fpWen!=rhs_.io_diffCommits_info_158_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_158_fpWen=0x%0h while the rhs_.io_diffCommits_info_158_fpWen=0x%0h",this.io_diffCommits_info_158_fpWen,rhs_.io_diffCommits_info_158_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_158_vecWen!=rhs_.io_diffCommits_info_158_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_158_vecWen=0x%0h while the rhs_.io_diffCommits_info_158_vecWen=0x%0h",this.io_diffCommits_info_158_vecWen,rhs_.io_diffCommits_info_158_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_158_v0Wen!=rhs_.io_diffCommits_info_158_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_158_v0Wen=0x%0h while the rhs_.io_diffCommits_info_158_v0Wen=0x%0h",this.io_diffCommits_info_158_v0Wen,rhs_.io_diffCommits_info_158_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_158_vlWen!=rhs_.io_diffCommits_info_158_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_158_vlWen=0x%0h while the rhs_.io_diffCommits_info_158_vlWen=0x%0h",this.io_diffCommits_info_158_vlWen,rhs_.io_diffCommits_info_158_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_159_ldest!=rhs_.io_diffCommits_info_159_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_159_ldest=0x%0h while the rhs_.io_diffCommits_info_159_ldest=0x%0h",this.io_diffCommits_info_159_ldest,rhs_.io_diffCommits_info_159_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_159_pdest!=rhs_.io_diffCommits_info_159_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_159_pdest=0x%0h while the rhs_.io_diffCommits_info_159_pdest=0x%0h",this.io_diffCommits_info_159_pdest,rhs_.io_diffCommits_info_159_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_159_rfWen!=rhs_.io_diffCommits_info_159_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_159_rfWen=0x%0h while the rhs_.io_diffCommits_info_159_rfWen=0x%0h",this.io_diffCommits_info_159_rfWen,rhs_.io_diffCommits_info_159_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_159_fpWen!=rhs_.io_diffCommits_info_159_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_159_fpWen=0x%0h while the rhs_.io_diffCommits_info_159_fpWen=0x%0h",this.io_diffCommits_info_159_fpWen,rhs_.io_diffCommits_info_159_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_159_vecWen!=rhs_.io_diffCommits_info_159_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_159_vecWen=0x%0h while the rhs_.io_diffCommits_info_159_vecWen=0x%0h",this.io_diffCommits_info_159_vecWen,rhs_.io_diffCommits_info_159_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_159_v0Wen!=rhs_.io_diffCommits_info_159_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_159_v0Wen=0x%0h while the rhs_.io_diffCommits_info_159_v0Wen=0x%0h",this.io_diffCommits_info_159_v0Wen,rhs_.io_diffCommits_info_159_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_159_vlWen!=rhs_.io_diffCommits_info_159_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_159_vlWen=0x%0h while the rhs_.io_diffCommits_info_159_vlWen=0x%0h",this.io_diffCommits_info_159_vlWen,rhs_.io_diffCommits_info_159_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_160_ldest!=rhs_.io_diffCommits_info_160_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_160_ldest=0x%0h while the rhs_.io_diffCommits_info_160_ldest=0x%0h",this.io_diffCommits_info_160_ldest,rhs_.io_diffCommits_info_160_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_160_pdest!=rhs_.io_diffCommits_info_160_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_160_pdest=0x%0h while the rhs_.io_diffCommits_info_160_pdest=0x%0h",this.io_diffCommits_info_160_pdest,rhs_.io_diffCommits_info_160_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_160_rfWen!=rhs_.io_diffCommits_info_160_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_160_rfWen=0x%0h while the rhs_.io_diffCommits_info_160_rfWen=0x%0h",this.io_diffCommits_info_160_rfWen,rhs_.io_diffCommits_info_160_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_160_fpWen!=rhs_.io_diffCommits_info_160_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_160_fpWen=0x%0h while the rhs_.io_diffCommits_info_160_fpWen=0x%0h",this.io_diffCommits_info_160_fpWen,rhs_.io_diffCommits_info_160_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_160_vecWen!=rhs_.io_diffCommits_info_160_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_160_vecWen=0x%0h while the rhs_.io_diffCommits_info_160_vecWen=0x%0h",this.io_diffCommits_info_160_vecWen,rhs_.io_diffCommits_info_160_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_160_v0Wen!=rhs_.io_diffCommits_info_160_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_160_v0Wen=0x%0h while the rhs_.io_diffCommits_info_160_v0Wen=0x%0h",this.io_diffCommits_info_160_v0Wen,rhs_.io_diffCommits_info_160_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_160_vlWen!=rhs_.io_diffCommits_info_160_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_160_vlWen=0x%0h while the rhs_.io_diffCommits_info_160_vlWen=0x%0h",this.io_diffCommits_info_160_vlWen,rhs_.io_diffCommits_info_160_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_161_ldest!=rhs_.io_diffCommits_info_161_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_161_ldest=0x%0h while the rhs_.io_diffCommits_info_161_ldest=0x%0h",this.io_diffCommits_info_161_ldest,rhs_.io_diffCommits_info_161_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_161_pdest!=rhs_.io_diffCommits_info_161_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_161_pdest=0x%0h while the rhs_.io_diffCommits_info_161_pdest=0x%0h",this.io_diffCommits_info_161_pdest,rhs_.io_diffCommits_info_161_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_161_rfWen!=rhs_.io_diffCommits_info_161_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_161_rfWen=0x%0h while the rhs_.io_diffCommits_info_161_rfWen=0x%0h",this.io_diffCommits_info_161_rfWen,rhs_.io_diffCommits_info_161_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_161_fpWen!=rhs_.io_diffCommits_info_161_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_161_fpWen=0x%0h while the rhs_.io_diffCommits_info_161_fpWen=0x%0h",this.io_diffCommits_info_161_fpWen,rhs_.io_diffCommits_info_161_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_161_vecWen!=rhs_.io_diffCommits_info_161_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_161_vecWen=0x%0h while the rhs_.io_diffCommits_info_161_vecWen=0x%0h",this.io_diffCommits_info_161_vecWen,rhs_.io_diffCommits_info_161_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_161_v0Wen!=rhs_.io_diffCommits_info_161_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_161_v0Wen=0x%0h while the rhs_.io_diffCommits_info_161_v0Wen=0x%0h",this.io_diffCommits_info_161_v0Wen,rhs_.io_diffCommits_info_161_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_161_vlWen!=rhs_.io_diffCommits_info_161_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_161_vlWen=0x%0h while the rhs_.io_diffCommits_info_161_vlWen=0x%0h",this.io_diffCommits_info_161_vlWen,rhs_.io_diffCommits_info_161_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_162_ldest!=rhs_.io_diffCommits_info_162_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_162_ldest=0x%0h while the rhs_.io_diffCommits_info_162_ldest=0x%0h",this.io_diffCommits_info_162_ldest,rhs_.io_diffCommits_info_162_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_162_pdest!=rhs_.io_diffCommits_info_162_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_162_pdest=0x%0h while the rhs_.io_diffCommits_info_162_pdest=0x%0h",this.io_diffCommits_info_162_pdest,rhs_.io_diffCommits_info_162_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_162_rfWen!=rhs_.io_diffCommits_info_162_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_162_rfWen=0x%0h while the rhs_.io_diffCommits_info_162_rfWen=0x%0h",this.io_diffCommits_info_162_rfWen,rhs_.io_diffCommits_info_162_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_162_fpWen!=rhs_.io_diffCommits_info_162_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_162_fpWen=0x%0h while the rhs_.io_diffCommits_info_162_fpWen=0x%0h",this.io_diffCommits_info_162_fpWen,rhs_.io_diffCommits_info_162_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_162_vecWen!=rhs_.io_diffCommits_info_162_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_162_vecWen=0x%0h while the rhs_.io_diffCommits_info_162_vecWen=0x%0h",this.io_diffCommits_info_162_vecWen,rhs_.io_diffCommits_info_162_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_162_v0Wen!=rhs_.io_diffCommits_info_162_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_162_v0Wen=0x%0h while the rhs_.io_diffCommits_info_162_v0Wen=0x%0h",this.io_diffCommits_info_162_v0Wen,rhs_.io_diffCommits_info_162_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_162_vlWen!=rhs_.io_diffCommits_info_162_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_162_vlWen=0x%0h while the rhs_.io_diffCommits_info_162_vlWen=0x%0h",this.io_diffCommits_info_162_vlWen,rhs_.io_diffCommits_info_162_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_163_ldest!=rhs_.io_diffCommits_info_163_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_163_ldest=0x%0h while the rhs_.io_diffCommits_info_163_ldest=0x%0h",this.io_diffCommits_info_163_ldest,rhs_.io_diffCommits_info_163_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_163_pdest!=rhs_.io_diffCommits_info_163_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_163_pdest=0x%0h while the rhs_.io_diffCommits_info_163_pdest=0x%0h",this.io_diffCommits_info_163_pdest,rhs_.io_diffCommits_info_163_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_163_rfWen!=rhs_.io_diffCommits_info_163_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_163_rfWen=0x%0h while the rhs_.io_diffCommits_info_163_rfWen=0x%0h",this.io_diffCommits_info_163_rfWen,rhs_.io_diffCommits_info_163_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_163_fpWen!=rhs_.io_diffCommits_info_163_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_163_fpWen=0x%0h while the rhs_.io_diffCommits_info_163_fpWen=0x%0h",this.io_diffCommits_info_163_fpWen,rhs_.io_diffCommits_info_163_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_163_vecWen!=rhs_.io_diffCommits_info_163_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_163_vecWen=0x%0h while the rhs_.io_diffCommits_info_163_vecWen=0x%0h",this.io_diffCommits_info_163_vecWen,rhs_.io_diffCommits_info_163_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_163_v0Wen!=rhs_.io_diffCommits_info_163_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_163_v0Wen=0x%0h while the rhs_.io_diffCommits_info_163_v0Wen=0x%0h",this.io_diffCommits_info_163_v0Wen,rhs_.io_diffCommits_info_163_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_163_vlWen!=rhs_.io_diffCommits_info_163_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_163_vlWen=0x%0h while the rhs_.io_diffCommits_info_163_vlWen=0x%0h",this.io_diffCommits_info_163_vlWen,rhs_.io_diffCommits_info_163_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_164_ldest!=rhs_.io_diffCommits_info_164_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_164_ldest=0x%0h while the rhs_.io_diffCommits_info_164_ldest=0x%0h",this.io_diffCommits_info_164_ldest,rhs_.io_diffCommits_info_164_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_164_pdest!=rhs_.io_diffCommits_info_164_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_164_pdest=0x%0h while the rhs_.io_diffCommits_info_164_pdest=0x%0h",this.io_diffCommits_info_164_pdest,rhs_.io_diffCommits_info_164_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_164_rfWen!=rhs_.io_diffCommits_info_164_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_164_rfWen=0x%0h while the rhs_.io_diffCommits_info_164_rfWen=0x%0h",this.io_diffCommits_info_164_rfWen,rhs_.io_diffCommits_info_164_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_164_fpWen!=rhs_.io_diffCommits_info_164_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_164_fpWen=0x%0h while the rhs_.io_diffCommits_info_164_fpWen=0x%0h",this.io_diffCommits_info_164_fpWen,rhs_.io_diffCommits_info_164_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_164_vecWen!=rhs_.io_diffCommits_info_164_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_164_vecWen=0x%0h while the rhs_.io_diffCommits_info_164_vecWen=0x%0h",this.io_diffCommits_info_164_vecWen,rhs_.io_diffCommits_info_164_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_164_v0Wen!=rhs_.io_diffCommits_info_164_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_164_v0Wen=0x%0h while the rhs_.io_diffCommits_info_164_v0Wen=0x%0h",this.io_diffCommits_info_164_v0Wen,rhs_.io_diffCommits_info_164_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_164_vlWen!=rhs_.io_diffCommits_info_164_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_164_vlWen=0x%0h while the rhs_.io_diffCommits_info_164_vlWen=0x%0h",this.io_diffCommits_info_164_vlWen,rhs_.io_diffCommits_info_164_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_165_ldest!=rhs_.io_diffCommits_info_165_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_165_ldest=0x%0h while the rhs_.io_diffCommits_info_165_ldest=0x%0h",this.io_diffCommits_info_165_ldest,rhs_.io_diffCommits_info_165_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_165_pdest!=rhs_.io_diffCommits_info_165_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_165_pdest=0x%0h while the rhs_.io_diffCommits_info_165_pdest=0x%0h",this.io_diffCommits_info_165_pdest,rhs_.io_diffCommits_info_165_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_165_rfWen!=rhs_.io_diffCommits_info_165_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_165_rfWen=0x%0h while the rhs_.io_diffCommits_info_165_rfWen=0x%0h",this.io_diffCommits_info_165_rfWen,rhs_.io_diffCommits_info_165_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_165_fpWen!=rhs_.io_diffCommits_info_165_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_165_fpWen=0x%0h while the rhs_.io_diffCommits_info_165_fpWen=0x%0h",this.io_diffCommits_info_165_fpWen,rhs_.io_diffCommits_info_165_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_165_vecWen!=rhs_.io_diffCommits_info_165_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_165_vecWen=0x%0h while the rhs_.io_diffCommits_info_165_vecWen=0x%0h",this.io_diffCommits_info_165_vecWen,rhs_.io_diffCommits_info_165_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_165_v0Wen!=rhs_.io_diffCommits_info_165_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_165_v0Wen=0x%0h while the rhs_.io_diffCommits_info_165_v0Wen=0x%0h",this.io_diffCommits_info_165_v0Wen,rhs_.io_diffCommits_info_165_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_165_vlWen!=rhs_.io_diffCommits_info_165_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_165_vlWen=0x%0h while the rhs_.io_diffCommits_info_165_vlWen=0x%0h",this.io_diffCommits_info_165_vlWen,rhs_.io_diffCommits_info_165_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_166_ldest!=rhs_.io_diffCommits_info_166_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_166_ldest=0x%0h while the rhs_.io_diffCommits_info_166_ldest=0x%0h",this.io_diffCommits_info_166_ldest,rhs_.io_diffCommits_info_166_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_166_pdest!=rhs_.io_diffCommits_info_166_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_166_pdest=0x%0h while the rhs_.io_diffCommits_info_166_pdest=0x%0h",this.io_diffCommits_info_166_pdest,rhs_.io_diffCommits_info_166_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_166_rfWen!=rhs_.io_diffCommits_info_166_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_166_rfWen=0x%0h while the rhs_.io_diffCommits_info_166_rfWen=0x%0h",this.io_diffCommits_info_166_rfWen,rhs_.io_diffCommits_info_166_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_166_fpWen!=rhs_.io_diffCommits_info_166_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_166_fpWen=0x%0h while the rhs_.io_diffCommits_info_166_fpWen=0x%0h",this.io_diffCommits_info_166_fpWen,rhs_.io_diffCommits_info_166_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_166_vecWen!=rhs_.io_diffCommits_info_166_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_166_vecWen=0x%0h while the rhs_.io_diffCommits_info_166_vecWen=0x%0h",this.io_diffCommits_info_166_vecWen,rhs_.io_diffCommits_info_166_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_166_v0Wen!=rhs_.io_diffCommits_info_166_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_166_v0Wen=0x%0h while the rhs_.io_diffCommits_info_166_v0Wen=0x%0h",this.io_diffCommits_info_166_v0Wen,rhs_.io_diffCommits_info_166_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_166_vlWen!=rhs_.io_diffCommits_info_166_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_166_vlWen=0x%0h while the rhs_.io_diffCommits_info_166_vlWen=0x%0h",this.io_diffCommits_info_166_vlWen,rhs_.io_diffCommits_info_166_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_167_ldest!=rhs_.io_diffCommits_info_167_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_167_ldest=0x%0h while the rhs_.io_diffCommits_info_167_ldest=0x%0h",this.io_diffCommits_info_167_ldest,rhs_.io_diffCommits_info_167_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_167_pdest!=rhs_.io_diffCommits_info_167_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_167_pdest=0x%0h while the rhs_.io_diffCommits_info_167_pdest=0x%0h",this.io_diffCommits_info_167_pdest,rhs_.io_diffCommits_info_167_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_167_rfWen!=rhs_.io_diffCommits_info_167_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_167_rfWen=0x%0h while the rhs_.io_diffCommits_info_167_rfWen=0x%0h",this.io_diffCommits_info_167_rfWen,rhs_.io_diffCommits_info_167_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_167_fpWen!=rhs_.io_diffCommits_info_167_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_167_fpWen=0x%0h while the rhs_.io_diffCommits_info_167_fpWen=0x%0h",this.io_diffCommits_info_167_fpWen,rhs_.io_diffCommits_info_167_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_167_vecWen!=rhs_.io_diffCommits_info_167_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_167_vecWen=0x%0h while the rhs_.io_diffCommits_info_167_vecWen=0x%0h",this.io_diffCommits_info_167_vecWen,rhs_.io_diffCommits_info_167_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_167_v0Wen!=rhs_.io_diffCommits_info_167_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_167_v0Wen=0x%0h while the rhs_.io_diffCommits_info_167_v0Wen=0x%0h",this.io_diffCommits_info_167_v0Wen,rhs_.io_diffCommits_info_167_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_167_vlWen!=rhs_.io_diffCommits_info_167_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_167_vlWen=0x%0h while the rhs_.io_diffCommits_info_167_vlWen=0x%0h",this.io_diffCommits_info_167_vlWen,rhs_.io_diffCommits_info_167_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_168_ldest!=rhs_.io_diffCommits_info_168_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_168_ldest=0x%0h while the rhs_.io_diffCommits_info_168_ldest=0x%0h",this.io_diffCommits_info_168_ldest,rhs_.io_diffCommits_info_168_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_168_pdest!=rhs_.io_diffCommits_info_168_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_168_pdest=0x%0h while the rhs_.io_diffCommits_info_168_pdest=0x%0h",this.io_diffCommits_info_168_pdest,rhs_.io_diffCommits_info_168_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_168_rfWen!=rhs_.io_diffCommits_info_168_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_168_rfWen=0x%0h while the rhs_.io_diffCommits_info_168_rfWen=0x%0h",this.io_diffCommits_info_168_rfWen,rhs_.io_diffCommits_info_168_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_168_fpWen!=rhs_.io_diffCommits_info_168_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_168_fpWen=0x%0h while the rhs_.io_diffCommits_info_168_fpWen=0x%0h",this.io_diffCommits_info_168_fpWen,rhs_.io_diffCommits_info_168_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_168_vecWen!=rhs_.io_diffCommits_info_168_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_168_vecWen=0x%0h while the rhs_.io_diffCommits_info_168_vecWen=0x%0h",this.io_diffCommits_info_168_vecWen,rhs_.io_diffCommits_info_168_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_168_v0Wen!=rhs_.io_diffCommits_info_168_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_168_v0Wen=0x%0h while the rhs_.io_diffCommits_info_168_v0Wen=0x%0h",this.io_diffCommits_info_168_v0Wen,rhs_.io_diffCommits_info_168_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_168_vlWen!=rhs_.io_diffCommits_info_168_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_168_vlWen=0x%0h while the rhs_.io_diffCommits_info_168_vlWen=0x%0h",this.io_diffCommits_info_168_vlWen,rhs_.io_diffCommits_info_168_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_169_ldest!=rhs_.io_diffCommits_info_169_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_169_ldest=0x%0h while the rhs_.io_diffCommits_info_169_ldest=0x%0h",this.io_diffCommits_info_169_ldest,rhs_.io_diffCommits_info_169_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_169_pdest!=rhs_.io_diffCommits_info_169_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_169_pdest=0x%0h while the rhs_.io_diffCommits_info_169_pdest=0x%0h",this.io_diffCommits_info_169_pdest,rhs_.io_diffCommits_info_169_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_169_rfWen!=rhs_.io_diffCommits_info_169_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_169_rfWen=0x%0h while the rhs_.io_diffCommits_info_169_rfWen=0x%0h",this.io_diffCommits_info_169_rfWen,rhs_.io_diffCommits_info_169_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_169_fpWen!=rhs_.io_diffCommits_info_169_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_169_fpWen=0x%0h while the rhs_.io_diffCommits_info_169_fpWen=0x%0h",this.io_diffCommits_info_169_fpWen,rhs_.io_diffCommits_info_169_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_169_vecWen!=rhs_.io_diffCommits_info_169_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_169_vecWen=0x%0h while the rhs_.io_diffCommits_info_169_vecWen=0x%0h",this.io_diffCommits_info_169_vecWen,rhs_.io_diffCommits_info_169_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_169_v0Wen!=rhs_.io_diffCommits_info_169_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_169_v0Wen=0x%0h while the rhs_.io_diffCommits_info_169_v0Wen=0x%0h",this.io_diffCommits_info_169_v0Wen,rhs_.io_diffCommits_info_169_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_169_vlWen!=rhs_.io_diffCommits_info_169_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_169_vlWen=0x%0h while the rhs_.io_diffCommits_info_169_vlWen=0x%0h",this.io_diffCommits_info_169_vlWen,rhs_.io_diffCommits_info_169_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_170_ldest!=rhs_.io_diffCommits_info_170_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_170_ldest=0x%0h while the rhs_.io_diffCommits_info_170_ldest=0x%0h",this.io_diffCommits_info_170_ldest,rhs_.io_diffCommits_info_170_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_170_pdest!=rhs_.io_diffCommits_info_170_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_170_pdest=0x%0h while the rhs_.io_diffCommits_info_170_pdest=0x%0h",this.io_diffCommits_info_170_pdest,rhs_.io_diffCommits_info_170_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_170_rfWen!=rhs_.io_diffCommits_info_170_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_170_rfWen=0x%0h while the rhs_.io_diffCommits_info_170_rfWen=0x%0h",this.io_diffCommits_info_170_rfWen,rhs_.io_diffCommits_info_170_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_170_fpWen!=rhs_.io_diffCommits_info_170_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_170_fpWen=0x%0h while the rhs_.io_diffCommits_info_170_fpWen=0x%0h",this.io_diffCommits_info_170_fpWen,rhs_.io_diffCommits_info_170_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_170_vecWen!=rhs_.io_diffCommits_info_170_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_170_vecWen=0x%0h while the rhs_.io_diffCommits_info_170_vecWen=0x%0h",this.io_diffCommits_info_170_vecWen,rhs_.io_diffCommits_info_170_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_170_v0Wen!=rhs_.io_diffCommits_info_170_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_170_v0Wen=0x%0h while the rhs_.io_diffCommits_info_170_v0Wen=0x%0h",this.io_diffCommits_info_170_v0Wen,rhs_.io_diffCommits_info_170_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_170_vlWen!=rhs_.io_diffCommits_info_170_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_170_vlWen=0x%0h while the rhs_.io_diffCommits_info_170_vlWen=0x%0h",this.io_diffCommits_info_170_vlWen,rhs_.io_diffCommits_info_170_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_171_ldest!=rhs_.io_diffCommits_info_171_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_171_ldest=0x%0h while the rhs_.io_diffCommits_info_171_ldest=0x%0h",this.io_diffCommits_info_171_ldest,rhs_.io_diffCommits_info_171_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_171_pdest!=rhs_.io_diffCommits_info_171_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_171_pdest=0x%0h while the rhs_.io_diffCommits_info_171_pdest=0x%0h",this.io_diffCommits_info_171_pdest,rhs_.io_diffCommits_info_171_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_171_rfWen!=rhs_.io_diffCommits_info_171_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_171_rfWen=0x%0h while the rhs_.io_diffCommits_info_171_rfWen=0x%0h",this.io_diffCommits_info_171_rfWen,rhs_.io_diffCommits_info_171_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_171_fpWen!=rhs_.io_diffCommits_info_171_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_171_fpWen=0x%0h while the rhs_.io_diffCommits_info_171_fpWen=0x%0h",this.io_diffCommits_info_171_fpWen,rhs_.io_diffCommits_info_171_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_171_vecWen!=rhs_.io_diffCommits_info_171_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_171_vecWen=0x%0h while the rhs_.io_diffCommits_info_171_vecWen=0x%0h",this.io_diffCommits_info_171_vecWen,rhs_.io_diffCommits_info_171_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_171_v0Wen!=rhs_.io_diffCommits_info_171_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_171_v0Wen=0x%0h while the rhs_.io_diffCommits_info_171_v0Wen=0x%0h",this.io_diffCommits_info_171_v0Wen,rhs_.io_diffCommits_info_171_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_171_vlWen!=rhs_.io_diffCommits_info_171_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_171_vlWen=0x%0h while the rhs_.io_diffCommits_info_171_vlWen=0x%0h",this.io_diffCommits_info_171_vlWen,rhs_.io_diffCommits_info_171_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_172_ldest!=rhs_.io_diffCommits_info_172_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_172_ldest=0x%0h while the rhs_.io_diffCommits_info_172_ldest=0x%0h",this.io_diffCommits_info_172_ldest,rhs_.io_diffCommits_info_172_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_172_pdest!=rhs_.io_diffCommits_info_172_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_172_pdest=0x%0h while the rhs_.io_diffCommits_info_172_pdest=0x%0h",this.io_diffCommits_info_172_pdest,rhs_.io_diffCommits_info_172_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_172_rfWen!=rhs_.io_diffCommits_info_172_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_172_rfWen=0x%0h while the rhs_.io_diffCommits_info_172_rfWen=0x%0h",this.io_diffCommits_info_172_rfWen,rhs_.io_diffCommits_info_172_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_172_fpWen!=rhs_.io_diffCommits_info_172_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_172_fpWen=0x%0h while the rhs_.io_diffCommits_info_172_fpWen=0x%0h",this.io_diffCommits_info_172_fpWen,rhs_.io_diffCommits_info_172_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_172_vecWen!=rhs_.io_diffCommits_info_172_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_172_vecWen=0x%0h while the rhs_.io_diffCommits_info_172_vecWen=0x%0h",this.io_diffCommits_info_172_vecWen,rhs_.io_diffCommits_info_172_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_172_v0Wen!=rhs_.io_diffCommits_info_172_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_172_v0Wen=0x%0h while the rhs_.io_diffCommits_info_172_v0Wen=0x%0h",this.io_diffCommits_info_172_v0Wen,rhs_.io_diffCommits_info_172_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_172_vlWen!=rhs_.io_diffCommits_info_172_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_172_vlWen=0x%0h while the rhs_.io_diffCommits_info_172_vlWen=0x%0h",this.io_diffCommits_info_172_vlWen,rhs_.io_diffCommits_info_172_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_173_ldest!=rhs_.io_diffCommits_info_173_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_173_ldest=0x%0h while the rhs_.io_diffCommits_info_173_ldest=0x%0h",this.io_diffCommits_info_173_ldest,rhs_.io_diffCommits_info_173_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_173_pdest!=rhs_.io_diffCommits_info_173_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_173_pdest=0x%0h while the rhs_.io_diffCommits_info_173_pdest=0x%0h",this.io_diffCommits_info_173_pdest,rhs_.io_diffCommits_info_173_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_173_rfWen!=rhs_.io_diffCommits_info_173_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_173_rfWen=0x%0h while the rhs_.io_diffCommits_info_173_rfWen=0x%0h",this.io_diffCommits_info_173_rfWen,rhs_.io_diffCommits_info_173_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_173_fpWen!=rhs_.io_diffCommits_info_173_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_173_fpWen=0x%0h while the rhs_.io_diffCommits_info_173_fpWen=0x%0h",this.io_diffCommits_info_173_fpWen,rhs_.io_diffCommits_info_173_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_173_vecWen!=rhs_.io_diffCommits_info_173_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_173_vecWen=0x%0h while the rhs_.io_diffCommits_info_173_vecWen=0x%0h",this.io_diffCommits_info_173_vecWen,rhs_.io_diffCommits_info_173_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_173_v0Wen!=rhs_.io_diffCommits_info_173_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_173_v0Wen=0x%0h while the rhs_.io_diffCommits_info_173_v0Wen=0x%0h",this.io_diffCommits_info_173_v0Wen,rhs_.io_diffCommits_info_173_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_173_vlWen!=rhs_.io_diffCommits_info_173_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_173_vlWen=0x%0h while the rhs_.io_diffCommits_info_173_vlWen=0x%0h",this.io_diffCommits_info_173_vlWen,rhs_.io_diffCommits_info_173_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_174_ldest!=rhs_.io_diffCommits_info_174_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_174_ldest=0x%0h while the rhs_.io_diffCommits_info_174_ldest=0x%0h",this.io_diffCommits_info_174_ldest,rhs_.io_diffCommits_info_174_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_174_pdest!=rhs_.io_diffCommits_info_174_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_174_pdest=0x%0h while the rhs_.io_diffCommits_info_174_pdest=0x%0h",this.io_diffCommits_info_174_pdest,rhs_.io_diffCommits_info_174_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_174_rfWen!=rhs_.io_diffCommits_info_174_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_174_rfWen=0x%0h while the rhs_.io_diffCommits_info_174_rfWen=0x%0h",this.io_diffCommits_info_174_rfWen,rhs_.io_diffCommits_info_174_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_174_fpWen!=rhs_.io_diffCommits_info_174_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_174_fpWen=0x%0h while the rhs_.io_diffCommits_info_174_fpWen=0x%0h",this.io_diffCommits_info_174_fpWen,rhs_.io_diffCommits_info_174_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_174_vecWen!=rhs_.io_diffCommits_info_174_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_174_vecWen=0x%0h while the rhs_.io_diffCommits_info_174_vecWen=0x%0h",this.io_diffCommits_info_174_vecWen,rhs_.io_diffCommits_info_174_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_174_v0Wen!=rhs_.io_diffCommits_info_174_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_174_v0Wen=0x%0h while the rhs_.io_diffCommits_info_174_v0Wen=0x%0h",this.io_diffCommits_info_174_v0Wen,rhs_.io_diffCommits_info_174_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_174_vlWen!=rhs_.io_diffCommits_info_174_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_174_vlWen=0x%0h while the rhs_.io_diffCommits_info_174_vlWen=0x%0h",this.io_diffCommits_info_174_vlWen,rhs_.io_diffCommits_info_174_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_175_ldest!=rhs_.io_diffCommits_info_175_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_175_ldest=0x%0h while the rhs_.io_diffCommits_info_175_ldest=0x%0h",this.io_diffCommits_info_175_ldest,rhs_.io_diffCommits_info_175_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_175_pdest!=rhs_.io_diffCommits_info_175_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_175_pdest=0x%0h while the rhs_.io_diffCommits_info_175_pdest=0x%0h",this.io_diffCommits_info_175_pdest,rhs_.io_diffCommits_info_175_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_175_rfWen!=rhs_.io_diffCommits_info_175_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_175_rfWen=0x%0h while the rhs_.io_diffCommits_info_175_rfWen=0x%0h",this.io_diffCommits_info_175_rfWen,rhs_.io_diffCommits_info_175_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_175_fpWen!=rhs_.io_diffCommits_info_175_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_175_fpWen=0x%0h while the rhs_.io_diffCommits_info_175_fpWen=0x%0h",this.io_diffCommits_info_175_fpWen,rhs_.io_diffCommits_info_175_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_175_vecWen!=rhs_.io_diffCommits_info_175_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_175_vecWen=0x%0h while the rhs_.io_diffCommits_info_175_vecWen=0x%0h",this.io_diffCommits_info_175_vecWen,rhs_.io_diffCommits_info_175_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_175_v0Wen!=rhs_.io_diffCommits_info_175_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_175_v0Wen=0x%0h while the rhs_.io_diffCommits_info_175_v0Wen=0x%0h",this.io_diffCommits_info_175_v0Wen,rhs_.io_diffCommits_info_175_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_175_vlWen!=rhs_.io_diffCommits_info_175_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_175_vlWen=0x%0h while the rhs_.io_diffCommits_info_175_vlWen=0x%0h",this.io_diffCommits_info_175_vlWen,rhs_.io_diffCommits_info_175_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_176_ldest!=rhs_.io_diffCommits_info_176_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_176_ldest=0x%0h while the rhs_.io_diffCommits_info_176_ldest=0x%0h",this.io_diffCommits_info_176_ldest,rhs_.io_diffCommits_info_176_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_176_pdest!=rhs_.io_diffCommits_info_176_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_176_pdest=0x%0h while the rhs_.io_diffCommits_info_176_pdest=0x%0h",this.io_diffCommits_info_176_pdest,rhs_.io_diffCommits_info_176_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_176_rfWen!=rhs_.io_diffCommits_info_176_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_176_rfWen=0x%0h while the rhs_.io_diffCommits_info_176_rfWen=0x%0h",this.io_diffCommits_info_176_rfWen,rhs_.io_diffCommits_info_176_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_176_fpWen!=rhs_.io_diffCommits_info_176_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_176_fpWen=0x%0h while the rhs_.io_diffCommits_info_176_fpWen=0x%0h",this.io_diffCommits_info_176_fpWen,rhs_.io_diffCommits_info_176_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_176_vecWen!=rhs_.io_diffCommits_info_176_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_176_vecWen=0x%0h while the rhs_.io_diffCommits_info_176_vecWen=0x%0h",this.io_diffCommits_info_176_vecWen,rhs_.io_diffCommits_info_176_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_176_v0Wen!=rhs_.io_diffCommits_info_176_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_176_v0Wen=0x%0h while the rhs_.io_diffCommits_info_176_v0Wen=0x%0h",this.io_diffCommits_info_176_v0Wen,rhs_.io_diffCommits_info_176_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_176_vlWen!=rhs_.io_diffCommits_info_176_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_176_vlWen=0x%0h while the rhs_.io_diffCommits_info_176_vlWen=0x%0h",this.io_diffCommits_info_176_vlWen,rhs_.io_diffCommits_info_176_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_177_ldest!=rhs_.io_diffCommits_info_177_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_177_ldest=0x%0h while the rhs_.io_diffCommits_info_177_ldest=0x%0h",this.io_diffCommits_info_177_ldest,rhs_.io_diffCommits_info_177_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_177_pdest!=rhs_.io_diffCommits_info_177_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_177_pdest=0x%0h while the rhs_.io_diffCommits_info_177_pdest=0x%0h",this.io_diffCommits_info_177_pdest,rhs_.io_diffCommits_info_177_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_177_rfWen!=rhs_.io_diffCommits_info_177_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_177_rfWen=0x%0h while the rhs_.io_diffCommits_info_177_rfWen=0x%0h",this.io_diffCommits_info_177_rfWen,rhs_.io_diffCommits_info_177_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_177_fpWen!=rhs_.io_diffCommits_info_177_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_177_fpWen=0x%0h while the rhs_.io_diffCommits_info_177_fpWen=0x%0h",this.io_diffCommits_info_177_fpWen,rhs_.io_diffCommits_info_177_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_177_vecWen!=rhs_.io_diffCommits_info_177_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_177_vecWen=0x%0h while the rhs_.io_diffCommits_info_177_vecWen=0x%0h",this.io_diffCommits_info_177_vecWen,rhs_.io_diffCommits_info_177_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_177_v0Wen!=rhs_.io_diffCommits_info_177_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_177_v0Wen=0x%0h while the rhs_.io_diffCommits_info_177_v0Wen=0x%0h",this.io_diffCommits_info_177_v0Wen,rhs_.io_diffCommits_info_177_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_177_vlWen!=rhs_.io_diffCommits_info_177_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_177_vlWen=0x%0h while the rhs_.io_diffCommits_info_177_vlWen=0x%0h",this.io_diffCommits_info_177_vlWen,rhs_.io_diffCommits_info_177_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_178_ldest!=rhs_.io_diffCommits_info_178_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_178_ldest=0x%0h while the rhs_.io_diffCommits_info_178_ldest=0x%0h",this.io_diffCommits_info_178_ldest,rhs_.io_diffCommits_info_178_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_178_pdest!=rhs_.io_diffCommits_info_178_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_178_pdest=0x%0h while the rhs_.io_diffCommits_info_178_pdest=0x%0h",this.io_diffCommits_info_178_pdest,rhs_.io_diffCommits_info_178_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_178_rfWen!=rhs_.io_diffCommits_info_178_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_178_rfWen=0x%0h while the rhs_.io_diffCommits_info_178_rfWen=0x%0h",this.io_diffCommits_info_178_rfWen,rhs_.io_diffCommits_info_178_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_178_fpWen!=rhs_.io_diffCommits_info_178_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_178_fpWen=0x%0h while the rhs_.io_diffCommits_info_178_fpWen=0x%0h",this.io_diffCommits_info_178_fpWen,rhs_.io_diffCommits_info_178_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_178_vecWen!=rhs_.io_diffCommits_info_178_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_178_vecWen=0x%0h while the rhs_.io_diffCommits_info_178_vecWen=0x%0h",this.io_diffCommits_info_178_vecWen,rhs_.io_diffCommits_info_178_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_178_v0Wen!=rhs_.io_diffCommits_info_178_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_178_v0Wen=0x%0h while the rhs_.io_diffCommits_info_178_v0Wen=0x%0h",this.io_diffCommits_info_178_v0Wen,rhs_.io_diffCommits_info_178_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_178_vlWen!=rhs_.io_diffCommits_info_178_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_178_vlWen=0x%0h while the rhs_.io_diffCommits_info_178_vlWen=0x%0h",this.io_diffCommits_info_178_vlWen,rhs_.io_diffCommits_info_178_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_179_ldest!=rhs_.io_diffCommits_info_179_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_179_ldest=0x%0h while the rhs_.io_diffCommits_info_179_ldest=0x%0h",this.io_diffCommits_info_179_ldest,rhs_.io_diffCommits_info_179_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_179_pdest!=rhs_.io_diffCommits_info_179_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_179_pdest=0x%0h while the rhs_.io_diffCommits_info_179_pdest=0x%0h",this.io_diffCommits_info_179_pdest,rhs_.io_diffCommits_info_179_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_179_rfWen!=rhs_.io_diffCommits_info_179_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_179_rfWen=0x%0h while the rhs_.io_diffCommits_info_179_rfWen=0x%0h",this.io_diffCommits_info_179_rfWen,rhs_.io_diffCommits_info_179_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_179_fpWen!=rhs_.io_diffCommits_info_179_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_179_fpWen=0x%0h while the rhs_.io_diffCommits_info_179_fpWen=0x%0h",this.io_diffCommits_info_179_fpWen,rhs_.io_diffCommits_info_179_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_179_vecWen!=rhs_.io_diffCommits_info_179_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_179_vecWen=0x%0h while the rhs_.io_diffCommits_info_179_vecWen=0x%0h",this.io_diffCommits_info_179_vecWen,rhs_.io_diffCommits_info_179_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_179_v0Wen!=rhs_.io_diffCommits_info_179_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_179_v0Wen=0x%0h while the rhs_.io_diffCommits_info_179_v0Wen=0x%0h",this.io_diffCommits_info_179_v0Wen,rhs_.io_diffCommits_info_179_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_179_vlWen!=rhs_.io_diffCommits_info_179_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_179_vlWen=0x%0h while the rhs_.io_diffCommits_info_179_vlWen=0x%0h",this.io_diffCommits_info_179_vlWen,rhs_.io_diffCommits_info_179_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_180_ldest!=rhs_.io_diffCommits_info_180_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_180_ldest=0x%0h while the rhs_.io_diffCommits_info_180_ldest=0x%0h",this.io_diffCommits_info_180_ldest,rhs_.io_diffCommits_info_180_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_180_pdest!=rhs_.io_diffCommits_info_180_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_180_pdest=0x%0h while the rhs_.io_diffCommits_info_180_pdest=0x%0h",this.io_diffCommits_info_180_pdest,rhs_.io_diffCommits_info_180_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_180_rfWen!=rhs_.io_diffCommits_info_180_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_180_rfWen=0x%0h while the rhs_.io_diffCommits_info_180_rfWen=0x%0h",this.io_diffCommits_info_180_rfWen,rhs_.io_diffCommits_info_180_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_180_fpWen!=rhs_.io_diffCommits_info_180_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_180_fpWen=0x%0h while the rhs_.io_diffCommits_info_180_fpWen=0x%0h",this.io_diffCommits_info_180_fpWen,rhs_.io_diffCommits_info_180_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_180_vecWen!=rhs_.io_diffCommits_info_180_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_180_vecWen=0x%0h while the rhs_.io_diffCommits_info_180_vecWen=0x%0h",this.io_diffCommits_info_180_vecWen,rhs_.io_diffCommits_info_180_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_180_v0Wen!=rhs_.io_diffCommits_info_180_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_180_v0Wen=0x%0h while the rhs_.io_diffCommits_info_180_v0Wen=0x%0h",this.io_diffCommits_info_180_v0Wen,rhs_.io_diffCommits_info_180_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_180_vlWen!=rhs_.io_diffCommits_info_180_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_180_vlWen=0x%0h while the rhs_.io_diffCommits_info_180_vlWen=0x%0h",this.io_diffCommits_info_180_vlWen,rhs_.io_diffCommits_info_180_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_181_ldest!=rhs_.io_diffCommits_info_181_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_181_ldest=0x%0h while the rhs_.io_diffCommits_info_181_ldest=0x%0h",this.io_diffCommits_info_181_ldest,rhs_.io_diffCommits_info_181_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_181_pdest!=rhs_.io_diffCommits_info_181_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_181_pdest=0x%0h while the rhs_.io_diffCommits_info_181_pdest=0x%0h",this.io_diffCommits_info_181_pdest,rhs_.io_diffCommits_info_181_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_181_rfWen!=rhs_.io_diffCommits_info_181_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_181_rfWen=0x%0h while the rhs_.io_diffCommits_info_181_rfWen=0x%0h",this.io_diffCommits_info_181_rfWen,rhs_.io_diffCommits_info_181_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_181_fpWen!=rhs_.io_diffCommits_info_181_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_181_fpWen=0x%0h while the rhs_.io_diffCommits_info_181_fpWen=0x%0h",this.io_diffCommits_info_181_fpWen,rhs_.io_diffCommits_info_181_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_181_vecWen!=rhs_.io_diffCommits_info_181_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_181_vecWen=0x%0h while the rhs_.io_diffCommits_info_181_vecWen=0x%0h",this.io_diffCommits_info_181_vecWen,rhs_.io_diffCommits_info_181_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_181_v0Wen!=rhs_.io_diffCommits_info_181_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_181_v0Wen=0x%0h while the rhs_.io_diffCommits_info_181_v0Wen=0x%0h",this.io_diffCommits_info_181_v0Wen,rhs_.io_diffCommits_info_181_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_181_vlWen!=rhs_.io_diffCommits_info_181_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_181_vlWen=0x%0h while the rhs_.io_diffCommits_info_181_vlWen=0x%0h",this.io_diffCommits_info_181_vlWen,rhs_.io_diffCommits_info_181_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_182_ldest!=rhs_.io_diffCommits_info_182_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_182_ldest=0x%0h while the rhs_.io_diffCommits_info_182_ldest=0x%0h",this.io_diffCommits_info_182_ldest,rhs_.io_diffCommits_info_182_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_182_pdest!=rhs_.io_diffCommits_info_182_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_182_pdest=0x%0h while the rhs_.io_diffCommits_info_182_pdest=0x%0h",this.io_diffCommits_info_182_pdest,rhs_.io_diffCommits_info_182_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_182_rfWen!=rhs_.io_diffCommits_info_182_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_182_rfWen=0x%0h while the rhs_.io_diffCommits_info_182_rfWen=0x%0h",this.io_diffCommits_info_182_rfWen,rhs_.io_diffCommits_info_182_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_182_fpWen!=rhs_.io_diffCommits_info_182_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_182_fpWen=0x%0h while the rhs_.io_diffCommits_info_182_fpWen=0x%0h",this.io_diffCommits_info_182_fpWen,rhs_.io_diffCommits_info_182_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_182_vecWen!=rhs_.io_diffCommits_info_182_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_182_vecWen=0x%0h while the rhs_.io_diffCommits_info_182_vecWen=0x%0h",this.io_diffCommits_info_182_vecWen,rhs_.io_diffCommits_info_182_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_182_v0Wen!=rhs_.io_diffCommits_info_182_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_182_v0Wen=0x%0h while the rhs_.io_diffCommits_info_182_v0Wen=0x%0h",this.io_diffCommits_info_182_v0Wen,rhs_.io_diffCommits_info_182_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_182_vlWen!=rhs_.io_diffCommits_info_182_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_182_vlWen=0x%0h while the rhs_.io_diffCommits_info_182_vlWen=0x%0h",this.io_diffCommits_info_182_vlWen,rhs_.io_diffCommits_info_182_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_183_ldest!=rhs_.io_diffCommits_info_183_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_183_ldest=0x%0h while the rhs_.io_diffCommits_info_183_ldest=0x%0h",this.io_diffCommits_info_183_ldest,rhs_.io_diffCommits_info_183_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_183_pdest!=rhs_.io_diffCommits_info_183_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_183_pdest=0x%0h while the rhs_.io_diffCommits_info_183_pdest=0x%0h",this.io_diffCommits_info_183_pdest,rhs_.io_diffCommits_info_183_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_183_rfWen!=rhs_.io_diffCommits_info_183_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_183_rfWen=0x%0h while the rhs_.io_diffCommits_info_183_rfWen=0x%0h",this.io_diffCommits_info_183_rfWen,rhs_.io_diffCommits_info_183_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_183_fpWen!=rhs_.io_diffCommits_info_183_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_183_fpWen=0x%0h while the rhs_.io_diffCommits_info_183_fpWen=0x%0h",this.io_diffCommits_info_183_fpWen,rhs_.io_diffCommits_info_183_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_183_vecWen!=rhs_.io_diffCommits_info_183_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_183_vecWen=0x%0h while the rhs_.io_diffCommits_info_183_vecWen=0x%0h",this.io_diffCommits_info_183_vecWen,rhs_.io_diffCommits_info_183_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_183_v0Wen!=rhs_.io_diffCommits_info_183_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_183_v0Wen=0x%0h while the rhs_.io_diffCommits_info_183_v0Wen=0x%0h",this.io_diffCommits_info_183_v0Wen,rhs_.io_diffCommits_info_183_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_183_vlWen!=rhs_.io_diffCommits_info_183_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_183_vlWen=0x%0h while the rhs_.io_diffCommits_info_183_vlWen=0x%0h",this.io_diffCommits_info_183_vlWen,rhs_.io_diffCommits_info_183_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_184_ldest!=rhs_.io_diffCommits_info_184_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_184_ldest=0x%0h while the rhs_.io_diffCommits_info_184_ldest=0x%0h",this.io_diffCommits_info_184_ldest,rhs_.io_diffCommits_info_184_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_184_pdest!=rhs_.io_diffCommits_info_184_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_184_pdest=0x%0h while the rhs_.io_diffCommits_info_184_pdest=0x%0h",this.io_diffCommits_info_184_pdest,rhs_.io_diffCommits_info_184_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_184_rfWen!=rhs_.io_diffCommits_info_184_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_184_rfWen=0x%0h while the rhs_.io_diffCommits_info_184_rfWen=0x%0h",this.io_diffCommits_info_184_rfWen,rhs_.io_diffCommits_info_184_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_184_fpWen!=rhs_.io_diffCommits_info_184_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_184_fpWen=0x%0h while the rhs_.io_diffCommits_info_184_fpWen=0x%0h",this.io_diffCommits_info_184_fpWen,rhs_.io_diffCommits_info_184_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_184_vecWen!=rhs_.io_diffCommits_info_184_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_184_vecWen=0x%0h while the rhs_.io_diffCommits_info_184_vecWen=0x%0h",this.io_diffCommits_info_184_vecWen,rhs_.io_diffCommits_info_184_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_184_v0Wen!=rhs_.io_diffCommits_info_184_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_184_v0Wen=0x%0h while the rhs_.io_diffCommits_info_184_v0Wen=0x%0h",this.io_diffCommits_info_184_v0Wen,rhs_.io_diffCommits_info_184_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_184_vlWen!=rhs_.io_diffCommits_info_184_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_184_vlWen=0x%0h while the rhs_.io_diffCommits_info_184_vlWen=0x%0h",this.io_diffCommits_info_184_vlWen,rhs_.io_diffCommits_info_184_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_185_ldest!=rhs_.io_diffCommits_info_185_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_185_ldest=0x%0h while the rhs_.io_diffCommits_info_185_ldest=0x%0h",this.io_diffCommits_info_185_ldest,rhs_.io_diffCommits_info_185_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_185_pdest!=rhs_.io_diffCommits_info_185_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_185_pdest=0x%0h while the rhs_.io_diffCommits_info_185_pdest=0x%0h",this.io_diffCommits_info_185_pdest,rhs_.io_diffCommits_info_185_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_185_rfWen!=rhs_.io_diffCommits_info_185_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_185_rfWen=0x%0h while the rhs_.io_diffCommits_info_185_rfWen=0x%0h",this.io_diffCommits_info_185_rfWen,rhs_.io_diffCommits_info_185_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_185_fpWen!=rhs_.io_diffCommits_info_185_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_185_fpWen=0x%0h while the rhs_.io_diffCommits_info_185_fpWen=0x%0h",this.io_diffCommits_info_185_fpWen,rhs_.io_diffCommits_info_185_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_185_vecWen!=rhs_.io_diffCommits_info_185_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_185_vecWen=0x%0h while the rhs_.io_diffCommits_info_185_vecWen=0x%0h",this.io_diffCommits_info_185_vecWen,rhs_.io_diffCommits_info_185_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_185_v0Wen!=rhs_.io_diffCommits_info_185_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_185_v0Wen=0x%0h while the rhs_.io_diffCommits_info_185_v0Wen=0x%0h",this.io_diffCommits_info_185_v0Wen,rhs_.io_diffCommits_info_185_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_185_vlWen!=rhs_.io_diffCommits_info_185_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_185_vlWen=0x%0h while the rhs_.io_diffCommits_info_185_vlWen=0x%0h",this.io_diffCommits_info_185_vlWen,rhs_.io_diffCommits_info_185_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_186_ldest!=rhs_.io_diffCommits_info_186_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_186_ldest=0x%0h while the rhs_.io_diffCommits_info_186_ldest=0x%0h",this.io_diffCommits_info_186_ldest,rhs_.io_diffCommits_info_186_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_186_pdest!=rhs_.io_diffCommits_info_186_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_186_pdest=0x%0h while the rhs_.io_diffCommits_info_186_pdest=0x%0h",this.io_diffCommits_info_186_pdest,rhs_.io_diffCommits_info_186_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_186_rfWen!=rhs_.io_diffCommits_info_186_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_186_rfWen=0x%0h while the rhs_.io_diffCommits_info_186_rfWen=0x%0h",this.io_diffCommits_info_186_rfWen,rhs_.io_diffCommits_info_186_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_186_fpWen!=rhs_.io_diffCommits_info_186_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_186_fpWen=0x%0h while the rhs_.io_diffCommits_info_186_fpWen=0x%0h",this.io_diffCommits_info_186_fpWen,rhs_.io_diffCommits_info_186_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_186_vecWen!=rhs_.io_diffCommits_info_186_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_186_vecWen=0x%0h while the rhs_.io_diffCommits_info_186_vecWen=0x%0h",this.io_diffCommits_info_186_vecWen,rhs_.io_diffCommits_info_186_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_186_v0Wen!=rhs_.io_diffCommits_info_186_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_186_v0Wen=0x%0h while the rhs_.io_diffCommits_info_186_v0Wen=0x%0h",this.io_diffCommits_info_186_v0Wen,rhs_.io_diffCommits_info_186_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_186_vlWen!=rhs_.io_diffCommits_info_186_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_186_vlWen=0x%0h while the rhs_.io_diffCommits_info_186_vlWen=0x%0h",this.io_diffCommits_info_186_vlWen,rhs_.io_diffCommits_info_186_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_187_ldest!=rhs_.io_diffCommits_info_187_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_187_ldest=0x%0h while the rhs_.io_diffCommits_info_187_ldest=0x%0h",this.io_diffCommits_info_187_ldest,rhs_.io_diffCommits_info_187_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_187_pdest!=rhs_.io_diffCommits_info_187_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_187_pdest=0x%0h while the rhs_.io_diffCommits_info_187_pdest=0x%0h",this.io_diffCommits_info_187_pdest,rhs_.io_diffCommits_info_187_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_187_rfWen!=rhs_.io_diffCommits_info_187_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_187_rfWen=0x%0h while the rhs_.io_diffCommits_info_187_rfWen=0x%0h",this.io_diffCommits_info_187_rfWen,rhs_.io_diffCommits_info_187_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_187_fpWen!=rhs_.io_diffCommits_info_187_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_187_fpWen=0x%0h while the rhs_.io_diffCommits_info_187_fpWen=0x%0h",this.io_diffCommits_info_187_fpWen,rhs_.io_diffCommits_info_187_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_187_vecWen!=rhs_.io_diffCommits_info_187_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_187_vecWen=0x%0h while the rhs_.io_diffCommits_info_187_vecWen=0x%0h",this.io_diffCommits_info_187_vecWen,rhs_.io_diffCommits_info_187_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_187_v0Wen!=rhs_.io_diffCommits_info_187_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_187_v0Wen=0x%0h while the rhs_.io_diffCommits_info_187_v0Wen=0x%0h",this.io_diffCommits_info_187_v0Wen,rhs_.io_diffCommits_info_187_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_187_vlWen!=rhs_.io_diffCommits_info_187_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_187_vlWen=0x%0h while the rhs_.io_diffCommits_info_187_vlWen=0x%0h",this.io_diffCommits_info_187_vlWen,rhs_.io_diffCommits_info_187_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_188_ldest!=rhs_.io_diffCommits_info_188_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_188_ldest=0x%0h while the rhs_.io_diffCommits_info_188_ldest=0x%0h",this.io_diffCommits_info_188_ldest,rhs_.io_diffCommits_info_188_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_188_pdest!=rhs_.io_diffCommits_info_188_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_188_pdest=0x%0h while the rhs_.io_diffCommits_info_188_pdest=0x%0h",this.io_diffCommits_info_188_pdest,rhs_.io_diffCommits_info_188_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_188_rfWen!=rhs_.io_diffCommits_info_188_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_188_rfWen=0x%0h while the rhs_.io_diffCommits_info_188_rfWen=0x%0h",this.io_diffCommits_info_188_rfWen,rhs_.io_diffCommits_info_188_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_188_fpWen!=rhs_.io_diffCommits_info_188_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_188_fpWen=0x%0h while the rhs_.io_diffCommits_info_188_fpWen=0x%0h",this.io_diffCommits_info_188_fpWen,rhs_.io_diffCommits_info_188_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_188_vecWen!=rhs_.io_diffCommits_info_188_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_188_vecWen=0x%0h while the rhs_.io_diffCommits_info_188_vecWen=0x%0h",this.io_diffCommits_info_188_vecWen,rhs_.io_diffCommits_info_188_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_188_v0Wen!=rhs_.io_diffCommits_info_188_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_188_v0Wen=0x%0h while the rhs_.io_diffCommits_info_188_v0Wen=0x%0h",this.io_diffCommits_info_188_v0Wen,rhs_.io_diffCommits_info_188_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_188_vlWen!=rhs_.io_diffCommits_info_188_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_188_vlWen=0x%0h while the rhs_.io_diffCommits_info_188_vlWen=0x%0h",this.io_diffCommits_info_188_vlWen,rhs_.io_diffCommits_info_188_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_189_ldest!=rhs_.io_diffCommits_info_189_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_189_ldest=0x%0h while the rhs_.io_diffCommits_info_189_ldest=0x%0h",this.io_diffCommits_info_189_ldest,rhs_.io_diffCommits_info_189_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_189_pdest!=rhs_.io_diffCommits_info_189_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_189_pdest=0x%0h while the rhs_.io_diffCommits_info_189_pdest=0x%0h",this.io_diffCommits_info_189_pdest,rhs_.io_diffCommits_info_189_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_189_rfWen!=rhs_.io_diffCommits_info_189_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_189_rfWen=0x%0h while the rhs_.io_diffCommits_info_189_rfWen=0x%0h",this.io_diffCommits_info_189_rfWen,rhs_.io_diffCommits_info_189_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_189_fpWen!=rhs_.io_diffCommits_info_189_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_189_fpWen=0x%0h while the rhs_.io_diffCommits_info_189_fpWen=0x%0h",this.io_diffCommits_info_189_fpWen,rhs_.io_diffCommits_info_189_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_189_vecWen!=rhs_.io_diffCommits_info_189_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_189_vecWen=0x%0h while the rhs_.io_diffCommits_info_189_vecWen=0x%0h",this.io_diffCommits_info_189_vecWen,rhs_.io_diffCommits_info_189_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_189_v0Wen!=rhs_.io_diffCommits_info_189_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_189_v0Wen=0x%0h while the rhs_.io_diffCommits_info_189_v0Wen=0x%0h",this.io_diffCommits_info_189_v0Wen,rhs_.io_diffCommits_info_189_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_189_vlWen!=rhs_.io_diffCommits_info_189_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_189_vlWen=0x%0h while the rhs_.io_diffCommits_info_189_vlWen=0x%0h",this.io_diffCommits_info_189_vlWen,rhs_.io_diffCommits_info_189_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_190_ldest!=rhs_.io_diffCommits_info_190_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_190_ldest=0x%0h while the rhs_.io_diffCommits_info_190_ldest=0x%0h",this.io_diffCommits_info_190_ldest,rhs_.io_diffCommits_info_190_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_190_pdest!=rhs_.io_diffCommits_info_190_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_190_pdest=0x%0h while the rhs_.io_diffCommits_info_190_pdest=0x%0h",this.io_diffCommits_info_190_pdest,rhs_.io_diffCommits_info_190_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_190_rfWen!=rhs_.io_diffCommits_info_190_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_190_rfWen=0x%0h while the rhs_.io_diffCommits_info_190_rfWen=0x%0h",this.io_diffCommits_info_190_rfWen,rhs_.io_diffCommits_info_190_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_190_fpWen!=rhs_.io_diffCommits_info_190_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_190_fpWen=0x%0h while the rhs_.io_diffCommits_info_190_fpWen=0x%0h",this.io_diffCommits_info_190_fpWen,rhs_.io_diffCommits_info_190_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_190_vecWen!=rhs_.io_diffCommits_info_190_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_190_vecWen=0x%0h while the rhs_.io_diffCommits_info_190_vecWen=0x%0h",this.io_diffCommits_info_190_vecWen,rhs_.io_diffCommits_info_190_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_190_v0Wen!=rhs_.io_diffCommits_info_190_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_190_v0Wen=0x%0h while the rhs_.io_diffCommits_info_190_v0Wen=0x%0h",this.io_diffCommits_info_190_v0Wen,rhs_.io_diffCommits_info_190_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_190_vlWen!=rhs_.io_diffCommits_info_190_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_190_vlWen=0x%0h while the rhs_.io_diffCommits_info_190_vlWen=0x%0h",this.io_diffCommits_info_190_vlWen,rhs_.io_diffCommits_info_190_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_191_ldest!=rhs_.io_diffCommits_info_191_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_191_ldest=0x%0h while the rhs_.io_diffCommits_info_191_ldest=0x%0h",this.io_diffCommits_info_191_ldest,rhs_.io_diffCommits_info_191_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_191_pdest!=rhs_.io_diffCommits_info_191_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_191_pdest=0x%0h while the rhs_.io_diffCommits_info_191_pdest=0x%0h",this.io_diffCommits_info_191_pdest,rhs_.io_diffCommits_info_191_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_191_rfWen!=rhs_.io_diffCommits_info_191_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_191_rfWen=0x%0h while the rhs_.io_diffCommits_info_191_rfWen=0x%0h",this.io_diffCommits_info_191_rfWen,rhs_.io_diffCommits_info_191_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_191_fpWen!=rhs_.io_diffCommits_info_191_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_191_fpWen=0x%0h while the rhs_.io_diffCommits_info_191_fpWen=0x%0h",this.io_diffCommits_info_191_fpWen,rhs_.io_diffCommits_info_191_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_191_vecWen!=rhs_.io_diffCommits_info_191_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_191_vecWen=0x%0h while the rhs_.io_diffCommits_info_191_vecWen=0x%0h",this.io_diffCommits_info_191_vecWen,rhs_.io_diffCommits_info_191_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_191_v0Wen!=rhs_.io_diffCommits_info_191_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_191_v0Wen=0x%0h while the rhs_.io_diffCommits_info_191_v0Wen=0x%0h",this.io_diffCommits_info_191_v0Wen,rhs_.io_diffCommits_info_191_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_191_vlWen!=rhs_.io_diffCommits_info_191_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_191_vlWen=0x%0h while the rhs_.io_diffCommits_info_191_vlWen=0x%0h",this.io_diffCommits_info_191_vlWen,rhs_.io_diffCommits_info_191_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_192_ldest!=rhs_.io_diffCommits_info_192_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_192_ldest=0x%0h while the rhs_.io_diffCommits_info_192_ldest=0x%0h",this.io_diffCommits_info_192_ldest,rhs_.io_diffCommits_info_192_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_192_pdest!=rhs_.io_diffCommits_info_192_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_192_pdest=0x%0h while the rhs_.io_diffCommits_info_192_pdest=0x%0h",this.io_diffCommits_info_192_pdest,rhs_.io_diffCommits_info_192_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_192_rfWen!=rhs_.io_diffCommits_info_192_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_192_rfWen=0x%0h while the rhs_.io_diffCommits_info_192_rfWen=0x%0h",this.io_diffCommits_info_192_rfWen,rhs_.io_diffCommits_info_192_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_192_fpWen!=rhs_.io_diffCommits_info_192_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_192_fpWen=0x%0h while the rhs_.io_diffCommits_info_192_fpWen=0x%0h",this.io_diffCommits_info_192_fpWen,rhs_.io_diffCommits_info_192_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_192_vecWen!=rhs_.io_diffCommits_info_192_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_192_vecWen=0x%0h while the rhs_.io_diffCommits_info_192_vecWen=0x%0h",this.io_diffCommits_info_192_vecWen,rhs_.io_diffCommits_info_192_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_192_v0Wen!=rhs_.io_diffCommits_info_192_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_192_v0Wen=0x%0h while the rhs_.io_diffCommits_info_192_v0Wen=0x%0h",this.io_diffCommits_info_192_v0Wen,rhs_.io_diffCommits_info_192_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_192_vlWen!=rhs_.io_diffCommits_info_192_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_192_vlWen=0x%0h while the rhs_.io_diffCommits_info_192_vlWen=0x%0h",this.io_diffCommits_info_192_vlWen,rhs_.io_diffCommits_info_192_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_193_ldest!=rhs_.io_diffCommits_info_193_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_193_ldest=0x%0h while the rhs_.io_diffCommits_info_193_ldest=0x%0h",this.io_diffCommits_info_193_ldest,rhs_.io_diffCommits_info_193_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_193_pdest!=rhs_.io_diffCommits_info_193_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_193_pdest=0x%0h while the rhs_.io_diffCommits_info_193_pdest=0x%0h",this.io_diffCommits_info_193_pdest,rhs_.io_diffCommits_info_193_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_193_rfWen!=rhs_.io_diffCommits_info_193_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_193_rfWen=0x%0h while the rhs_.io_diffCommits_info_193_rfWen=0x%0h",this.io_diffCommits_info_193_rfWen,rhs_.io_diffCommits_info_193_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_193_fpWen!=rhs_.io_diffCommits_info_193_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_193_fpWen=0x%0h while the rhs_.io_diffCommits_info_193_fpWen=0x%0h",this.io_diffCommits_info_193_fpWen,rhs_.io_diffCommits_info_193_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_193_vecWen!=rhs_.io_diffCommits_info_193_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_193_vecWen=0x%0h while the rhs_.io_diffCommits_info_193_vecWen=0x%0h",this.io_diffCommits_info_193_vecWen,rhs_.io_diffCommits_info_193_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_193_v0Wen!=rhs_.io_diffCommits_info_193_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_193_v0Wen=0x%0h while the rhs_.io_diffCommits_info_193_v0Wen=0x%0h",this.io_diffCommits_info_193_v0Wen,rhs_.io_diffCommits_info_193_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_193_vlWen!=rhs_.io_diffCommits_info_193_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_193_vlWen=0x%0h while the rhs_.io_diffCommits_info_193_vlWen=0x%0h",this.io_diffCommits_info_193_vlWen,rhs_.io_diffCommits_info_193_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_194_ldest!=rhs_.io_diffCommits_info_194_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_194_ldest=0x%0h while the rhs_.io_diffCommits_info_194_ldest=0x%0h",this.io_diffCommits_info_194_ldest,rhs_.io_diffCommits_info_194_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_194_pdest!=rhs_.io_diffCommits_info_194_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_194_pdest=0x%0h while the rhs_.io_diffCommits_info_194_pdest=0x%0h",this.io_diffCommits_info_194_pdest,rhs_.io_diffCommits_info_194_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_194_rfWen!=rhs_.io_diffCommits_info_194_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_194_rfWen=0x%0h while the rhs_.io_diffCommits_info_194_rfWen=0x%0h",this.io_diffCommits_info_194_rfWen,rhs_.io_diffCommits_info_194_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_194_fpWen!=rhs_.io_diffCommits_info_194_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_194_fpWen=0x%0h while the rhs_.io_diffCommits_info_194_fpWen=0x%0h",this.io_diffCommits_info_194_fpWen,rhs_.io_diffCommits_info_194_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_194_vecWen!=rhs_.io_diffCommits_info_194_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_194_vecWen=0x%0h while the rhs_.io_diffCommits_info_194_vecWen=0x%0h",this.io_diffCommits_info_194_vecWen,rhs_.io_diffCommits_info_194_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_194_v0Wen!=rhs_.io_diffCommits_info_194_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_194_v0Wen=0x%0h while the rhs_.io_diffCommits_info_194_v0Wen=0x%0h",this.io_diffCommits_info_194_v0Wen,rhs_.io_diffCommits_info_194_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_194_vlWen!=rhs_.io_diffCommits_info_194_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_194_vlWen=0x%0h while the rhs_.io_diffCommits_info_194_vlWen=0x%0h",this.io_diffCommits_info_194_vlWen,rhs_.io_diffCommits_info_194_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_195_ldest!=rhs_.io_diffCommits_info_195_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_195_ldest=0x%0h while the rhs_.io_diffCommits_info_195_ldest=0x%0h",this.io_diffCommits_info_195_ldest,rhs_.io_diffCommits_info_195_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_195_pdest!=rhs_.io_diffCommits_info_195_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_195_pdest=0x%0h while the rhs_.io_diffCommits_info_195_pdest=0x%0h",this.io_diffCommits_info_195_pdest,rhs_.io_diffCommits_info_195_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_195_rfWen!=rhs_.io_diffCommits_info_195_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_195_rfWen=0x%0h while the rhs_.io_diffCommits_info_195_rfWen=0x%0h",this.io_diffCommits_info_195_rfWen,rhs_.io_diffCommits_info_195_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_195_fpWen!=rhs_.io_diffCommits_info_195_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_195_fpWen=0x%0h while the rhs_.io_diffCommits_info_195_fpWen=0x%0h",this.io_diffCommits_info_195_fpWen,rhs_.io_diffCommits_info_195_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_195_vecWen!=rhs_.io_diffCommits_info_195_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_195_vecWen=0x%0h while the rhs_.io_diffCommits_info_195_vecWen=0x%0h",this.io_diffCommits_info_195_vecWen,rhs_.io_diffCommits_info_195_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_195_v0Wen!=rhs_.io_diffCommits_info_195_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_195_v0Wen=0x%0h while the rhs_.io_diffCommits_info_195_v0Wen=0x%0h",this.io_diffCommits_info_195_v0Wen,rhs_.io_diffCommits_info_195_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_195_vlWen!=rhs_.io_diffCommits_info_195_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_195_vlWen=0x%0h while the rhs_.io_diffCommits_info_195_vlWen=0x%0h",this.io_diffCommits_info_195_vlWen,rhs_.io_diffCommits_info_195_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_196_ldest!=rhs_.io_diffCommits_info_196_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_196_ldest=0x%0h while the rhs_.io_diffCommits_info_196_ldest=0x%0h",this.io_diffCommits_info_196_ldest,rhs_.io_diffCommits_info_196_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_196_pdest!=rhs_.io_diffCommits_info_196_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_196_pdest=0x%0h while the rhs_.io_diffCommits_info_196_pdest=0x%0h",this.io_diffCommits_info_196_pdest,rhs_.io_diffCommits_info_196_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_196_rfWen!=rhs_.io_diffCommits_info_196_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_196_rfWen=0x%0h while the rhs_.io_diffCommits_info_196_rfWen=0x%0h",this.io_diffCommits_info_196_rfWen,rhs_.io_diffCommits_info_196_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_196_fpWen!=rhs_.io_diffCommits_info_196_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_196_fpWen=0x%0h while the rhs_.io_diffCommits_info_196_fpWen=0x%0h",this.io_diffCommits_info_196_fpWen,rhs_.io_diffCommits_info_196_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_196_vecWen!=rhs_.io_diffCommits_info_196_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_196_vecWen=0x%0h while the rhs_.io_diffCommits_info_196_vecWen=0x%0h",this.io_diffCommits_info_196_vecWen,rhs_.io_diffCommits_info_196_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_196_v0Wen!=rhs_.io_diffCommits_info_196_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_196_v0Wen=0x%0h while the rhs_.io_diffCommits_info_196_v0Wen=0x%0h",this.io_diffCommits_info_196_v0Wen,rhs_.io_diffCommits_info_196_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_196_vlWen!=rhs_.io_diffCommits_info_196_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_196_vlWen=0x%0h while the rhs_.io_diffCommits_info_196_vlWen=0x%0h",this.io_diffCommits_info_196_vlWen,rhs_.io_diffCommits_info_196_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_197_ldest!=rhs_.io_diffCommits_info_197_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_197_ldest=0x%0h while the rhs_.io_diffCommits_info_197_ldest=0x%0h",this.io_diffCommits_info_197_ldest,rhs_.io_diffCommits_info_197_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_197_pdest!=rhs_.io_diffCommits_info_197_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_197_pdest=0x%0h while the rhs_.io_diffCommits_info_197_pdest=0x%0h",this.io_diffCommits_info_197_pdest,rhs_.io_diffCommits_info_197_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_197_rfWen!=rhs_.io_diffCommits_info_197_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_197_rfWen=0x%0h while the rhs_.io_diffCommits_info_197_rfWen=0x%0h",this.io_diffCommits_info_197_rfWen,rhs_.io_diffCommits_info_197_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_197_fpWen!=rhs_.io_diffCommits_info_197_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_197_fpWen=0x%0h while the rhs_.io_diffCommits_info_197_fpWen=0x%0h",this.io_diffCommits_info_197_fpWen,rhs_.io_diffCommits_info_197_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_197_vecWen!=rhs_.io_diffCommits_info_197_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_197_vecWen=0x%0h while the rhs_.io_diffCommits_info_197_vecWen=0x%0h",this.io_diffCommits_info_197_vecWen,rhs_.io_diffCommits_info_197_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_197_v0Wen!=rhs_.io_diffCommits_info_197_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_197_v0Wen=0x%0h while the rhs_.io_diffCommits_info_197_v0Wen=0x%0h",this.io_diffCommits_info_197_v0Wen,rhs_.io_diffCommits_info_197_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_197_vlWen!=rhs_.io_diffCommits_info_197_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_197_vlWen=0x%0h while the rhs_.io_diffCommits_info_197_vlWen=0x%0h",this.io_diffCommits_info_197_vlWen,rhs_.io_diffCommits_info_197_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_198_ldest!=rhs_.io_diffCommits_info_198_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_198_ldest=0x%0h while the rhs_.io_diffCommits_info_198_ldest=0x%0h",this.io_diffCommits_info_198_ldest,rhs_.io_diffCommits_info_198_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_198_pdest!=rhs_.io_diffCommits_info_198_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_198_pdest=0x%0h while the rhs_.io_diffCommits_info_198_pdest=0x%0h",this.io_diffCommits_info_198_pdest,rhs_.io_diffCommits_info_198_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_198_rfWen!=rhs_.io_diffCommits_info_198_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_198_rfWen=0x%0h while the rhs_.io_diffCommits_info_198_rfWen=0x%0h",this.io_diffCommits_info_198_rfWen,rhs_.io_diffCommits_info_198_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_198_fpWen!=rhs_.io_diffCommits_info_198_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_198_fpWen=0x%0h while the rhs_.io_diffCommits_info_198_fpWen=0x%0h",this.io_diffCommits_info_198_fpWen,rhs_.io_diffCommits_info_198_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_198_vecWen!=rhs_.io_diffCommits_info_198_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_198_vecWen=0x%0h while the rhs_.io_diffCommits_info_198_vecWen=0x%0h",this.io_diffCommits_info_198_vecWen,rhs_.io_diffCommits_info_198_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_198_v0Wen!=rhs_.io_diffCommits_info_198_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_198_v0Wen=0x%0h while the rhs_.io_diffCommits_info_198_v0Wen=0x%0h",this.io_diffCommits_info_198_v0Wen,rhs_.io_diffCommits_info_198_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_198_vlWen!=rhs_.io_diffCommits_info_198_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_198_vlWen=0x%0h while the rhs_.io_diffCommits_info_198_vlWen=0x%0h",this.io_diffCommits_info_198_vlWen,rhs_.io_diffCommits_info_198_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_199_ldest!=rhs_.io_diffCommits_info_199_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_199_ldest=0x%0h while the rhs_.io_diffCommits_info_199_ldest=0x%0h",this.io_diffCommits_info_199_ldest,rhs_.io_diffCommits_info_199_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_199_pdest!=rhs_.io_diffCommits_info_199_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_199_pdest=0x%0h while the rhs_.io_diffCommits_info_199_pdest=0x%0h",this.io_diffCommits_info_199_pdest,rhs_.io_diffCommits_info_199_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_199_rfWen!=rhs_.io_diffCommits_info_199_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_199_rfWen=0x%0h while the rhs_.io_diffCommits_info_199_rfWen=0x%0h",this.io_diffCommits_info_199_rfWen,rhs_.io_diffCommits_info_199_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_199_fpWen!=rhs_.io_diffCommits_info_199_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_199_fpWen=0x%0h while the rhs_.io_diffCommits_info_199_fpWen=0x%0h",this.io_diffCommits_info_199_fpWen,rhs_.io_diffCommits_info_199_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_199_vecWen!=rhs_.io_diffCommits_info_199_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_199_vecWen=0x%0h while the rhs_.io_diffCommits_info_199_vecWen=0x%0h",this.io_diffCommits_info_199_vecWen,rhs_.io_diffCommits_info_199_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_199_v0Wen!=rhs_.io_diffCommits_info_199_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_199_v0Wen=0x%0h while the rhs_.io_diffCommits_info_199_v0Wen=0x%0h",this.io_diffCommits_info_199_v0Wen,rhs_.io_diffCommits_info_199_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_199_vlWen!=rhs_.io_diffCommits_info_199_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_199_vlWen=0x%0h while the rhs_.io_diffCommits_info_199_vlWen=0x%0h",this.io_diffCommits_info_199_vlWen,rhs_.io_diffCommits_info_199_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_200_ldest!=rhs_.io_diffCommits_info_200_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_200_ldest=0x%0h while the rhs_.io_diffCommits_info_200_ldest=0x%0h",this.io_diffCommits_info_200_ldest,rhs_.io_diffCommits_info_200_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_200_pdest!=rhs_.io_diffCommits_info_200_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_200_pdest=0x%0h while the rhs_.io_diffCommits_info_200_pdest=0x%0h",this.io_diffCommits_info_200_pdest,rhs_.io_diffCommits_info_200_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_200_rfWen!=rhs_.io_diffCommits_info_200_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_200_rfWen=0x%0h while the rhs_.io_diffCommits_info_200_rfWen=0x%0h",this.io_diffCommits_info_200_rfWen,rhs_.io_diffCommits_info_200_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_200_fpWen!=rhs_.io_diffCommits_info_200_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_200_fpWen=0x%0h while the rhs_.io_diffCommits_info_200_fpWen=0x%0h",this.io_diffCommits_info_200_fpWen,rhs_.io_diffCommits_info_200_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_200_vecWen!=rhs_.io_diffCommits_info_200_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_200_vecWen=0x%0h while the rhs_.io_diffCommits_info_200_vecWen=0x%0h",this.io_diffCommits_info_200_vecWen,rhs_.io_diffCommits_info_200_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_200_v0Wen!=rhs_.io_diffCommits_info_200_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_200_v0Wen=0x%0h while the rhs_.io_diffCommits_info_200_v0Wen=0x%0h",this.io_diffCommits_info_200_v0Wen,rhs_.io_diffCommits_info_200_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_200_vlWen!=rhs_.io_diffCommits_info_200_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_200_vlWen=0x%0h while the rhs_.io_diffCommits_info_200_vlWen=0x%0h",this.io_diffCommits_info_200_vlWen,rhs_.io_diffCommits_info_200_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_201_ldest!=rhs_.io_diffCommits_info_201_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_201_ldest=0x%0h while the rhs_.io_diffCommits_info_201_ldest=0x%0h",this.io_diffCommits_info_201_ldest,rhs_.io_diffCommits_info_201_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_201_pdest!=rhs_.io_diffCommits_info_201_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_201_pdest=0x%0h while the rhs_.io_diffCommits_info_201_pdest=0x%0h",this.io_diffCommits_info_201_pdest,rhs_.io_diffCommits_info_201_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_201_rfWen!=rhs_.io_diffCommits_info_201_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_201_rfWen=0x%0h while the rhs_.io_diffCommits_info_201_rfWen=0x%0h",this.io_diffCommits_info_201_rfWen,rhs_.io_diffCommits_info_201_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_201_fpWen!=rhs_.io_diffCommits_info_201_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_201_fpWen=0x%0h while the rhs_.io_diffCommits_info_201_fpWen=0x%0h",this.io_diffCommits_info_201_fpWen,rhs_.io_diffCommits_info_201_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_201_vecWen!=rhs_.io_diffCommits_info_201_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_201_vecWen=0x%0h while the rhs_.io_diffCommits_info_201_vecWen=0x%0h",this.io_diffCommits_info_201_vecWen,rhs_.io_diffCommits_info_201_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_201_v0Wen!=rhs_.io_diffCommits_info_201_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_201_v0Wen=0x%0h while the rhs_.io_diffCommits_info_201_v0Wen=0x%0h",this.io_diffCommits_info_201_v0Wen,rhs_.io_diffCommits_info_201_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_201_vlWen!=rhs_.io_diffCommits_info_201_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_201_vlWen=0x%0h while the rhs_.io_diffCommits_info_201_vlWen=0x%0h",this.io_diffCommits_info_201_vlWen,rhs_.io_diffCommits_info_201_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_202_ldest!=rhs_.io_diffCommits_info_202_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_202_ldest=0x%0h while the rhs_.io_diffCommits_info_202_ldest=0x%0h",this.io_diffCommits_info_202_ldest,rhs_.io_diffCommits_info_202_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_202_pdest!=rhs_.io_diffCommits_info_202_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_202_pdest=0x%0h while the rhs_.io_diffCommits_info_202_pdest=0x%0h",this.io_diffCommits_info_202_pdest,rhs_.io_diffCommits_info_202_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_202_rfWen!=rhs_.io_diffCommits_info_202_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_202_rfWen=0x%0h while the rhs_.io_diffCommits_info_202_rfWen=0x%0h",this.io_diffCommits_info_202_rfWen,rhs_.io_diffCommits_info_202_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_202_fpWen!=rhs_.io_diffCommits_info_202_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_202_fpWen=0x%0h while the rhs_.io_diffCommits_info_202_fpWen=0x%0h",this.io_diffCommits_info_202_fpWen,rhs_.io_diffCommits_info_202_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_202_vecWen!=rhs_.io_diffCommits_info_202_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_202_vecWen=0x%0h while the rhs_.io_diffCommits_info_202_vecWen=0x%0h",this.io_diffCommits_info_202_vecWen,rhs_.io_diffCommits_info_202_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_202_v0Wen!=rhs_.io_diffCommits_info_202_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_202_v0Wen=0x%0h while the rhs_.io_diffCommits_info_202_v0Wen=0x%0h",this.io_diffCommits_info_202_v0Wen,rhs_.io_diffCommits_info_202_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_202_vlWen!=rhs_.io_diffCommits_info_202_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_202_vlWen=0x%0h while the rhs_.io_diffCommits_info_202_vlWen=0x%0h",this.io_diffCommits_info_202_vlWen,rhs_.io_diffCommits_info_202_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_203_ldest!=rhs_.io_diffCommits_info_203_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_203_ldest=0x%0h while the rhs_.io_diffCommits_info_203_ldest=0x%0h",this.io_diffCommits_info_203_ldest,rhs_.io_diffCommits_info_203_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_203_pdest!=rhs_.io_diffCommits_info_203_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_203_pdest=0x%0h while the rhs_.io_diffCommits_info_203_pdest=0x%0h",this.io_diffCommits_info_203_pdest,rhs_.io_diffCommits_info_203_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_203_rfWen!=rhs_.io_diffCommits_info_203_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_203_rfWen=0x%0h while the rhs_.io_diffCommits_info_203_rfWen=0x%0h",this.io_diffCommits_info_203_rfWen,rhs_.io_diffCommits_info_203_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_203_fpWen!=rhs_.io_diffCommits_info_203_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_203_fpWen=0x%0h while the rhs_.io_diffCommits_info_203_fpWen=0x%0h",this.io_diffCommits_info_203_fpWen,rhs_.io_diffCommits_info_203_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_203_vecWen!=rhs_.io_diffCommits_info_203_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_203_vecWen=0x%0h while the rhs_.io_diffCommits_info_203_vecWen=0x%0h",this.io_diffCommits_info_203_vecWen,rhs_.io_diffCommits_info_203_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_203_v0Wen!=rhs_.io_diffCommits_info_203_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_203_v0Wen=0x%0h while the rhs_.io_diffCommits_info_203_v0Wen=0x%0h",this.io_diffCommits_info_203_v0Wen,rhs_.io_diffCommits_info_203_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_203_vlWen!=rhs_.io_diffCommits_info_203_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_203_vlWen=0x%0h while the rhs_.io_diffCommits_info_203_vlWen=0x%0h",this.io_diffCommits_info_203_vlWen,rhs_.io_diffCommits_info_203_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_204_ldest!=rhs_.io_diffCommits_info_204_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_204_ldest=0x%0h while the rhs_.io_diffCommits_info_204_ldest=0x%0h",this.io_diffCommits_info_204_ldest,rhs_.io_diffCommits_info_204_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_204_pdest!=rhs_.io_diffCommits_info_204_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_204_pdest=0x%0h while the rhs_.io_diffCommits_info_204_pdest=0x%0h",this.io_diffCommits_info_204_pdest,rhs_.io_diffCommits_info_204_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_204_rfWen!=rhs_.io_diffCommits_info_204_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_204_rfWen=0x%0h while the rhs_.io_diffCommits_info_204_rfWen=0x%0h",this.io_diffCommits_info_204_rfWen,rhs_.io_diffCommits_info_204_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_204_fpWen!=rhs_.io_diffCommits_info_204_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_204_fpWen=0x%0h while the rhs_.io_diffCommits_info_204_fpWen=0x%0h",this.io_diffCommits_info_204_fpWen,rhs_.io_diffCommits_info_204_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_204_vecWen!=rhs_.io_diffCommits_info_204_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_204_vecWen=0x%0h while the rhs_.io_diffCommits_info_204_vecWen=0x%0h",this.io_diffCommits_info_204_vecWen,rhs_.io_diffCommits_info_204_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_204_v0Wen!=rhs_.io_diffCommits_info_204_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_204_v0Wen=0x%0h while the rhs_.io_diffCommits_info_204_v0Wen=0x%0h",this.io_diffCommits_info_204_v0Wen,rhs_.io_diffCommits_info_204_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_204_vlWen!=rhs_.io_diffCommits_info_204_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_204_vlWen=0x%0h while the rhs_.io_diffCommits_info_204_vlWen=0x%0h",this.io_diffCommits_info_204_vlWen,rhs_.io_diffCommits_info_204_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_205_ldest!=rhs_.io_diffCommits_info_205_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_205_ldest=0x%0h while the rhs_.io_diffCommits_info_205_ldest=0x%0h",this.io_diffCommits_info_205_ldest,rhs_.io_diffCommits_info_205_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_205_pdest!=rhs_.io_diffCommits_info_205_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_205_pdest=0x%0h while the rhs_.io_diffCommits_info_205_pdest=0x%0h",this.io_diffCommits_info_205_pdest,rhs_.io_diffCommits_info_205_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_205_rfWen!=rhs_.io_diffCommits_info_205_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_205_rfWen=0x%0h while the rhs_.io_diffCommits_info_205_rfWen=0x%0h",this.io_diffCommits_info_205_rfWen,rhs_.io_diffCommits_info_205_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_205_fpWen!=rhs_.io_diffCommits_info_205_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_205_fpWen=0x%0h while the rhs_.io_diffCommits_info_205_fpWen=0x%0h",this.io_diffCommits_info_205_fpWen,rhs_.io_diffCommits_info_205_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_205_vecWen!=rhs_.io_diffCommits_info_205_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_205_vecWen=0x%0h while the rhs_.io_diffCommits_info_205_vecWen=0x%0h",this.io_diffCommits_info_205_vecWen,rhs_.io_diffCommits_info_205_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_205_v0Wen!=rhs_.io_diffCommits_info_205_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_205_v0Wen=0x%0h while the rhs_.io_diffCommits_info_205_v0Wen=0x%0h",this.io_diffCommits_info_205_v0Wen,rhs_.io_diffCommits_info_205_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_205_vlWen!=rhs_.io_diffCommits_info_205_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_205_vlWen=0x%0h while the rhs_.io_diffCommits_info_205_vlWen=0x%0h",this.io_diffCommits_info_205_vlWen,rhs_.io_diffCommits_info_205_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_206_ldest!=rhs_.io_diffCommits_info_206_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_206_ldest=0x%0h while the rhs_.io_diffCommits_info_206_ldest=0x%0h",this.io_diffCommits_info_206_ldest,rhs_.io_diffCommits_info_206_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_206_pdest!=rhs_.io_diffCommits_info_206_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_206_pdest=0x%0h while the rhs_.io_diffCommits_info_206_pdest=0x%0h",this.io_diffCommits_info_206_pdest,rhs_.io_diffCommits_info_206_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_206_rfWen!=rhs_.io_diffCommits_info_206_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_206_rfWen=0x%0h while the rhs_.io_diffCommits_info_206_rfWen=0x%0h",this.io_diffCommits_info_206_rfWen,rhs_.io_diffCommits_info_206_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_206_fpWen!=rhs_.io_diffCommits_info_206_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_206_fpWen=0x%0h while the rhs_.io_diffCommits_info_206_fpWen=0x%0h",this.io_diffCommits_info_206_fpWen,rhs_.io_diffCommits_info_206_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_206_vecWen!=rhs_.io_diffCommits_info_206_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_206_vecWen=0x%0h while the rhs_.io_diffCommits_info_206_vecWen=0x%0h",this.io_diffCommits_info_206_vecWen,rhs_.io_diffCommits_info_206_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_206_v0Wen!=rhs_.io_diffCommits_info_206_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_206_v0Wen=0x%0h while the rhs_.io_diffCommits_info_206_v0Wen=0x%0h",this.io_diffCommits_info_206_v0Wen,rhs_.io_diffCommits_info_206_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_206_vlWen!=rhs_.io_diffCommits_info_206_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_206_vlWen=0x%0h while the rhs_.io_diffCommits_info_206_vlWen=0x%0h",this.io_diffCommits_info_206_vlWen,rhs_.io_diffCommits_info_206_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_207_ldest!=rhs_.io_diffCommits_info_207_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_207_ldest=0x%0h while the rhs_.io_diffCommits_info_207_ldest=0x%0h",this.io_diffCommits_info_207_ldest,rhs_.io_diffCommits_info_207_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_207_pdest!=rhs_.io_diffCommits_info_207_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_207_pdest=0x%0h while the rhs_.io_diffCommits_info_207_pdest=0x%0h",this.io_diffCommits_info_207_pdest,rhs_.io_diffCommits_info_207_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_207_rfWen!=rhs_.io_diffCommits_info_207_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_207_rfWen=0x%0h while the rhs_.io_diffCommits_info_207_rfWen=0x%0h",this.io_diffCommits_info_207_rfWen,rhs_.io_diffCommits_info_207_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_207_fpWen!=rhs_.io_diffCommits_info_207_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_207_fpWen=0x%0h while the rhs_.io_diffCommits_info_207_fpWen=0x%0h",this.io_diffCommits_info_207_fpWen,rhs_.io_diffCommits_info_207_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_207_vecWen!=rhs_.io_diffCommits_info_207_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_207_vecWen=0x%0h while the rhs_.io_diffCommits_info_207_vecWen=0x%0h",this.io_diffCommits_info_207_vecWen,rhs_.io_diffCommits_info_207_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_207_v0Wen!=rhs_.io_diffCommits_info_207_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_207_v0Wen=0x%0h while the rhs_.io_diffCommits_info_207_v0Wen=0x%0h",this.io_diffCommits_info_207_v0Wen,rhs_.io_diffCommits_info_207_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_207_vlWen!=rhs_.io_diffCommits_info_207_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_207_vlWen=0x%0h while the rhs_.io_diffCommits_info_207_vlWen=0x%0h",this.io_diffCommits_info_207_vlWen,rhs_.io_diffCommits_info_207_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_208_ldest!=rhs_.io_diffCommits_info_208_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_208_ldest=0x%0h while the rhs_.io_diffCommits_info_208_ldest=0x%0h",this.io_diffCommits_info_208_ldest,rhs_.io_diffCommits_info_208_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_208_pdest!=rhs_.io_diffCommits_info_208_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_208_pdest=0x%0h while the rhs_.io_diffCommits_info_208_pdest=0x%0h",this.io_diffCommits_info_208_pdest,rhs_.io_diffCommits_info_208_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_208_rfWen!=rhs_.io_diffCommits_info_208_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_208_rfWen=0x%0h while the rhs_.io_diffCommits_info_208_rfWen=0x%0h",this.io_diffCommits_info_208_rfWen,rhs_.io_diffCommits_info_208_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_208_fpWen!=rhs_.io_diffCommits_info_208_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_208_fpWen=0x%0h while the rhs_.io_diffCommits_info_208_fpWen=0x%0h",this.io_diffCommits_info_208_fpWen,rhs_.io_diffCommits_info_208_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_208_vecWen!=rhs_.io_diffCommits_info_208_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_208_vecWen=0x%0h while the rhs_.io_diffCommits_info_208_vecWen=0x%0h",this.io_diffCommits_info_208_vecWen,rhs_.io_diffCommits_info_208_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_208_v0Wen!=rhs_.io_diffCommits_info_208_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_208_v0Wen=0x%0h while the rhs_.io_diffCommits_info_208_v0Wen=0x%0h",this.io_diffCommits_info_208_v0Wen,rhs_.io_diffCommits_info_208_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_208_vlWen!=rhs_.io_diffCommits_info_208_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_208_vlWen=0x%0h while the rhs_.io_diffCommits_info_208_vlWen=0x%0h",this.io_diffCommits_info_208_vlWen,rhs_.io_diffCommits_info_208_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_209_ldest!=rhs_.io_diffCommits_info_209_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_209_ldest=0x%0h while the rhs_.io_diffCommits_info_209_ldest=0x%0h",this.io_diffCommits_info_209_ldest,rhs_.io_diffCommits_info_209_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_209_pdest!=rhs_.io_diffCommits_info_209_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_209_pdest=0x%0h while the rhs_.io_diffCommits_info_209_pdest=0x%0h",this.io_diffCommits_info_209_pdest,rhs_.io_diffCommits_info_209_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_209_rfWen!=rhs_.io_diffCommits_info_209_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_209_rfWen=0x%0h while the rhs_.io_diffCommits_info_209_rfWen=0x%0h",this.io_diffCommits_info_209_rfWen,rhs_.io_diffCommits_info_209_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_209_fpWen!=rhs_.io_diffCommits_info_209_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_209_fpWen=0x%0h while the rhs_.io_diffCommits_info_209_fpWen=0x%0h",this.io_diffCommits_info_209_fpWen,rhs_.io_diffCommits_info_209_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_209_vecWen!=rhs_.io_diffCommits_info_209_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_209_vecWen=0x%0h while the rhs_.io_diffCommits_info_209_vecWen=0x%0h",this.io_diffCommits_info_209_vecWen,rhs_.io_diffCommits_info_209_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_209_v0Wen!=rhs_.io_diffCommits_info_209_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_209_v0Wen=0x%0h while the rhs_.io_diffCommits_info_209_v0Wen=0x%0h",this.io_diffCommits_info_209_v0Wen,rhs_.io_diffCommits_info_209_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_209_vlWen!=rhs_.io_diffCommits_info_209_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_209_vlWen=0x%0h while the rhs_.io_diffCommits_info_209_vlWen=0x%0h",this.io_diffCommits_info_209_vlWen,rhs_.io_diffCommits_info_209_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_210_ldest!=rhs_.io_diffCommits_info_210_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_210_ldest=0x%0h while the rhs_.io_diffCommits_info_210_ldest=0x%0h",this.io_diffCommits_info_210_ldest,rhs_.io_diffCommits_info_210_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_210_pdest!=rhs_.io_diffCommits_info_210_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_210_pdest=0x%0h while the rhs_.io_diffCommits_info_210_pdest=0x%0h",this.io_diffCommits_info_210_pdest,rhs_.io_diffCommits_info_210_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_210_rfWen!=rhs_.io_diffCommits_info_210_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_210_rfWen=0x%0h while the rhs_.io_diffCommits_info_210_rfWen=0x%0h",this.io_diffCommits_info_210_rfWen,rhs_.io_diffCommits_info_210_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_210_fpWen!=rhs_.io_diffCommits_info_210_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_210_fpWen=0x%0h while the rhs_.io_diffCommits_info_210_fpWen=0x%0h",this.io_diffCommits_info_210_fpWen,rhs_.io_diffCommits_info_210_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_210_vecWen!=rhs_.io_diffCommits_info_210_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_210_vecWen=0x%0h while the rhs_.io_diffCommits_info_210_vecWen=0x%0h",this.io_diffCommits_info_210_vecWen,rhs_.io_diffCommits_info_210_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_210_v0Wen!=rhs_.io_diffCommits_info_210_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_210_v0Wen=0x%0h while the rhs_.io_diffCommits_info_210_v0Wen=0x%0h",this.io_diffCommits_info_210_v0Wen,rhs_.io_diffCommits_info_210_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_210_vlWen!=rhs_.io_diffCommits_info_210_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_210_vlWen=0x%0h while the rhs_.io_diffCommits_info_210_vlWen=0x%0h",this.io_diffCommits_info_210_vlWen,rhs_.io_diffCommits_info_210_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_211_ldest!=rhs_.io_diffCommits_info_211_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_211_ldest=0x%0h while the rhs_.io_diffCommits_info_211_ldest=0x%0h",this.io_diffCommits_info_211_ldest,rhs_.io_diffCommits_info_211_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_211_pdest!=rhs_.io_diffCommits_info_211_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_211_pdest=0x%0h while the rhs_.io_diffCommits_info_211_pdest=0x%0h",this.io_diffCommits_info_211_pdest,rhs_.io_diffCommits_info_211_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_211_rfWen!=rhs_.io_diffCommits_info_211_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_211_rfWen=0x%0h while the rhs_.io_diffCommits_info_211_rfWen=0x%0h",this.io_diffCommits_info_211_rfWen,rhs_.io_diffCommits_info_211_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_211_fpWen!=rhs_.io_diffCommits_info_211_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_211_fpWen=0x%0h while the rhs_.io_diffCommits_info_211_fpWen=0x%0h",this.io_diffCommits_info_211_fpWen,rhs_.io_diffCommits_info_211_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_211_vecWen!=rhs_.io_diffCommits_info_211_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_211_vecWen=0x%0h while the rhs_.io_diffCommits_info_211_vecWen=0x%0h",this.io_diffCommits_info_211_vecWen,rhs_.io_diffCommits_info_211_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_211_v0Wen!=rhs_.io_diffCommits_info_211_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_211_v0Wen=0x%0h while the rhs_.io_diffCommits_info_211_v0Wen=0x%0h",this.io_diffCommits_info_211_v0Wen,rhs_.io_diffCommits_info_211_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_211_vlWen!=rhs_.io_diffCommits_info_211_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_211_vlWen=0x%0h while the rhs_.io_diffCommits_info_211_vlWen=0x%0h",this.io_diffCommits_info_211_vlWen,rhs_.io_diffCommits_info_211_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_212_ldest!=rhs_.io_diffCommits_info_212_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_212_ldest=0x%0h while the rhs_.io_diffCommits_info_212_ldest=0x%0h",this.io_diffCommits_info_212_ldest,rhs_.io_diffCommits_info_212_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_212_pdest!=rhs_.io_diffCommits_info_212_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_212_pdest=0x%0h while the rhs_.io_diffCommits_info_212_pdest=0x%0h",this.io_diffCommits_info_212_pdest,rhs_.io_diffCommits_info_212_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_212_rfWen!=rhs_.io_diffCommits_info_212_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_212_rfWen=0x%0h while the rhs_.io_diffCommits_info_212_rfWen=0x%0h",this.io_diffCommits_info_212_rfWen,rhs_.io_diffCommits_info_212_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_212_fpWen!=rhs_.io_diffCommits_info_212_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_212_fpWen=0x%0h while the rhs_.io_diffCommits_info_212_fpWen=0x%0h",this.io_diffCommits_info_212_fpWen,rhs_.io_diffCommits_info_212_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_212_vecWen!=rhs_.io_diffCommits_info_212_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_212_vecWen=0x%0h while the rhs_.io_diffCommits_info_212_vecWen=0x%0h",this.io_diffCommits_info_212_vecWen,rhs_.io_diffCommits_info_212_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_212_v0Wen!=rhs_.io_diffCommits_info_212_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_212_v0Wen=0x%0h while the rhs_.io_diffCommits_info_212_v0Wen=0x%0h",this.io_diffCommits_info_212_v0Wen,rhs_.io_diffCommits_info_212_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_212_vlWen!=rhs_.io_diffCommits_info_212_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_212_vlWen=0x%0h while the rhs_.io_diffCommits_info_212_vlWen=0x%0h",this.io_diffCommits_info_212_vlWen,rhs_.io_diffCommits_info_212_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_213_ldest!=rhs_.io_diffCommits_info_213_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_213_ldest=0x%0h while the rhs_.io_diffCommits_info_213_ldest=0x%0h",this.io_diffCommits_info_213_ldest,rhs_.io_diffCommits_info_213_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_213_pdest!=rhs_.io_diffCommits_info_213_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_213_pdest=0x%0h while the rhs_.io_diffCommits_info_213_pdest=0x%0h",this.io_diffCommits_info_213_pdest,rhs_.io_diffCommits_info_213_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_213_rfWen!=rhs_.io_diffCommits_info_213_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_213_rfWen=0x%0h while the rhs_.io_diffCommits_info_213_rfWen=0x%0h",this.io_diffCommits_info_213_rfWen,rhs_.io_diffCommits_info_213_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_213_fpWen!=rhs_.io_diffCommits_info_213_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_213_fpWen=0x%0h while the rhs_.io_diffCommits_info_213_fpWen=0x%0h",this.io_diffCommits_info_213_fpWen,rhs_.io_diffCommits_info_213_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_213_vecWen!=rhs_.io_diffCommits_info_213_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_213_vecWen=0x%0h while the rhs_.io_diffCommits_info_213_vecWen=0x%0h",this.io_diffCommits_info_213_vecWen,rhs_.io_diffCommits_info_213_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_213_v0Wen!=rhs_.io_diffCommits_info_213_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_213_v0Wen=0x%0h while the rhs_.io_diffCommits_info_213_v0Wen=0x%0h",this.io_diffCommits_info_213_v0Wen,rhs_.io_diffCommits_info_213_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_213_vlWen!=rhs_.io_diffCommits_info_213_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_213_vlWen=0x%0h while the rhs_.io_diffCommits_info_213_vlWen=0x%0h",this.io_diffCommits_info_213_vlWen,rhs_.io_diffCommits_info_213_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_214_ldest!=rhs_.io_diffCommits_info_214_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_214_ldest=0x%0h while the rhs_.io_diffCommits_info_214_ldest=0x%0h",this.io_diffCommits_info_214_ldest,rhs_.io_diffCommits_info_214_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_214_pdest!=rhs_.io_diffCommits_info_214_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_214_pdest=0x%0h while the rhs_.io_diffCommits_info_214_pdest=0x%0h",this.io_diffCommits_info_214_pdest,rhs_.io_diffCommits_info_214_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_214_rfWen!=rhs_.io_diffCommits_info_214_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_214_rfWen=0x%0h while the rhs_.io_diffCommits_info_214_rfWen=0x%0h",this.io_diffCommits_info_214_rfWen,rhs_.io_diffCommits_info_214_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_214_fpWen!=rhs_.io_diffCommits_info_214_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_214_fpWen=0x%0h while the rhs_.io_diffCommits_info_214_fpWen=0x%0h",this.io_diffCommits_info_214_fpWen,rhs_.io_diffCommits_info_214_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_214_vecWen!=rhs_.io_diffCommits_info_214_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_214_vecWen=0x%0h while the rhs_.io_diffCommits_info_214_vecWen=0x%0h",this.io_diffCommits_info_214_vecWen,rhs_.io_diffCommits_info_214_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_214_v0Wen!=rhs_.io_diffCommits_info_214_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_214_v0Wen=0x%0h while the rhs_.io_diffCommits_info_214_v0Wen=0x%0h",this.io_diffCommits_info_214_v0Wen,rhs_.io_diffCommits_info_214_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_214_vlWen!=rhs_.io_diffCommits_info_214_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_214_vlWen=0x%0h while the rhs_.io_diffCommits_info_214_vlWen=0x%0h",this.io_diffCommits_info_214_vlWen,rhs_.io_diffCommits_info_214_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_215_ldest!=rhs_.io_diffCommits_info_215_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_215_ldest=0x%0h while the rhs_.io_diffCommits_info_215_ldest=0x%0h",this.io_diffCommits_info_215_ldest,rhs_.io_diffCommits_info_215_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_215_pdest!=rhs_.io_diffCommits_info_215_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_215_pdest=0x%0h while the rhs_.io_diffCommits_info_215_pdest=0x%0h",this.io_diffCommits_info_215_pdest,rhs_.io_diffCommits_info_215_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_215_rfWen!=rhs_.io_diffCommits_info_215_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_215_rfWen=0x%0h while the rhs_.io_diffCommits_info_215_rfWen=0x%0h",this.io_diffCommits_info_215_rfWen,rhs_.io_diffCommits_info_215_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_215_fpWen!=rhs_.io_diffCommits_info_215_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_215_fpWen=0x%0h while the rhs_.io_diffCommits_info_215_fpWen=0x%0h",this.io_diffCommits_info_215_fpWen,rhs_.io_diffCommits_info_215_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_215_vecWen!=rhs_.io_diffCommits_info_215_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_215_vecWen=0x%0h while the rhs_.io_diffCommits_info_215_vecWen=0x%0h",this.io_diffCommits_info_215_vecWen,rhs_.io_diffCommits_info_215_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_215_v0Wen!=rhs_.io_diffCommits_info_215_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_215_v0Wen=0x%0h while the rhs_.io_diffCommits_info_215_v0Wen=0x%0h",this.io_diffCommits_info_215_v0Wen,rhs_.io_diffCommits_info_215_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_215_vlWen!=rhs_.io_diffCommits_info_215_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_215_vlWen=0x%0h while the rhs_.io_diffCommits_info_215_vlWen=0x%0h",this.io_diffCommits_info_215_vlWen,rhs_.io_diffCommits_info_215_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_216_ldest!=rhs_.io_diffCommits_info_216_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_216_ldest=0x%0h while the rhs_.io_diffCommits_info_216_ldest=0x%0h",this.io_diffCommits_info_216_ldest,rhs_.io_diffCommits_info_216_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_216_pdest!=rhs_.io_diffCommits_info_216_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_216_pdest=0x%0h while the rhs_.io_diffCommits_info_216_pdest=0x%0h",this.io_diffCommits_info_216_pdest,rhs_.io_diffCommits_info_216_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_216_rfWen!=rhs_.io_diffCommits_info_216_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_216_rfWen=0x%0h while the rhs_.io_diffCommits_info_216_rfWen=0x%0h",this.io_diffCommits_info_216_rfWen,rhs_.io_diffCommits_info_216_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_216_fpWen!=rhs_.io_diffCommits_info_216_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_216_fpWen=0x%0h while the rhs_.io_diffCommits_info_216_fpWen=0x%0h",this.io_diffCommits_info_216_fpWen,rhs_.io_diffCommits_info_216_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_216_vecWen!=rhs_.io_diffCommits_info_216_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_216_vecWen=0x%0h while the rhs_.io_diffCommits_info_216_vecWen=0x%0h",this.io_diffCommits_info_216_vecWen,rhs_.io_diffCommits_info_216_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_216_v0Wen!=rhs_.io_diffCommits_info_216_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_216_v0Wen=0x%0h while the rhs_.io_diffCommits_info_216_v0Wen=0x%0h",this.io_diffCommits_info_216_v0Wen,rhs_.io_diffCommits_info_216_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_216_vlWen!=rhs_.io_diffCommits_info_216_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_216_vlWen=0x%0h while the rhs_.io_diffCommits_info_216_vlWen=0x%0h",this.io_diffCommits_info_216_vlWen,rhs_.io_diffCommits_info_216_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_217_ldest!=rhs_.io_diffCommits_info_217_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_217_ldest=0x%0h while the rhs_.io_diffCommits_info_217_ldest=0x%0h",this.io_diffCommits_info_217_ldest,rhs_.io_diffCommits_info_217_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_217_pdest!=rhs_.io_diffCommits_info_217_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_217_pdest=0x%0h while the rhs_.io_diffCommits_info_217_pdest=0x%0h",this.io_diffCommits_info_217_pdest,rhs_.io_diffCommits_info_217_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_217_rfWen!=rhs_.io_diffCommits_info_217_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_217_rfWen=0x%0h while the rhs_.io_diffCommits_info_217_rfWen=0x%0h",this.io_diffCommits_info_217_rfWen,rhs_.io_diffCommits_info_217_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_217_fpWen!=rhs_.io_diffCommits_info_217_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_217_fpWen=0x%0h while the rhs_.io_diffCommits_info_217_fpWen=0x%0h",this.io_diffCommits_info_217_fpWen,rhs_.io_diffCommits_info_217_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_217_vecWen!=rhs_.io_diffCommits_info_217_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_217_vecWen=0x%0h while the rhs_.io_diffCommits_info_217_vecWen=0x%0h",this.io_diffCommits_info_217_vecWen,rhs_.io_diffCommits_info_217_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_217_v0Wen!=rhs_.io_diffCommits_info_217_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_217_v0Wen=0x%0h while the rhs_.io_diffCommits_info_217_v0Wen=0x%0h",this.io_diffCommits_info_217_v0Wen,rhs_.io_diffCommits_info_217_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_217_vlWen!=rhs_.io_diffCommits_info_217_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_217_vlWen=0x%0h while the rhs_.io_diffCommits_info_217_vlWen=0x%0h",this.io_diffCommits_info_217_vlWen,rhs_.io_diffCommits_info_217_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_218_ldest!=rhs_.io_diffCommits_info_218_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_218_ldest=0x%0h while the rhs_.io_diffCommits_info_218_ldest=0x%0h",this.io_diffCommits_info_218_ldest,rhs_.io_diffCommits_info_218_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_218_pdest!=rhs_.io_diffCommits_info_218_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_218_pdest=0x%0h while the rhs_.io_diffCommits_info_218_pdest=0x%0h",this.io_diffCommits_info_218_pdest,rhs_.io_diffCommits_info_218_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_218_rfWen!=rhs_.io_diffCommits_info_218_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_218_rfWen=0x%0h while the rhs_.io_diffCommits_info_218_rfWen=0x%0h",this.io_diffCommits_info_218_rfWen,rhs_.io_diffCommits_info_218_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_218_fpWen!=rhs_.io_diffCommits_info_218_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_218_fpWen=0x%0h while the rhs_.io_diffCommits_info_218_fpWen=0x%0h",this.io_diffCommits_info_218_fpWen,rhs_.io_diffCommits_info_218_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_218_vecWen!=rhs_.io_diffCommits_info_218_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_218_vecWen=0x%0h while the rhs_.io_diffCommits_info_218_vecWen=0x%0h",this.io_diffCommits_info_218_vecWen,rhs_.io_diffCommits_info_218_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_218_v0Wen!=rhs_.io_diffCommits_info_218_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_218_v0Wen=0x%0h while the rhs_.io_diffCommits_info_218_v0Wen=0x%0h",this.io_diffCommits_info_218_v0Wen,rhs_.io_diffCommits_info_218_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_218_vlWen!=rhs_.io_diffCommits_info_218_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_218_vlWen=0x%0h while the rhs_.io_diffCommits_info_218_vlWen=0x%0h",this.io_diffCommits_info_218_vlWen,rhs_.io_diffCommits_info_218_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_219_ldest!=rhs_.io_diffCommits_info_219_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_219_ldest=0x%0h while the rhs_.io_diffCommits_info_219_ldest=0x%0h",this.io_diffCommits_info_219_ldest,rhs_.io_diffCommits_info_219_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_219_pdest!=rhs_.io_diffCommits_info_219_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_219_pdest=0x%0h while the rhs_.io_diffCommits_info_219_pdest=0x%0h",this.io_diffCommits_info_219_pdest,rhs_.io_diffCommits_info_219_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_219_rfWen!=rhs_.io_diffCommits_info_219_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_219_rfWen=0x%0h while the rhs_.io_diffCommits_info_219_rfWen=0x%0h",this.io_diffCommits_info_219_rfWen,rhs_.io_diffCommits_info_219_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_219_fpWen!=rhs_.io_diffCommits_info_219_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_219_fpWen=0x%0h while the rhs_.io_diffCommits_info_219_fpWen=0x%0h",this.io_diffCommits_info_219_fpWen,rhs_.io_diffCommits_info_219_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_219_vecWen!=rhs_.io_diffCommits_info_219_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_219_vecWen=0x%0h while the rhs_.io_diffCommits_info_219_vecWen=0x%0h",this.io_diffCommits_info_219_vecWen,rhs_.io_diffCommits_info_219_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_219_v0Wen!=rhs_.io_diffCommits_info_219_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_219_v0Wen=0x%0h while the rhs_.io_diffCommits_info_219_v0Wen=0x%0h",this.io_diffCommits_info_219_v0Wen,rhs_.io_diffCommits_info_219_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_219_vlWen!=rhs_.io_diffCommits_info_219_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_219_vlWen=0x%0h while the rhs_.io_diffCommits_info_219_vlWen=0x%0h",this.io_diffCommits_info_219_vlWen,rhs_.io_diffCommits_info_219_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_220_ldest!=rhs_.io_diffCommits_info_220_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_220_ldest=0x%0h while the rhs_.io_diffCommits_info_220_ldest=0x%0h",this.io_diffCommits_info_220_ldest,rhs_.io_diffCommits_info_220_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_220_pdest!=rhs_.io_diffCommits_info_220_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_220_pdest=0x%0h while the rhs_.io_diffCommits_info_220_pdest=0x%0h",this.io_diffCommits_info_220_pdest,rhs_.io_diffCommits_info_220_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_220_rfWen!=rhs_.io_diffCommits_info_220_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_220_rfWen=0x%0h while the rhs_.io_diffCommits_info_220_rfWen=0x%0h",this.io_diffCommits_info_220_rfWen,rhs_.io_diffCommits_info_220_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_220_fpWen!=rhs_.io_diffCommits_info_220_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_220_fpWen=0x%0h while the rhs_.io_diffCommits_info_220_fpWen=0x%0h",this.io_diffCommits_info_220_fpWen,rhs_.io_diffCommits_info_220_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_220_vecWen!=rhs_.io_diffCommits_info_220_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_220_vecWen=0x%0h while the rhs_.io_diffCommits_info_220_vecWen=0x%0h",this.io_diffCommits_info_220_vecWen,rhs_.io_diffCommits_info_220_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_220_v0Wen!=rhs_.io_diffCommits_info_220_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_220_v0Wen=0x%0h while the rhs_.io_diffCommits_info_220_v0Wen=0x%0h",this.io_diffCommits_info_220_v0Wen,rhs_.io_diffCommits_info_220_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_220_vlWen!=rhs_.io_diffCommits_info_220_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_220_vlWen=0x%0h while the rhs_.io_diffCommits_info_220_vlWen=0x%0h",this.io_diffCommits_info_220_vlWen,rhs_.io_diffCommits_info_220_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_221_ldest!=rhs_.io_diffCommits_info_221_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_221_ldest=0x%0h while the rhs_.io_diffCommits_info_221_ldest=0x%0h",this.io_diffCommits_info_221_ldest,rhs_.io_diffCommits_info_221_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_221_pdest!=rhs_.io_diffCommits_info_221_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_221_pdest=0x%0h while the rhs_.io_diffCommits_info_221_pdest=0x%0h",this.io_diffCommits_info_221_pdest,rhs_.io_diffCommits_info_221_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_221_rfWen!=rhs_.io_diffCommits_info_221_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_221_rfWen=0x%0h while the rhs_.io_diffCommits_info_221_rfWen=0x%0h",this.io_diffCommits_info_221_rfWen,rhs_.io_diffCommits_info_221_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_221_fpWen!=rhs_.io_diffCommits_info_221_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_221_fpWen=0x%0h while the rhs_.io_diffCommits_info_221_fpWen=0x%0h",this.io_diffCommits_info_221_fpWen,rhs_.io_diffCommits_info_221_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_221_vecWen!=rhs_.io_diffCommits_info_221_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_221_vecWen=0x%0h while the rhs_.io_diffCommits_info_221_vecWen=0x%0h",this.io_diffCommits_info_221_vecWen,rhs_.io_diffCommits_info_221_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_221_v0Wen!=rhs_.io_diffCommits_info_221_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_221_v0Wen=0x%0h while the rhs_.io_diffCommits_info_221_v0Wen=0x%0h",this.io_diffCommits_info_221_v0Wen,rhs_.io_diffCommits_info_221_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_221_vlWen!=rhs_.io_diffCommits_info_221_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_221_vlWen=0x%0h while the rhs_.io_diffCommits_info_221_vlWen=0x%0h",this.io_diffCommits_info_221_vlWen,rhs_.io_diffCommits_info_221_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_222_ldest!=rhs_.io_diffCommits_info_222_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_222_ldest=0x%0h while the rhs_.io_diffCommits_info_222_ldest=0x%0h",this.io_diffCommits_info_222_ldest,rhs_.io_diffCommits_info_222_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_222_pdest!=rhs_.io_diffCommits_info_222_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_222_pdest=0x%0h while the rhs_.io_diffCommits_info_222_pdest=0x%0h",this.io_diffCommits_info_222_pdest,rhs_.io_diffCommits_info_222_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_222_rfWen!=rhs_.io_diffCommits_info_222_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_222_rfWen=0x%0h while the rhs_.io_diffCommits_info_222_rfWen=0x%0h",this.io_diffCommits_info_222_rfWen,rhs_.io_diffCommits_info_222_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_222_fpWen!=rhs_.io_diffCommits_info_222_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_222_fpWen=0x%0h while the rhs_.io_diffCommits_info_222_fpWen=0x%0h",this.io_diffCommits_info_222_fpWen,rhs_.io_diffCommits_info_222_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_222_vecWen!=rhs_.io_diffCommits_info_222_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_222_vecWen=0x%0h while the rhs_.io_diffCommits_info_222_vecWen=0x%0h",this.io_diffCommits_info_222_vecWen,rhs_.io_diffCommits_info_222_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_222_v0Wen!=rhs_.io_diffCommits_info_222_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_222_v0Wen=0x%0h while the rhs_.io_diffCommits_info_222_v0Wen=0x%0h",this.io_diffCommits_info_222_v0Wen,rhs_.io_diffCommits_info_222_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_222_vlWen!=rhs_.io_diffCommits_info_222_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_222_vlWen=0x%0h while the rhs_.io_diffCommits_info_222_vlWen=0x%0h",this.io_diffCommits_info_222_vlWen,rhs_.io_diffCommits_info_222_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_223_ldest!=rhs_.io_diffCommits_info_223_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_223_ldest=0x%0h while the rhs_.io_diffCommits_info_223_ldest=0x%0h",this.io_diffCommits_info_223_ldest,rhs_.io_diffCommits_info_223_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_223_pdest!=rhs_.io_diffCommits_info_223_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_223_pdest=0x%0h while the rhs_.io_diffCommits_info_223_pdest=0x%0h",this.io_diffCommits_info_223_pdest,rhs_.io_diffCommits_info_223_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_223_rfWen!=rhs_.io_diffCommits_info_223_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_223_rfWen=0x%0h while the rhs_.io_diffCommits_info_223_rfWen=0x%0h",this.io_diffCommits_info_223_rfWen,rhs_.io_diffCommits_info_223_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_223_fpWen!=rhs_.io_diffCommits_info_223_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_223_fpWen=0x%0h while the rhs_.io_diffCommits_info_223_fpWen=0x%0h",this.io_diffCommits_info_223_fpWen,rhs_.io_diffCommits_info_223_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_223_vecWen!=rhs_.io_diffCommits_info_223_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_223_vecWen=0x%0h while the rhs_.io_diffCommits_info_223_vecWen=0x%0h",this.io_diffCommits_info_223_vecWen,rhs_.io_diffCommits_info_223_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_223_v0Wen!=rhs_.io_diffCommits_info_223_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_223_v0Wen=0x%0h while the rhs_.io_diffCommits_info_223_v0Wen=0x%0h",this.io_diffCommits_info_223_v0Wen,rhs_.io_diffCommits_info_223_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_223_vlWen!=rhs_.io_diffCommits_info_223_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_223_vlWen=0x%0h while the rhs_.io_diffCommits_info_223_vlWen=0x%0h",this.io_diffCommits_info_223_vlWen,rhs_.io_diffCommits_info_223_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_224_ldest!=rhs_.io_diffCommits_info_224_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_224_ldest=0x%0h while the rhs_.io_diffCommits_info_224_ldest=0x%0h",this.io_diffCommits_info_224_ldest,rhs_.io_diffCommits_info_224_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_224_pdest!=rhs_.io_diffCommits_info_224_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_224_pdest=0x%0h while the rhs_.io_diffCommits_info_224_pdest=0x%0h",this.io_diffCommits_info_224_pdest,rhs_.io_diffCommits_info_224_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_224_rfWen!=rhs_.io_diffCommits_info_224_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_224_rfWen=0x%0h while the rhs_.io_diffCommits_info_224_rfWen=0x%0h",this.io_diffCommits_info_224_rfWen,rhs_.io_diffCommits_info_224_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_224_fpWen!=rhs_.io_diffCommits_info_224_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_224_fpWen=0x%0h while the rhs_.io_diffCommits_info_224_fpWen=0x%0h",this.io_diffCommits_info_224_fpWen,rhs_.io_diffCommits_info_224_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_224_vecWen!=rhs_.io_diffCommits_info_224_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_224_vecWen=0x%0h while the rhs_.io_diffCommits_info_224_vecWen=0x%0h",this.io_diffCommits_info_224_vecWen,rhs_.io_diffCommits_info_224_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_224_v0Wen!=rhs_.io_diffCommits_info_224_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_224_v0Wen=0x%0h while the rhs_.io_diffCommits_info_224_v0Wen=0x%0h",this.io_diffCommits_info_224_v0Wen,rhs_.io_diffCommits_info_224_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_224_vlWen!=rhs_.io_diffCommits_info_224_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_224_vlWen=0x%0h while the rhs_.io_diffCommits_info_224_vlWen=0x%0h",this.io_diffCommits_info_224_vlWen,rhs_.io_diffCommits_info_224_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_225_ldest!=rhs_.io_diffCommits_info_225_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_225_ldest=0x%0h while the rhs_.io_diffCommits_info_225_ldest=0x%0h",this.io_diffCommits_info_225_ldest,rhs_.io_diffCommits_info_225_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_225_pdest!=rhs_.io_diffCommits_info_225_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_225_pdest=0x%0h while the rhs_.io_diffCommits_info_225_pdest=0x%0h",this.io_diffCommits_info_225_pdest,rhs_.io_diffCommits_info_225_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_225_rfWen!=rhs_.io_diffCommits_info_225_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_225_rfWen=0x%0h while the rhs_.io_diffCommits_info_225_rfWen=0x%0h",this.io_diffCommits_info_225_rfWen,rhs_.io_diffCommits_info_225_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_225_fpWen!=rhs_.io_diffCommits_info_225_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_225_fpWen=0x%0h while the rhs_.io_diffCommits_info_225_fpWen=0x%0h",this.io_diffCommits_info_225_fpWen,rhs_.io_diffCommits_info_225_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_225_vecWen!=rhs_.io_diffCommits_info_225_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_225_vecWen=0x%0h while the rhs_.io_diffCommits_info_225_vecWen=0x%0h",this.io_diffCommits_info_225_vecWen,rhs_.io_diffCommits_info_225_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_225_v0Wen!=rhs_.io_diffCommits_info_225_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_225_v0Wen=0x%0h while the rhs_.io_diffCommits_info_225_v0Wen=0x%0h",this.io_diffCommits_info_225_v0Wen,rhs_.io_diffCommits_info_225_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_225_vlWen!=rhs_.io_diffCommits_info_225_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_225_vlWen=0x%0h while the rhs_.io_diffCommits_info_225_vlWen=0x%0h",this.io_diffCommits_info_225_vlWen,rhs_.io_diffCommits_info_225_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_226_ldest!=rhs_.io_diffCommits_info_226_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_226_ldest=0x%0h while the rhs_.io_diffCommits_info_226_ldest=0x%0h",this.io_diffCommits_info_226_ldest,rhs_.io_diffCommits_info_226_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_226_pdest!=rhs_.io_diffCommits_info_226_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_226_pdest=0x%0h while the rhs_.io_diffCommits_info_226_pdest=0x%0h",this.io_diffCommits_info_226_pdest,rhs_.io_diffCommits_info_226_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_226_rfWen!=rhs_.io_diffCommits_info_226_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_226_rfWen=0x%0h while the rhs_.io_diffCommits_info_226_rfWen=0x%0h",this.io_diffCommits_info_226_rfWen,rhs_.io_diffCommits_info_226_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_226_fpWen!=rhs_.io_diffCommits_info_226_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_226_fpWen=0x%0h while the rhs_.io_diffCommits_info_226_fpWen=0x%0h",this.io_diffCommits_info_226_fpWen,rhs_.io_diffCommits_info_226_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_226_vecWen!=rhs_.io_diffCommits_info_226_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_226_vecWen=0x%0h while the rhs_.io_diffCommits_info_226_vecWen=0x%0h",this.io_diffCommits_info_226_vecWen,rhs_.io_diffCommits_info_226_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_226_v0Wen!=rhs_.io_diffCommits_info_226_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_226_v0Wen=0x%0h while the rhs_.io_diffCommits_info_226_v0Wen=0x%0h",this.io_diffCommits_info_226_v0Wen,rhs_.io_diffCommits_info_226_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_226_vlWen!=rhs_.io_diffCommits_info_226_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_226_vlWen=0x%0h while the rhs_.io_diffCommits_info_226_vlWen=0x%0h",this.io_diffCommits_info_226_vlWen,rhs_.io_diffCommits_info_226_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_227_ldest!=rhs_.io_diffCommits_info_227_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_227_ldest=0x%0h while the rhs_.io_diffCommits_info_227_ldest=0x%0h",this.io_diffCommits_info_227_ldest,rhs_.io_diffCommits_info_227_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_227_pdest!=rhs_.io_diffCommits_info_227_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_227_pdest=0x%0h while the rhs_.io_diffCommits_info_227_pdest=0x%0h",this.io_diffCommits_info_227_pdest,rhs_.io_diffCommits_info_227_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_227_rfWen!=rhs_.io_diffCommits_info_227_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_227_rfWen=0x%0h while the rhs_.io_diffCommits_info_227_rfWen=0x%0h",this.io_diffCommits_info_227_rfWen,rhs_.io_diffCommits_info_227_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_227_fpWen!=rhs_.io_diffCommits_info_227_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_227_fpWen=0x%0h while the rhs_.io_diffCommits_info_227_fpWen=0x%0h",this.io_diffCommits_info_227_fpWen,rhs_.io_diffCommits_info_227_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_227_vecWen!=rhs_.io_diffCommits_info_227_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_227_vecWen=0x%0h while the rhs_.io_diffCommits_info_227_vecWen=0x%0h",this.io_diffCommits_info_227_vecWen,rhs_.io_diffCommits_info_227_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_227_v0Wen!=rhs_.io_diffCommits_info_227_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_227_v0Wen=0x%0h while the rhs_.io_diffCommits_info_227_v0Wen=0x%0h",this.io_diffCommits_info_227_v0Wen,rhs_.io_diffCommits_info_227_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_227_vlWen!=rhs_.io_diffCommits_info_227_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_227_vlWen=0x%0h while the rhs_.io_diffCommits_info_227_vlWen=0x%0h",this.io_diffCommits_info_227_vlWen,rhs_.io_diffCommits_info_227_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_228_ldest!=rhs_.io_diffCommits_info_228_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_228_ldest=0x%0h while the rhs_.io_diffCommits_info_228_ldest=0x%0h",this.io_diffCommits_info_228_ldest,rhs_.io_diffCommits_info_228_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_228_pdest!=rhs_.io_diffCommits_info_228_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_228_pdest=0x%0h while the rhs_.io_diffCommits_info_228_pdest=0x%0h",this.io_diffCommits_info_228_pdest,rhs_.io_diffCommits_info_228_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_228_rfWen!=rhs_.io_diffCommits_info_228_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_228_rfWen=0x%0h while the rhs_.io_diffCommits_info_228_rfWen=0x%0h",this.io_diffCommits_info_228_rfWen,rhs_.io_diffCommits_info_228_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_228_fpWen!=rhs_.io_diffCommits_info_228_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_228_fpWen=0x%0h while the rhs_.io_diffCommits_info_228_fpWen=0x%0h",this.io_diffCommits_info_228_fpWen,rhs_.io_diffCommits_info_228_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_228_vecWen!=rhs_.io_diffCommits_info_228_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_228_vecWen=0x%0h while the rhs_.io_diffCommits_info_228_vecWen=0x%0h",this.io_diffCommits_info_228_vecWen,rhs_.io_diffCommits_info_228_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_228_v0Wen!=rhs_.io_diffCommits_info_228_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_228_v0Wen=0x%0h while the rhs_.io_diffCommits_info_228_v0Wen=0x%0h",this.io_diffCommits_info_228_v0Wen,rhs_.io_diffCommits_info_228_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_228_vlWen!=rhs_.io_diffCommits_info_228_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_228_vlWen=0x%0h while the rhs_.io_diffCommits_info_228_vlWen=0x%0h",this.io_diffCommits_info_228_vlWen,rhs_.io_diffCommits_info_228_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_229_ldest!=rhs_.io_diffCommits_info_229_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_229_ldest=0x%0h while the rhs_.io_diffCommits_info_229_ldest=0x%0h",this.io_diffCommits_info_229_ldest,rhs_.io_diffCommits_info_229_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_229_pdest!=rhs_.io_diffCommits_info_229_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_229_pdest=0x%0h while the rhs_.io_diffCommits_info_229_pdest=0x%0h",this.io_diffCommits_info_229_pdest,rhs_.io_diffCommits_info_229_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_229_rfWen!=rhs_.io_diffCommits_info_229_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_229_rfWen=0x%0h while the rhs_.io_diffCommits_info_229_rfWen=0x%0h",this.io_diffCommits_info_229_rfWen,rhs_.io_diffCommits_info_229_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_229_fpWen!=rhs_.io_diffCommits_info_229_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_229_fpWen=0x%0h while the rhs_.io_diffCommits_info_229_fpWen=0x%0h",this.io_diffCommits_info_229_fpWen,rhs_.io_diffCommits_info_229_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_229_vecWen!=rhs_.io_diffCommits_info_229_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_229_vecWen=0x%0h while the rhs_.io_diffCommits_info_229_vecWen=0x%0h",this.io_diffCommits_info_229_vecWen,rhs_.io_diffCommits_info_229_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_229_v0Wen!=rhs_.io_diffCommits_info_229_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_229_v0Wen=0x%0h while the rhs_.io_diffCommits_info_229_v0Wen=0x%0h",this.io_diffCommits_info_229_v0Wen,rhs_.io_diffCommits_info_229_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_229_vlWen!=rhs_.io_diffCommits_info_229_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_229_vlWen=0x%0h while the rhs_.io_diffCommits_info_229_vlWen=0x%0h",this.io_diffCommits_info_229_vlWen,rhs_.io_diffCommits_info_229_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_230_ldest!=rhs_.io_diffCommits_info_230_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_230_ldest=0x%0h while the rhs_.io_diffCommits_info_230_ldest=0x%0h",this.io_diffCommits_info_230_ldest,rhs_.io_diffCommits_info_230_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_230_pdest!=rhs_.io_diffCommits_info_230_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_230_pdest=0x%0h while the rhs_.io_diffCommits_info_230_pdest=0x%0h",this.io_diffCommits_info_230_pdest,rhs_.io_diffCommits_info_230_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_230_rfWen!=rhs_.io_diffCommits_info_230_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_230_rfWen=0x%0h while the rhs_.io_diffCommits_info_230_rfWen=0x%0h",this.io_diffCommits_info_230_rfWen,rhs_.io_diffCommits_info_230_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_230_fpWen!=rhs_.io_diffCommits_info_230_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_230_fpWen=0x%0h while the rhs_.io_diffCommits_info_230_fpWen=0x%0h",this.io_diffCommits_info_230_fpWen,rhs_.io_diffCommits_info_230_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_230_vecWen!=rhs_.io_diffCommits_info_230_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_230_vecWen=0x%0h while the rhs_.io_diffCommits_info_230_vecWen=0x%0h",this.io_diffCommits_info_230_vecWen,rhs_.io_diffCommits_info_230_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_230_v0Wen!=rhs_.io_diffCommits_info_230_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_230_v0Wen=0x%0h while the rhs_.io_diffCommits_info_230_v0Wen=0x%0h",this.io_diffCommits_info_230_v0Wen,rhs_.io_diffCommits_info_230_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_230_vlWen!=rhs_.io_diffCommits_info_230_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_230_vlWen=0x%0h while the rhs_.io_diffCommits_info_230_vlWen=0x%0h",this.io_diffCommits_info_230_vlWen,rhs_.io_diffCommits_info_230_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_231_ldest!=rhs_.io_diffCommits_info_231_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_231_ldest=0x%0h while the rhs_.io_diffCommits_info_231_ldest=0x%0h",this.io_diffCommits_info_231_ldest,rhs_.io_diffCommits_info_231_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_231_pdest!=rhs_.io_diffCommits_info_231_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_231_pdest=0x%0h while the rhs_.io_diffCommits_info_231_pdest=0x%0h",this.io_diffCommits_info_231_pdest,rhs_.io_diffCommits_info_231_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_231_rfWen!=rhs_.io_diffCommits_info_231_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_231_rfWen=0x%0h while the rhs_.io_diffCommits_info_231_rfWen=0x%0h",this.io_diffCommits_info_231_rfWen,rhs_.io_diffCommits_info_231_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_231_fpWen!=rhs_.io_diffCommits_info_231_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_231_fpWen=0x%0h while the rhs_.io_diffCommits_info_231_fpWen=0x%0h",this.io_diffCommits_info_231_fpWen,rhs_.io_diffCommits_info_231_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_231_vecWen!=rhs_.io_diffCommits_info_231_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_231_vecWen=0x%0h while the rhs_.io_diffCommits_info_231_vecWen=0x%0h",this.io_diffCommits_info_231_vecWen,rhs_.io_diffCommits_info_231_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_231_v0Wen!=rhs_.io_diffCommits_info_231_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_231_v0Wen=0x%0h while the rhs_.io_diffCommits_info_231_v0Wen=0x%0h",this.io_diffCommits_info_231_v0Wen,rhs_.io_diffCommits_info_231_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_231_vlWen!=rhs_.io_diffCommits_info_231_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_231_vlWen=0x%0h while the rhs_.io_diffCommits_info_231_vlWen=0x%0h",this.io_diffCommits_info_231_vlWen,rhs_.io_diffCommits_info_231_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_232_ldest!=rhs_.io_diffCommits_info_232_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_232_ldest=0x%0h while the rhs_.io_diffCommits_info_232_ldest=0x%0h",this.io_diffCommits_info_232_ldest,rhs_.io_diffCommits_info_232_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_232_pdest!=rhs_.io_diffCommits_info_232_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_232_pdest=0x%0h while the rhs_.io_diffCommits_info_232_pdest=0x%0h",this.io_diffCommits_info_232_pdest,rhs_.io_diffCommits_info_232_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_232_rfWen!=rhs_.io_diffCommits_info_232_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_232_rfWen=0x%0h while the rhs_.io_diffCommits_info_232_rfWen=0x%0h",this.io_diffCommits_info_232_rfWen,rhs_.io_diffCommits_info_232_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_232_fpWen!=rhs_.io_diffCommits_info_232_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_232_fpWen=0x%0h while the rhs_.io_diffCommits_info_232_fpWen=0x%0h",this.io_diffCommits_info_232_fpWen,rhs_.io_diffCommits_info_232_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_232_vecWen!=rhs_.io_diffCommits_info_232_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_232_vecWen=0x%0h while the rhs_.io_diffCommits_info_232_vecWen=0x%0h",this.io_diffCommits_info_232_vecWen,rhs_.io_diffCommits_info_232_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_232_v0Wen!=rhs_.io_diffCommits_info_232_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_232_v0Wen=0x%0h while the rhs_.io_diffCommits_info_232_v0Wen=0x%0h",this.io_diffCommits_info_232_v0Wen,rhs_.io_diffCommits_info_232_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_232_vlWen!=rhs_.io_diffCommits_info_232_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_232_vlWen=0x%0h while the rhs_.io_diffCommits_info_232_vlWen=0x%0h",this.io_diffCommits_info_232_vlWen,rhs_.io_diffCommits_info_232_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_233_ldest!=rhs_.io_diffCommits_info_233_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_233_ldest=0x%0h while the rhs_.io_diffCommits_info_233_ldest=0x%0h",this.io_diffCommits_info_233_ldest,rhs_.io_diffCommits_info_233_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_233_pdest!=rhs_.io_diffCommits_info_233_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_233_pdest=0x%0h while the rhs_.io_diffCommits_info_233_pdest=0x%0h",this.io_diffCommits_info_233_pdest,rhs_.io_diffCommits_info_233_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_233_rfWen!=rhs_.io_diffCommits_info_233_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_233_rfWen=0x%0h while the rhs_.io_diffCommits_info_233_rfWen=0x%0h",this.io_diffCommits_info_233_rfWen,rhs_.io_diffCommits_info_233_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_233_fpWen!=rhs_.io_diffCommits_info_233_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_233_fpWen=0x%0h while the rhs_.io_diffCommits_info_233_fpWen=0x%0h",this.io_diffCommits_info_233_fpWen,rhs_.io_diffCommits_info_233_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_233_vecWen!=rhs_.io_diffCommits_info_233_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_233_vecWen=0x%0h while the rhs_.io_diffCommits_info_233_vecWen=0x%0h",this.io_diffCommits_info_233_vecWen,rhs_.io_diffCommits_info_233_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_233_v0Wen!=rhs_.io_diffCommits_info_233_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_233_v0Wen=0x%0h while the rhs_.io_diffCommits_info_233_v0Wen=0x%0h",this.io_diffCommits_info_233_v0Wen,rhs_.io_diffCommits_info_233_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_233_vlWen!=rhs_.io_diffCommits_info_233_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_233_vlWen=0x%0h while the rhs_.io_diffCommits_info_233_vlWen=0x%0h",this.io_diffCommits_info_233_vlWen,rhs_.io_diffCommits_info_233_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_234_ldest!=rhs_.io_diffCommits_info_234_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_234_ldest=0x%0h while the rhs_.io_diffCommits_info_234_ldest=0x%0h",this.io_diffCommits_info_234_ldest,rhs_.io_diffCommits_info_234_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_234_pdest!=rhs_.io_diffCommits_info_234_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_234_pdest=0x%0h while the rhs_.io_diffCommits_info_234_pdest=0x%0h",this.io_diffCommits_info_234_pdest,rhs_.io_diffCommits_info_234_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_234_rfWen!=rhs_.io_diffCommits_info_234_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_234_rfWen=0x%0h while the rhs_.io_diffCommits_info_234_rfWen=0x%0h",this.io_diffCommits_info_234_rfWen,rhs_.io_diffCommits_info_234_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_234_fpWen!=rhs_.io_diffCommits_info_234_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_234_fpWen=0x%0h while the rhs_.io_diffCommits_info_234_fpWen=0x%0h",this.io_diffCommits_info_234_fpWen,rhs_.io_diffCommits_info_234_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_234_vecWen!=rhs_.io_diffCommits_info_234_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_234_vecWen=0x%0h while the rhs_.io_diffCommits_info_234_vecWen=0x%0h",this.io_diffCommits_info_234_vecWen,rhs_.io_diffCommits_info_234_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_234_v0Wen!=rhs_.io_diffCommits_info_234_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_234_v0Wen=0x%0h while the rhs_.io_diffCommits_info_234_v0Wen=0x%0h",this.io_diffCommits_info_234_v0Wen,rhs_.io_diffCommits_info_234_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_234_vlWen!=rhs_.io_diffCommits_info_234_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_234_vlWen=0x%0h while the rhs_.io_diffCommits_info_234_vlWen=0x%0h",this.io_diffCommits_info_234_vlWen,rhs_.io_diffCommits_info_234_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_235_ldest!=rhs_.io_diffCommits_info_235_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_235_ldest=0x%0h while the rhs_.io_diffCommits_info_235_ldest=0x%0h",this.io_diffCommits_info_235_ldest,rhs_.io_diffCommits_info_235_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_235_pdest!=rhs_.io_diffCommits_info_235_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_235_pdest=0x%0h while the rhs_.io_diffCommits_info_235_pdest=0x%0h",this.io_diffCommits_info_235_pdest,rhs_.io_diffCommits_info_235_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_235_rfWen!=rhs_.io_diffCommits_info_235_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_235_rfWen=0x%0h while the rhs_.io_diffCommits_info_235_rfWen=0x%0h",this.io_diffCommits_info_235_rfWen,rhs_.io_diffCommits_info_235_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_235_fpWen!=rhs_.io_diffCommits_info_235_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_235_fpWen=0x%0h while the rhs_.io_diffCommits_info_235_fpWen=0x%0h",this.io_diffCommits_info_235_fpWen,rhs_.io_diffCommits_info_235_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_235_vecWen!=rhs_.io_diffCommits_info_235_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_235_vecWen=0x%0h while the rhs_.io_diffCommits_info_235_vecWen=0x%0h",this.io_diffCommits_info_235_vecWen,rhs_.io_diffCommits_info_235_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_235_v0Wen!=rhs_.io_diffCommits_info_235_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_235_v0Wen=0x%0h while the rhs_.io_diffCommits_info_235_v0Wen=0x%0h",this.io_diffCommits_info_235_v0Wen,rhs_.io_diffCommits_info_235_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_235_vlWen!=rhs_.io_diffCommits_info_235_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_235_vlWen=0x%0h while the rhs_.io_diffCommits_info_235_vlWen=0x%0h",this.io_diffCommits_info_235_vlWen,rhs_.io_diffCommits_info_235_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_236_ldest!=rhs_.io_diffCommits_info_236_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_236_ldest=0x%0h while the rhs_.io_diffCommits_info_236_ldest=0x%0h",this.io_diffCommits_info_236_ldest,rhs_.io_diffCommits_info_236_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_236_pdest!=rhs_.io_diffCommits_info_236_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_236_pdest=0x%0h while the rhs_.io_diffCommits_info_236_pdest=0x%0h",this.io_diffCommits_info_236_pdest,rhs_.io_diffCommits_info_236_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_236_rfWen!=rhs_.io_diffCommits_info_236_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_236_rfWen=0x%0h while the rhs_.io_diffCommits_info_236_rfWen=0x%0h",this.io_diffCommits_info_236_rfWen,rhs_.io_diffCommits_info_236_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_236_fpWen!=rhs_.io_diffCommits_info_236_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_236_fpWen=0x%0h while the rhs_.io_diffCommits_info_236_fpWen=0x%0h",this.io_diffCommits_info_236_fpWen,rhs_.io_diffCommits_info_236_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_236_vecWen!=rhs_.io_diffCommits_info_236_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_236_vecWen=0x%0h while the rhs_.io_diffCommits_info_236_vecWen=0x%0h",this.io_diffCommits_info_236_vecWen,rhs_.io_diffCommits_info_236_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_236_v0Wen!=rhs_.io_diffCommits_info_236_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_236_v0Wen=0x%0h while the rhs_.io_diffCommits_info_236_v0Wen=0x%0h",this.io_diffCommits_info_236_v0Wen,rhs_.io_diffCommits_info_236_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_236_vlWen!=rhs_.io_diffCommits_info_236_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_236_vlWen=0x%0h while the rhs_.io_diffCommits_info_236_vlWen=0x%0h",this.io_diffCommits_info_236_vlWen,rhs_.io_diffCommits_info_236_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_237_ldest!=rhs_.io_diffCommits_info_237_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_237_ldest=0x%0h while the rhs_.io_diffCommits_info_237_ldest=0x%0h",this.io_diffCommits_info_237_ldest,rhs_.io_diffCommits_info_237_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_237_pdest!=rhs_.io_diffCommits_info_237_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_237_pdest=0x%0h while the rhs_.io_diffCommits_info_237_pdest=0x%0h",this.io_diffCommits_info_237_pdest,rhs_.io_diffCommits_info_237_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_237_rfWen!=rhs_.io_diffCommits_info_237_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_237_rfWen=0x%0h while the rhs_.io_diffCommits_info_237_rfWen=0x%0h",this.io_diffCommits_info_237_rfWen,rhs_.io_diffCommits_info_237_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_237_fpWen!=rhs_.io_diffCommits_info_237_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_237_fpWen=0x%0h while the rhs_.io_diffCommits_info_237_fpWen=0x%0h",this.io_diffCommits_info_237_fpWen,rhs_.io_diffCommits_info_237_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_237_vecWen!=rhs_.io_diffCommits_info_237_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_237_vecWen=0x%0h while the rhs_.io_diffCommits_info_237_vecWen=0x%0h",this.io_diffCommits_info_237_vecWen,rhs_.io_diffCommits_info_237_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_237_v0Wen!=rhs_.io_diffCommits_info_237_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_237_v0Wen=0x%0h while the rhs_.io_diffCommits_info_237_v0Wen=0x%0h",this.io_diffCommits_info_237_v0Wen,rhs_.io_diffCommits_info_237_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_237_vlWen!=rhs_.io_diffCommits_info_237_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_237_vlWen=0x%0h while the rhs_.io_diffCommits_info_237_vlWen=0x%0h",this.io_diffCommits_info_237_vlWen,rhs_.io_diffCommits_info_237_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_238_ldest!=rhs_.io_diffCommits_info_238_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_238_ldest=0x%0h while the rhs_.io_diffCommits_info_238_ldest=0x%0h",this.io_diffCommits_info_238_ldest,rhs_.io_diffCommits_info_238_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_238_pdest!=rhs_.io_diffCommits_info_238_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_238_pdest=0x%0h while the rhs_.io_diffCommits_info_238_pdest=0x%0h",this.io_diffCommits_info_238_pdest,rhs_.io_diffCommits_info_238_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_238_rfWen!=rhs_.io_diffCommits_info_238_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_238_rfWen=0x%0h while the rhs_.io_diffCommits_info_238_rfWen=0x%0h",this.io_diffCommits_info_238_rfWen,rhs_.io_diffCommits_info_238_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_238_fpWen!=rhs_.io_diffCommits_info_238_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_238_fpWen=0x%0h while the rhs_.io_diffCommits_info_238_fpWen=0x%0h",this.io_diffCommits_info_238_fpWen,rhs_.io_diffCommits_info_238_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_238_vecWen!=rhs_.io_diffCommits_info_238_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_238_vecWen=0x%0h while the rhs_.io_diffCommits_info_238_vecWen=0x%0h",this.io_diffCommits_info_238_vecWen,rhs_.io_diffCommits_info_238_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_238_v0Wen!=rhs_.io_diffCommits_info_238_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_238_v0Wen=0x%0h while the rhs_.io_diffCommits_info_238_v0Wen=0x%0h",this.io_diffCommits_info_238_v0Wen,rhs_.io_diffCommits_info_238_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_238_vlWen!=rhs_.io_diffCommits_info_238_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_238_vlWen=0x%0h while the rhs_.io_diffCommits_info_238_vlWen=0x%0h",this.io_diffCommits_info_238_vlWen,rhs_.io_diffCommits_info_238_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_239_ldest!=rhs_.io_diffCommits_info_239_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_239_ldest=0x%0h while the rhs_.io_diffCommits_info_239_ldest=0x%0h",this.io_diffCommits_info_239_ldest,rhs_.io_diffCommits_info_239_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_239_pdest!=rhs_.io_diffCommits_info_239_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_239_pdest=0x%0h while the rhs_.io_diffCommits_info_239_pdest=0x%0h",this.io_diffCommits_info_239_pdest,rhs_.io_diffCommits_info_239_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_239_rfWen!=rhs_.io_diffCommits_info_239_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_239_rfWen=0x%0h while the rhs_.io_diffCommits_info_239_rfWen=0x%0h",this.io_diffCommits_info_239_rfWen,rhs_.io_diffCommits_info_239_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_239_fpWen!=rhs_.io_diffCommits_info_239_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_239_fpWen=0x%0h while the rhs_.io_diffCommits_info_239_fpWen=0x%0h",this.io_diffCommits_info_239_fpWen,rhs_.io_diffCommits_info_239_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_239_vecWen!=rhs_.io_diffCommits_info_239_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_239_vecWen=0x%0h while the rhs_.io_diffCommits_info_239_vecWen=0x%0h",this.io_diffCommits_info_239_vecWen,rhs_.io_diffCommits_info_239_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_239_v0Wen!=rhs_.io_diffCommits_info_239_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_239_v0Wen=0x%0h while the rhs_.io_diffCommits_info_239_v0Wen=0x%0h",this.io_diffCommits_info_239_v0Wen,rhs_.io_diffCommits_info_239_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_239_vlWen!=rhs_.io_diffCommits_info_239_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_239_vlWen=0x%0h while the rhs_.io_diffCommits_info_239_vlWen=0x%0h",this.io_diffCommits_info_239_vlWen,rhs_.io_diffCommits_info_239_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_240_ldest!=rhs_.io_diffCommits_info_240_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_240_ldest=0x%0h while the rhs_.io_diffCommits_info_240_ldest=0x%0h",this.io_diffCommits_info_240_ldest,rhs_.io_diffCommits_info_240_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_240_pdest!=rhs_.io_diffCommits_info_240_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_240_pdest=0x%0h while the rhs_.io_diffCommits_info_240_pdest=0x%0h",this.io_diffCommits_info_240_pdest,rhs_.io_diffCommits_info_240_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_240_rfWen!=rhs_.io_diffCommits_info_240_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_240_rfWen=0x%0h while the rhs_.io_diffCommits_info_240_rfWen=0x%0h",this.io_diffCommits_info_240_rfWen,rhs_.io_diffCommits_info_240_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_240_fpWen!=rhs_.io_diffCommits_info_240_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_240_fpWen=0x%0h while the rhs_.io_diffCommits_info_240_fpWen=0x%0h",this.io_diffCommits_info_240_fpWen,rhs_.io_diffCommits_info_240_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_240_vecWen!=rhs_.io_diffCommits_info_240_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_240_vecWen=0x%0h while the rhs_.io_diffCommits_info_240_vecWen=0x%0h",this.io_diffCommits_info_240_vecWen,rhs_.io_diffCommits_info_240_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_240_v0Wen!=rhs_.io_diffCommits_info_240_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_240_v0Wen=0x%0h while the rhs_.io_diffCommits_info_240_v0Wen=0x%0h",this.io_diffCommits_info_240_v0Wen,rhs_.io_diffCommits_info_240_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_240_vlWen!=rhs_.io_diffCommits_info_240_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_240_vlWen=0x%0h while the rhs_.io_diffCommits_info_240_vlWen=0x%0h",this.io_diffCommits_info_240_vlWen,rhs_.io_diffCommits_info_240_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_241_ldest!=rhs_.io_diffCommits_info_241_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_241_ldest=0x%0h while the rhs_.io_diffCommits_info_241_ldest=0x%0h",this.io_diffCommits_info_241_ldest,rhs_.io_diffCommits_info_241_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_241_pdest!=rhs_.io_diffCommits_info_241_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_241_pdest=0x%0h while the rhs_.io_diffCommits_info_241_pdest=0x%0h",this.io_diffCommits_info_241_pdest,rhs_.io_diffCommits_info_241_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_241_rfWen!=rhs_.io_diffCommits_info_241_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_241_rfWen=0x%0h while the rhs_.io_diffCommits_info_241_rfWen=0x%0h",this.io_diffCommits_info_241_rfWen,rhs_.io_diffCommits_info_241_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_241_fpWen!=rhs_.io_diffCommits_info_241_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_241_fpWen=0x%0h while the rhs_.io_diffCommits_info_241_fpWen=0x%0h",this.io_diffCommits_info_241_fpWen,rhs_.io_diffCommits_info_241_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_241_vecWen!=rhs_.io_diffCommits_info_241_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_241_vecWen=0x%0h while the rhs_.io_diffCommits_info_241_vecWen=0x%0h",this.io_diffCommits_info_241_vecWen,rhs_.io_diffCommits_info_241_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_241_v0Wen!=rhs_.io_diffCommits_info_241_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_241_v0Wen=0x%0h while the rhs_.io_diffCommits_info_241_v0Wen=0x%0h",this.io_diffCommits_info_241_v0Wen,rhs_.io_diffCommits_info_241_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_241_vlWen!=rhs_.io_diffCommits_info_241_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_241_vlWen=0x%0h while the rhs_.io_diffCommits_info_241_vlWen=0x%0h",this.io_diffCommits_info_241_vlWen,rhs_.io_diffCommits_info_241_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_242_ldest!=rhs_.io_diffCommits_info_242_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_242_ldest=0x%0h while the rhs_.io_diffCommits_info_242_ldest=0x%0h",this.io_diffCommits_info_242_ldest,rhs_.io_diffCommits_info_242_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_242_pdest!=rhs_.io_diffCommits_info_242_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_242_pdest=0x%0h while the rhs_.io_diffCommits_info_242_pdest=0x%0h",this.io_diffCommits_info_242_pdest,rhs_.io_diffCommits_info_242_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_242_rfWen!=rhs_.io_diffCommits_info_242_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_242_rfWen=0x%0h while the rhs_.io_diffCommits_info_242_rfWen=0x%0h",this.io_diffCommits_info_242_rfWen,rhs_.io_diffCommits_info_242_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_242_fpWen!=rhs_.io_diffCommits_info_242_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_242_fpWen=0x%0h while the rhs_.io_diffCommits_info_242_fpWen=0x%0h",this.io_diffCommits_info_242_fpWen,rhs_.io_diffCommits_info_242_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_242_vecWen!=rhs_.io_diffCommits_info_242_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_242_vecWen=0x%0h while the rhs_.io_diffCommits_info_242_vecWen=0x%0h",this.io_diffCommits_info_242_vecWen,rhs_.io_diffCommits_info_242_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_242_v0Wen!=rhs_.io_diffCommits_info_242_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_242_v0Wen=0x%0h while the rhs_.io_diffCommits_info_242_v0Wen=0x%0h",this.io_diffCommits_info_242_v0Wen,rhs_.io_diffCommits_info_242_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_242_vlWen!=rhs_.io_diffCommits_info_242_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_242_vlWen=0x%0h while the rhs_.io_diffCommits_info_242_vlWen=0x%0h",this.io_diffCommits_info_242_vlWen,rhs_.io_diffCommits_info_242_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_243_ldest!=rhs_.io_diffCommits_info_243_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_243_ldest=0x%0h while the rhs_.io_diffCommits_info_243_ldest=0x%0h",this.io_diffCommits_info_243_ldest,rhs_.io_diffCommits_info_243_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_243_pdest!=rhs_.io_diffCommits_info_243_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_243_pdest=0x%0h while the rhs_.io_diffCommits_info_243_pdest=0x%0h",this.io_diffCommits_info_243_pdest,rhs_.io_diffCommits_info_243_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_243_rfWen!=rhs_.io_diffCommits_info_243_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_243_rfWen=0x%0h while the rhs_.io_diffCommits_info_243_rfWen=0x%0h",this.io_diffCommits_info_243_rfWen,rhs_.io_diffCommits_info_243_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_243_fpWen!=rhs_.io_diffCommits_info_243_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_243_fpWen=0x%0h while the rhs_.io_diffCommits_info_243_fpWen=0x%0h",this.io_diffCommits_info_243_fpWen,rhs_.io_diffCommits_info_243_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_243_vecWen!=rhs_.io_diffCommits_info_243_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_243_vecWen=0x%0h while the rhs_.io_diffCommits_info_243_vecWen=0x%0h",this.io_diffCommits_info_243_vecWen,rhs_.io_diffCommits_info_243_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_243_v0Wen!=rhs_.io_diffCommits_info_243_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_243_v0Wen=0x%0h while the rhs_.io_diffCommits_info_243_v0Wen=0x%0h",this.io_diffCommits_info_243_v0Wen,rhs_.io_diffCommits_info_243_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_243_vlWen!=rhs_.io_diffCommits_info_243_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_243_vlWen=0x%0h while the rhs_.io_diffCommits_info_243_vlWen=0x%0h",this.io_diffCommits_info_243_vlWen,rhs_.io_diffCommits_info_243_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_244_ldest!=rhs_.io_diffCommits_info_244_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_244_ldest=0x%0h while the rhs_.io_diffCommits_info_244_ldest=0x%0h",this.io_diffCommits_info_244_ldest,rhs_.io_diffCommits_info_244_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_244_pdest!=rhs_.io_diffCommits_info_244_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_244_pdest=0x%0h while the rhs_.io_diffCommits_info_244_pdest=0x%0h",this.io_diffCommits_info_244_pdest,rhs_.io_diffCommits_info_244_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_244_rfWen!=rhs_.io_diffCommits_info_244_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_244_rfWen=0x%0h while the rhs_.io_diffCommits_info_244_rfWen=0x%0h",this.io_diffCommits_info_244_rfWen,rhs_.io_diffCommits_info_244_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_244_fpWen!=rhs_.io_diffCommits_info_244_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_244_fpWen=0x%0h while the rhs_.io_diffCommits_info_244_fpWen=0x%0h",this.io_diffCommits_info_244_fpWen,rhs_.io_diffCommits_info_244_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_244_vecWen!=rhs_.io_diffCommits_info_244_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_244_vecWen=0x%0h while the rhs_.io_diffCommits_info_244_vecWen=0x%0h",this.io_diffCommits_info_244_vecWen,rhs_.io_diffCommits_info_244_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_244_v0Wen!=rhs_.io_diffCommits_info_244_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_244_v0Wen=0x%0h while the rhs_.io_diffCommits_info_244_v0Wen=0x%0h",this.io_diffCommits_info_244_v0Wen,rhs_.io_diffCommits_info_244_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_244_vlWen!=rhs_.io_diffCommits_info_244_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_244_vlWen=0x%0h while the rhs_.io_diffCommits_info_244_vlWen=0x%0h",this.io_diffCommits_info_244_vlWen,rhs_.io_diffCommits_info_244_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_245_ldest!=rhs_.io_diffCommits_info_245_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_245_ldest=0x%0h while the rhs_.io_diffCommits_info_245_ldest=0x%0h",this.io_diffCommits_info_245_ldest,rhs_.io_diffCommits_info_245_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_245_pdest!=rhs_.io_diffCommits_info_245_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_245_pdest=0x%0h while the rhs_.io_diffCommits_info_245_pdest=0x%0h",this.io_diffCommits_info_245_pdest,rhs_.io_diffCommits_info_245_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_245_rfWen!=rhs_.io_diffCommits_info_245_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_245_rfWen=0x%0h while the rhs_.io_diffCommits_info_245_rfWen=0x%0h",this.io_diffCommits_info_245_rfWen,rhs_.io_diffCommits_info_245_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_245_fpWen!=rhs_.io_diffCommits_info_245_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_245_fpWen=0x%0h while the rhs_.io_diffCommits_info_245_fpWen=0x%0h",this.io_diffCommits_info_245_fpWen,rhs_.io_diffCommits_info_245_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_245_vecWen!=rhs_.io_diffCommits_info_245_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_245_vecWen=0x%0h while the rhs_.io_diffCommits_info_245_vecWen=0x%0h",this.io_diffCommits_info_245_vecWen,rhs_.io_diffCommits_info_245_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_245_v0Wen!=rhs_.io_diffCommits_info_245_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_245_v0Wen=0x%0h while the rhs_.io_diffCommits_info_245_v0Wen=0x%0h",this.io_diffCommits_info_245_v0Wen,rhs_.io_diffCommits_info_245_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_245_vlWen!=rhs_.io_diffCommits_info_245_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_245_vlWen=0x%0h while the rhs_.io_diffCommits_info_245_vlWen=0x%0h",this.io_diffCommits_info_245_vlWen,rhs_.io_diffCommits_info_245_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_246_ldest!=rhs_.io_diffCommits_info_246_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_246_ldest=0x%0h while the rhs_.io_diffCommits_info_246_ldest=0x%0h",this.io_diffCommits_info_246_ldest,rhs_.io_diffCommits_info_246_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_246_pdest!=rhs_.io_diffCommits_info_246_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_246_pdest=0x%0h while the rhs_.io_diffCommits_info_246_pdest=0x%0h",this.io_diffCommits_info_246_pdest,rhs_.io_diffCommits_info_246_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_246_rfWen!=rhs_.io_diffCommits_info_246_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_246_rfWen=0x%0h while the rhs_.io_diffCommits_info_246_rfWen=0x%0h",this.io_diffCommits_info_246_rfWen,rhs_.io_diffCommits_info_246_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_246_fpWen!=rhs_.io_diffCommits_info_246_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_246_fpWen=0x%0h while the rhs_.io_diffCommits_info_246_fpWen=0x%0h",this.io_diffCommits_info_246_fpWen,rhs_.io_diffCommits_info_246_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_246_vecWen!=rhs_.io_diffCommits_info_246_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_246_vecWen=0x%0h while the rhs_.io_diffCommits_info_246_vecWen=0x%0h",this.io_diffCommits_info_246_vecWen,rhs_.io_diffCommits_info_246_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_246_v0Wen!=rhs_.io_diffCommits_info_246_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_246_v0Wen=0x%0h while the rhs_.io_diffCommits_info_246_v0Wen=0x%0h",this.io_diffCommits_info_246_v0Wen,rhs_.io_diffCommits_info_246_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_246_vlWen!=rhs_.io_diffCommits_info_246_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_246_vlWen=0x%0h while the rhs_.io_diffCommits_info_246_vlWen=0x%0h",this.io_diffCommits_info_246_vlWen,rhs_.io_diffCommits_info_246_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_247_ldest!=rhs_.io_diffCommits_info_247_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_247_ldest=0x%0h while the rhs_.io_diffCommits_info_247_ldest=0x%0h",this.io_diffCommits_info_247_ldest,rhs_.io_diffCommits_info_247_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_247_pdest!=rhs_.io_diffCommits_info_247_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_247_pdest=0x%0h while the rhs_.io_diffCommits_info_247_pdest=0x%0h",this.io_diffCommits_info_247_pdest,rhs_.io_diffCommits_info_247_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_247_rfWen!=rhs_.io_diffCommits_info_247_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_247_rfWen=0x%0h while the rhs_.io_diffCommits_info_247_rfWen=0x%0h",this.io_diffCommits_info_247_rfWen,rhs_.io_diffCommits_info_247_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_247_fpWen!=rhs_.io_diffCommits_info_247_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_247_fpWen=0x%0h while the rhs_.io_diffCommits_info_247_fpWen=0x%0h",this.io_diffCommits_info_247_fpWen,rhs_.io_diffCommits_info_247_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_247_vecWen!=rhs_.io_diffCommits_info_247_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_247_vecWen=0x%0h while the rhs_.io_diffCommits_info_247_vecWen=0x%0h",this.io_diffCommits_info_247_vecWen,rhs_.io_diffCommits_info_247_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_247_v0Wen!=rhs_.io_diffCommits_info_247_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_247_v0Wen=0x%0h while the rhs_.io_diffCommits_info_247_v0Wen=0x%0h",this.io_diffCommits_info_247_v0Wen,rhs_.io_diffCommits_info_247_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_247_vlWen!=rhs_.io_diffCommits_info_247_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_247_vlWen=0x%0h while the rhs_.io_diffCommits_info_247_vlWen=0x%0h",this.io_diffCommits_info_247_vlWen,rhs_.io_diffCommits_info_247_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_248_ldest!=rhs_.io_diffCommits_info_248_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_248_ldest=0x%0h while the rhs_.io_diffCommits_info_248_ldest=0x%0h",this.io_diffCommits_info_248_ldest,rhs_.io_diffCommits_info_248_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_248_pdest!=rhs_.io_diffCommits_info_248_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_248_pdest=0x%0h while the rhs_.io_diffCommits_info_248_pdest=0x%0h",this.io_diffCommits_info_248_pdest,rhs_.io_diffCommits_info_248_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_248_rfWen!=rhs_.io_diffCommits_info_248_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_248_rfWen=0x%0h while the rhs_.io_diffCommits_info_248_rfWen=0x%0h",this.io_diffCommits_info_248_rfWen,rhs_.io_diffCommits_info_248_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_248_fpWen!=rhs_.io_diffCommits_info_248_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_248_fpWen=0x%0h while the rhs_.io_diffCommits_info_248_fpWen=0x%0h",this.io_diffCommits_info_248_fpWen,rhs_.io_diffCommits_info_248_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_248_vecWen!=rhs_.io_diffCommits_info_248_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_248_vecWen=0x%0h while the rhs_.io_diffCommits_info_248_vecWen=0x%0h",this.io_diffCommits_info_248_vecWen,rhs_.io_diffCommits_info_248_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_248_v0Wen!=rhs_.io_diffCommits_info_248_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_248_v0Wen=0x%0h while the rhs_.io_diffCommits_info_248_v0Wen=0x%0h",this.io_diffCommits_info_248_v0Wen,rhs_.io_diffCommits_info_248_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_248_vlWen!=rhs_.io_diffCommits_info_248_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_248_vlWen=0x%0h while the rhs_.io_diffCommits_info_248_vlWen=0x%0h",this.io_diffCommits_info_248_vlWen,rhs_.io_diffCommits_info_248_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_249_ldest!=rhs_.io_diffCommits_info_249_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_249_ldest=0x%0h while the rhs_.io_diffCommits_info_249_ldest=0x%0h",this.io_diffCommits_info_249_ldest,rhs_.io_diffCommits_info_249_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_249_pdest!=rhs_.io_diffCommits_info_249_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_249_pdest=0x%0h while the rhs_.io_diffCommits_info_249_pdest=0x%0h",this.io_diffCommits_info_249_pdest,rhs_.io_diffCommits_info_249_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_249_rfWen!=rhs_.io_diffCommits_info_249_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_249_rfWen=0x%0h while the rhs_.io_diffCommits_info_249_rfWen=0x%0h",this.io_diffCommits_info_249_rfWen,rhs_.io_diffCommits_info_249_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_249_fpWen!=rhs_.io_diffCommits_info_249_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_249_fpWen=0x%0h while the rhs_.io_diffCommits_info_249_fpWen=0x%0h",this.io_diffCommits_info_249_fpWen,rhs_.io_diffCommits_info_249_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_249_vecWen!=rhs_.io_diffCommits_info_249_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_249_vecWen=0x%0h while the rhs_.io_diffCommits_info_249_vecWen=0x%0h",this.io_diffCommits_info_249_vecWen,rhs_.io_diffCommits_info_249_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_249_v0Wen!=rhs_.io_diffCommits_info_249_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_249_v0Wen=0x%0h while the rhs_.io_diffCommits_info_249_v0Wen=0x%0h",this.io_diffCommits_info_249_v0Wen,rhs_.io_diffCommits_info_249_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_249_vlWen!=rhs_.io_diffCommits_info_249_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_249_vlWen=0x%0h while the rhs_.io_diffCommits_info_249_vlWen=0x%0h",this.io_diffCommits_info_249_vlWen,rhs_.io_diffCommits_info_249_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_250_ldest!=rhs_.io_diffCommits_info_250_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_250_ldest=0x%0h while the rhs_.io_diffCommits_info_250_ldest=0x%0h",this.io_diffCommits_info_250_ldest,rhs_.io_diffCommits_info_250_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_250_pdest!=rhs_.io_diffCommits_info_250_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_250_pdest=0x%0h while the rhs_.io_diffCommits_info_250_pdest=0x%0h",this.io_diffCommits_info_250_pdest,rhs_.io_diffCommits_info_250_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_250_rfWen!=rhs_.io_diffCommits_info_250_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_250_rfWen=0x%0h while the rhs_.io_diffCommits_info_250_rfWen=0x%0h",this.io_diffCommits_info_250_rfWen,rhs_.io_diffCommits_info_250_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_250_fpWen!=rhs_.io_diffCommits_info_250_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_250_fpWen=0x%0h while the rhs_.io_diffCommits_info_250_fpWen=0x%0h",this.io_diffCommits_info_250_fpWen,rhs_.io_diffCommits_info_250_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_250_vecWen!=rhs_.io_diffCommits_info_250_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_250_vecWen=0x%0h while the rhs_.io_diffCommits_info_250_vecWen=0x%0h",this.io_diffCommits_info_250_vecWen,rhs_.io_diffCommits_info_250_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_250_v0Wen!=rhs_.io_diffCommits_info_250_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_250_v0Wen=0x%0h while the rhs_.io_diffCommits_info_250_v0Wen=0x%0h",this.io_diffCommits_info_250_v0Wen,rhs_.io_diffCommits_info_250_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_250_vlWen!=rhs_.io_diffCommits_info_250_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_250_vlWen=0x%0h while the rhs_.io_diffCommits_info_250_vlWen=0x%0h",this.io_diffCommits_info_250_vlWen,rhs_.io_diffCommits_info_250_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_251_ldest!=rhs_.io_diffCommits_info_251_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_251_ldest=0x%0h while the rhs_.io_diffCommits_info_251_ldest=0x%0h",this.io_diffCommits_info_251_ldest,rhs_.io_diffCommits_info_251_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_251_pdest!=rhs_.io_diffCommits_info_251_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_251_pdest=0x%0h while the rhs_.io_diffCommits_info_251_pdest=0x%0h",this.io_diffCommits_info_251_pdest,rhs_.io_diffCommits_info_251_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_251_rfWen!=rhs_.io_diffCommits_info_251_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_251_rfWen=0x%0h while the rhs_.io_diffCommits_info_251_rfWen=0x%0h",this.io_diffCommits_info_251_rfWen,rhs_.io_diffCommits_info_251_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_251_fpWen!=rhs_.io_diffCommits_info_251_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_251_fpWen=0x%0h while the rhs_.io_diffCommits_info_251_fpWen=0x%0h",this.io_diffCommits_info_251_fpWen,rhs_.io_diffCommits_info_251_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_251_vecWen!=rhs_.io_diffCommits_info_251_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_251_vecWen=0x%0h while the rhs_.io_diffCommits_info_251_vecWen=0x%0h",this.io_diffCommits_info_251_vecWen,rhs_.io_diffCommits_info_251_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_251_v0Wen!=rhs_.io_diffCommits_info_251_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_251_v0Wen=0x%0h while the rhs_.io_diffCommits_info_251_v0Wen=0x%0h",this.io_diffCommits_info_251_v0Wen,rhs_.io_diffCommits_info_251_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_251_vlWen!=rhs_.io_diffCommits_info_251_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_251_vlWen=0x%0h while the rhs_.io_diffCommits_info_251_vlWen=0x%0h",this.io_diffCommits_info_251_vlWen,rhs_.io_diffCommits_info_251_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_252_ldest!=rhs_.io_diffCommits_info_252_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_252_ldest=0x%0h while the rhs_.io_diffCommits_info_252_ldest=0x%0h",this.io_diffCommits_info_252_ldest,rhs_.io_diffCommits_info_252_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_252_pdest!=rhs_.io_diffCommits_info_252_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_252_pdest=0x%0h while the rhs_.io_diffCommits_info_252_pdest=0x%0h",this.io_diffCommits_info_252_pdest,rhs_.io_diffCommits_info_252_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_252_rfWen!=rhs_.io_diffCommits_info_252_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_252_rfWen=0x%0h while the rhs_.io_diffCommits_info_252_rfWen=0x%0h",this.io_diffCommits_info_252_rfWen,rhs_.io_diffCommits_info_252_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_252_fpWen!=rhs_.io_diffCommits_info_252_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_252_fpWen=0x%0h while the rhs_.io_diffCommits_info_252_fpWen=0x%0h",this.io_diffCommits_info_252_fpWen,rhs_.io_diffCommits_info_252_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_252_vecWen!=rhs_.io_diffCommits_info_252_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_252_vecWen=0x%0h while the rhs_.io_diffCommits_info_252_vecWen=0x%0h",this.io_diffCommits_info_252_vecWen,rhs_.io_diffCommits_info_252_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_252_v0Wen!=rhs_.io_diffCommits_info_252_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_252_v0Wen=0x%0h while the rhs_.io_diffCommits_info_252_v0Wen=0x%0h",this.io_diffCommits_info_252_v0Wen,rhs_.io_diffCommits_info_252_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_252_vlWen!=rhs_.io_diffCommits_info_252_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_252_vlWen=0x%0h while the rhs_.io_diffCommits_info_252_vlWen=0x%0h",this.io_diffCommits_info_252_vlWen,rhs_.io_diffCommits_info_252_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_253_ldest!=rhs_.io_diffCommits_info_253_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_253_ldest=0x%0h while the rhs_.io_diffCommits_info_253_ldest=0x%0h",this.io_diffCommits_info_253_ldest,rhs_.io_diffCommits_info_253_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_253_pdest!=rhs_.io_diffCommits_info_253_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_253_pdest=0x%0h while the rhs_.io_diffCommits_info_253_pdest=0x%0h",this.io_diffCommits_info_253_pdest,rhs_.io_diffCommits_info_253_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_253_rfWen!=rhs_.io_diffCommits_info_253_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_253_rfWen=0x%0h while the rhs_.io_diffCommits_info_253_rfWen=0x%0h",this.io_diffCommits_info_253_rfWen,rhs_.io_diffCommits_info_253_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_253_fpWen!=rhs_.io_diffCommits_info_253_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_253_fpWen=0x%0h while the rhs_.io_diffCommits_info_253_fpWen=0x%0h",this.io_diffCommits_info_253_fpWen,rhs_.io_diffCommits_info_253_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_253_vecWen!=rhs_.io_diffCommits_info_253_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_253_vecWen=0x%0h while the rhs_.io_diffCommits_info_253_vecWen=0x%0h",this.io_diffCommits_info_253_vecWen,rhs_.io_diffCommits_info_253_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_253_v0Wen!=rhs_.io_diffCommits_info_253_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_253_v0Wen=0x%0h while the rhs_.io_diffCommits_info_253_v0Wen=0x%0h",this.io_diffCommits_info_253_v0Wen,rhs_.io_diffCommits_info_253_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_253_vlWen!=rhs_.io_diffCommits_info_253_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_253_vlWen=0x%0h while the rhs_.io_diffCommits_info_253_vlWen=0x%0h",this.io_diffCommits_info_253_vlWen,rhs_.io_diffCommits_info_253_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_254_ldest!=rhs_.io_diffCommits_info_254_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_254_ldest=0x%0h while the rhs_.io_diffCommits_info_254_ldest=0x%0h",this.io_diffCommits_info_254_ldest,rhs_.io_diffCommits_info_254_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_254_pdest!=rhs_.io_diffCommits_info_254_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_254_pdest=0x%0h while the rhs_.io_diffCommits_info_254_pdest=0x%0h",this.io_diffCommits_info_254_pdest,rhs_.io_diffCommits_info_254_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_254_rfWen!=rhs_.io_diffCommits_info_254_rfWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_254_rfWen=0x%0h while the rhs_.io_diffCommits_info_254_rfWen=0x%0h",this.io_diffCommits_info_254_rfWen,rhs_.io_diffCommits_info_254_rfWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_254_fpWen!=rhs_.io_diffCommits_info_254_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_254_fpWen=0x%0h while the rhs_.io_diffCommits_info_254_fpWen=0x%0h",this.io_diffCommits_info_254_fpWen,rhs_.io_diffCommits_info_254_fpWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_254_vecWen!=rhs_.io_diffCommits_info_254_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_254_vecWen=0x%0h while the rhs_.io_diffCommits_info_254_vecWen=0x%0h",this.io_diffCommits_info_254_vecWen,rhs_.io_diffCommits_info_254_vecWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_254_v0Wen!=rhs_.io_diffCommits_info_254_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_254_v0Wen=0x%0h while the rhs_.io_diffCommits_info_254_v0Wen=0x%0h",this.io_diffCommits_info_254_v0Wen,rhs_.io_diffCommits_info_254_v0Wen),UVM_NONE)
        end

        if(this.io_diffCommits_info_254_vlWen!=rhs_.io_diffCommits_info_254_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_254_vlWen=0x%0h while the rhs_.io_diffCommits_info_254_vlWen=0x%0h",this.io_diffCommits_info_254_vlWen,rhs_.io_diffCommits_info_254_vlWen),UVM_NONE)
        end

        if(this.io_diffCommits_info_255_ldest!=rhs_.io_diffCommits_info_255_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_255_ldest=0x%0h while the rhs_.io_diffCommits_info_255_ldest=0x%0h",this.io_diffCommits_info_255_ldest,rhs_.io_diffCommits_info_255_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_255_pdest!=rhs_.io_diffCommits_info_255_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_255_pdest=0x%0h while the rhs_.io_diffCommits_info_255_pdest=0x%0h",this.io_diffCommits_info_255_pdest,rhs_.io_diffCommits_info_255_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_256_ldest!=rhs_.io_diffCommits_info_256_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_256_ldest=0x%0h while the rhs_.io_diffCommits_info_256_ldest=0x%0h",this.io_diffCommits_info_256_ldest,rhs_.io_diffCommits_info_256_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_256_pdest!=rhs_.io_diffCommits_info_256_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_256_pdest=0x%0h while the rhs_.io_diffCommits_info_256_pdest=0x%0h",this.io_diffCommits_info_256_pdest,rhs_.io_diffCommits_info_256_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_257_ldest!=rhs_.io_diffCommits_info_257_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_257_ldest=0x%0h while the rhs_.io_diffCommits_info_257_ldest=0x%0h",this.io_diffCommits_info_257_ldest,rhs_.io_diffCommits_info_257_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_257_pdest!=rhs_.io_diffCommits_info_257_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_257_pdest=0x%0h while the rhs_.io_diffCommits_info_257_pdest=0x%0h",this.io_diffCommits_info_257_pdest,rhs_.io_diffCommits_info_257_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_258_ldest!=rhs_.io_diffCommits_info_258_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_258_ldest=0x%0h while the rhs_.io_diffCommits_info_258_ldest=0x%0h",this.io_diffCommits_info_258_ldest,rhs_.io_diffCommits_info_258_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_258_pdest!=rhs_.io_diffCommits_info_258_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_258_pdest=0x%0h while the rhs_.io_diffCommits_info_258_pdest=0x%0h",this.io_diffCommits_info_258_pdest,rhs_.io_diffCommits_info_258_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_259_ldest!=rhs_.io_diffCommits_info_259_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_259_ldest=0x%0h while the rhs_.io_diffCommits_info_259_ldest=0x%0h",this.io_diffCommits_info_259_ldest,rhs_.io_diffCommits_info_259_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_259_pdest!=rhs_.io_diffCommits_info_259_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_259_pdest=0x%0h while the rhs_.io_diffCommits_info_259_pdest=0x%0h",this.io_diffCommits_info_259_pdest,rhs_.io_diffCommits_info_259_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_260_ldest!=rhs_.io_diffCommits_info_260_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_260_ldest=0x%0h while the rhs_.io_diffCommits_info_260_ldest=0x%0h",this.io_diffCommits_info_260_ldest,rhs_.io_diffCommits_info_260_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_260_pdest!=rhs_.io_diffCommits_info_260_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_260_pdest=0x%0h while the rhs_.io_diffCommits_info_260_pdest=0x%0h",this.io_diffCommits_info_260_pdest,rhs_.io_diffCommits_info_260_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_261_ldest!=rhs_.io_diffCommits_info_261_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_261_ldest=0x%0h while the rhs_.io_diffCommits_info_261_ldest=0x%0h",this.io_diffCommits_info_261_ldest,rhs_.io_diffCommits_info_261_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_261_pdest!=rhs_.io_diffCommits_info_261_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_261_pdest=0x%0h while the rhs_.io_diffCommits_info_261_pdest=0x%0h",this.io_diffCommits_info_261_pdest,rhs_.io_diffCommits_info_261_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_262_ldest!=rhs_.io_diffCommits_info_262_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_262_ldest=0x%0h while the rhs_.io_diffCommits_info_262_ldest=0x%0h",this.io_diffCommits_info_262_ldest,rhs_.io_diffCommits_info_262_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_262_pdest!=rhs_.io_diffCommits_info_262_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_262_pdest=0x%0h while the rhs_.io_diffCommits_info_262_pdest=0x%0h",this.io_diffCommits_info_262_pdest,rhs_.io_diffCommits_info_262_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_263_ldest!=rhs_.io_diffCommits_info_263_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_263_ldest=0x%0h while the rhs_.io_diffCommits_info_263_ldest=0x%0h",this.io_diffCommits_info_263_ldest,rhs_.io_diffCommits_info_263_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_263_pdest!=rhs_.io_diffCommits_info_263_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_263_pdest=0x%0h while the rhs_.io_diffCommits_info_263_pdest=0x%0h",this.io_diffCommits_info_263_pdest,rhs_.io_diffCommits_info_263_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_264_ldest!=rhs_.io_diffCommits_info_264_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_264_ldest=0x%0h while the rhs_.io_diffCommits_info_264_ldest=0x%0h",this.io_diffCommits_info_264_ldest,rhs_.io_diffCommits_info_264_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_264_pdest!=rhs_.io_diffCommits_info_264_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_264_pdest=0x%0h while the rhs_.io_diffCommits_info_264_pdest=0x%0h",this.io_diffCommits_info_264_pdest,rhs_.io_diffCommits_info_264_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_265_ldest!=rhs_.io_diffCommits_info_265_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_265_ldest=0x%0h while the rhs_.io_diffCommits_info_265_ldest=0x%0h",this.io_diffCommits_info_265_ldest,rhs_.io_diffCommits_info_265_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_265_pdest!=rhs_.io_diffCommits_info_265_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_265_pdest=0x%0h while the rhs_.io_diffCommits_info_265_pdest=0x%0h",this.io_diffCommits_info_265_pdest,rhs_.io_diffCommits_info_265_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_266_ldest!=rhs_.io_diffCommits_info_266_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_266_ldest=0x%0h while the rhs_.io_diffCommits_info_266_ldest=0x%0h",this.io_diffCommits_info_266_ldest,rhs_.io_diffCommits_info_266_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_266_pdest!=rhs_.io_diffCommits_info_266_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_266_pdest=0x%0h while the rhs_.io_diffCommits_info_266_pdest=0x%0h",this.io_diffCommits_info_266_pdest,rhs_.io_diffCommits_info_266_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_267_ldest!=rhs_.io_diffCommits_info_267_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_267_ldest=0x%0h while the rhs_.io_diffCommits_info_267_ldest=0x%0h",this.io_diffCommits_info_267_ldest,rhs_.io_diffCommits_info_267_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_267_pdest!=rhs_.io_diffCommits_info_267_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_267_pdest=0x%0h while the rhs_.io_diffCommits_info_267_pdest=0x%0h",this.io_diffCommits_info_267_pdest,rhs_.io_diffCommits_info_267_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_268_ldest!=rhs_.io_diffCommits_info_268_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_268_ldest=0x%0h while the rhs_.io_diffCommits_info_268_ldest=0x%0h",this.io_diffCommits_info_268_ldest,rhs_.io_diffCommits_info_268_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_268_pdest!=rhs_.io_diffCommits_info_268_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_268_pdest=0x%0h while the rhs_.io_diffCommits_info_268_pdest=0x%0h",this.io_diffCommits_info_268_pdest,rhs_.io_diffCommits_info_268_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_269_ldest!=rhs_.io_diffCommits_info_269_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_269_ldest=0x%0h while the rhs_.io_diffCommits_info_269_ldest=0x%0h",this.io_diffCommits_info_269_ldest,rhs_.io_diffCommits_info_269_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_269_pdest!=rhs_.io_diffCommits_info_269_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_269_pdest=0x%0h while the rhs_.io_diffCommits_info_269_pdest=0x%0h",this.io_diffCommits_info_269_pdest,rhs_.io_diffCommits_info_269_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_270_ldest!=rhs_.io_diffCommits_info_270_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_270_ldest=0x%0h while the rhs_.io_diffCommits_info_270_ldest=0x%0h",this.io_diffCommits_info_270_ldest,rhs_.io_diffCommits_info_270_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_270_pdest!=rhs_.io_diffCommits_info_270_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_270_pdest=0x%0h while the rhs_.io_diffCommits_info_270_pdest=0x%0h",this.io_diffCommits_info_270_pdest,rhs_.io_diffCommits_info_270_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_271_ldest!=rhs_.io_diffCommits_info_271_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_271_ldest=0x%0h while the rhs_.io_diffCommits_info_271_ldest=0x%0h",this.io_diffCommits_info_271_ldest,rhs_.io_diffCommits_info_271_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_271_pdest!=rhs_.io_diffCommits_info_271_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_271_pdest=0x%0h while the rhs_.io_diffCommits_info_271_pdest=0x%0h",this.io_diffCommits_info_271_pdest,rhs_.io_diffCommits_info_271_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_272_ldest!=rhs_.io_diffCommits_info_272_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_272_ldest=0x%0h while the rhs_.io_diffCommits_info_272_ldest=0x%0h",this.io_diffCommits_info_272_ldest,rhs_.io_diffCommits_info_272_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_272_pdest!=rhs_.io_diffCommits_info_272_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_272_pdest=0x%0h while the rhs_.io_diffCommits_info_272_pdest=0x%0h",this.io_diffCommits_info_272_pdest,rhs_.io_diffCommits_info_272_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_273_ldest!=rhs_.io_diffCommits_info_273_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_273_ldest=0x%0h while the rhs_.io_diffCommits_info_273_ldest=0x%0h",this.io_diffCommits_info_273_ldest,rhs_.io_diffCommits_info_273_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_273_pdest!=rhs_.io_diffCommits_info_273_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_273_pdest=0x%0h while the rhs_.io_diffCommits_info_273_pdest=0x%0h",this.io_diffCommits_info_273_pdest,rhs_.io_diffCommits_info_273_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_274_ldest!=rhs_.io_diffCommits_info_274_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_274_ldest=0x%0h while the rhs_.io_diffCommits_info_274_ldest=0x%0h",this.io_diffCommits_info_274_ldest,rhs_.io_diffCommits_info_274_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_274_pdest!=rhs_.io_diffCommits_info_274_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_274_pdest=0x%0h while the rhs_.io_diffCommits_info_274_pdest=0x%0h",this.io_diffCommits_info_274_pdest,rhs_.io_diffCommits_info_274_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_275_ldest!=rhs_.io_diffCommits_info_275_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_275_ldest=0x%0h while the rhs_.io_diffCommits_info_275_ldest=0x%0h",this.io_diffCommits_info_275_ldest,rhs_.io_diffCommits_info_275_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_275_pdest!=rhs_.io_diffCommits_info_275_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_275_pdest=0x%0h while the rhs_.io_diffCommits_info_275_pdest=0x%0h",this.io_diffCommits_info_275_pdest,rhs_.io_diffCommits_info_275_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_276_ldest!=rhs_.io_diffCommits_info_276_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_276_ldest=0x%0h while the rhs_.io_diffCommits_info_276_ldest=0x%0h",this.io_diffCommits_info_276_ldest,rhs_.io_diffCommits_info_276_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_276_pdest!=rhs_.io_diffCommits_info_276_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_276_pdest=0x%0h while the rhs_.io_diffCommits_info_276_pdest=0x%0h",this.io_diffCommits_info_276_pdest,rhs_.io_diffCommits_info_276_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_277_ldest!=rhs_.io_diffCommits_info_277_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_277_ldest=0x%0h while the rhs_.io_diffCommits_info_277_ldest=0x%0h",this.io_diffCommits_info_277_ldest,rhs_.io_diffCommits_info_277_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_277_pdest!=rhs_.io_diffCommits_info_277_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_277_pdest=0x%0h while the rhs_.io_diffCommits_info_277_pdest=0x%0h",this.io_diffCommits_info_277_pdest,rhs_.io_diffCommits_info_277_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_278_ldest!=rhs_.io_diffCommits_info_278_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_278_ldest=0x%0h while the rhs_.io_diffCommits_info_278_ldest=0x%0h",this.io_diffCommits_info_278_ldest,rhs_.io_diffCommits_info_278_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_278_pdest!=rhs_.io_diffCommits_info_278_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_278_pdest=0x%0h while the rhs_.io_diffCommits_info_278_pdest=0x%0h",this.io_diffCommits_info_278_pdest,rhs_.io_diffCommits_info_278_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_279_ldest!=rhs_.io_diffCommits_info_279_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_279_ldest=0x%0h while the rhs_.io_diffCommits_info_279_ldest=0x%0h",this.io_diffCommits_info_279_ldest,rhs_.io_diffCommits_info_279_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_279_pdest!=rhs_.io_diffCommits_info_279_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_279_pdest=0x%0h while the rhs_.io_diffCommits_info_279_pdest=0x%0h",this.io_diffCommits_info_279_pdest,rhs_.io_diffCommits_info_279_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_280_ldest!=rhs_.io_diffCommits_info_280_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_280_ldest=0x%0h while the rhs_.io_diffCommits_info_280_ldest=0x%0h",this.io_diffCommits_info_280_ldest,rhs_.io_diffCommits_info_280_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_280_pdest!=rhs_.io_diffCommits_info_280_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_280_pdest=0x%0h while the rhs_.io_diffCommits_info_280_pdest=0x%0h",this.io_diffCommits_info_280_pdest,rhs_.io_diffCommits_info_280_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_281_ldest!=rhs_.io_diffCommits_info_281_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_281_ldest=0x%0h while the rhs_.io_diffCommits_info_281_ldest=0x%0h",this.io_diffCommits_info_281_ldest,rhs_.io_diffCommits_info_281_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_281_pdest!=rhs_.io_diffCommits_info_281_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_281_pdest=0x%0h while the rhs_.io_diffCommits_info_281_pdest=0x%0h",this.io_diffCommits_info_281_pdest,rhs_.io_diffCommits_info_281_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_282_ldest!=rhs_.io_diffCommits_info_282_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_282_ldest=0x%0h while the rhs_.io_diffCommits_info_282_ldest=0x%0h",this.io_diffCommits_info_282_ldest,rhs_.io_diffCommits_info_282_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_282_pdest!=rhs_.io_diffCommits_info_282_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_282_pdest=0x%0h while the rhs_.io_diffCommits_info_282_pdest=0x%0h",this.io_diffCommits_info_282_pdest,rhs_.io_diffCommits_info_282_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_283_ldest!=rhs_.io_diffCommits_info_283_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_283_ldest=0x%0h while the rhs_.io_diffCommits_info_283_ldest=0x%0h",this.io_diffCommits_info_283_ldest,rhs_.io_diffCommits_info_283_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_283_pdest!=rhs_.io_diffCommits_info_283_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_283_pdest=0x%0h while the rhs_.io_diffCommits_info_283_pdest=0x%0h",this.io_diffCommits_info_283_pdest,rhs_.io_diffCommits_info_283_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_284_ldest!=rhs_.io_diffCommits_info_284_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_284_ldest=0x%0h while the rhs_.io_diffCommits_info_284_ldest=0x%0h",this.io_diffCommits_info_284_ldest,rhs_.io_diffCommits_info_284_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_284_pdest!=rhs_.io_diffCommits_info_284_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_284_pdest=0x%0h while the rhs_.io_diffCommits_info_284_pdest=0x%0h",this.io_diffCommits_info_284_pdest,rhs_.io_diffCommits_info_284_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_285_ldest!=rhs_.io_diffCommits_info_285_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_285_ldest=0x%0h while the rhs_.io_diffCommits_info_285_ldest=0x%0h",this.io_diffCommits_info_285_ldest,rhs_.io_diffCommits_info_285_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_285_pdest!=rhs_.io_diffCommits_info_285_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_285_pdest=0x%0h while the rhs_.io_diffCommits_info_285_pdest=0x%0h",this.io_diffCommits_info_285_pdest,rhs_.io_diffCommits_info_285_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_286_ldest!=rhs_.io_diffCommits_info_286_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_286_ldest=0x%0h while the rhs_.io_diffCommits_info_286_ldest=0x%0h",this.io_diffCommits_info_286_ldest,rhs_.io_diffCommits_info_286_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_286_pdest!=rhs_.io_diffCommits_info_286_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_286_pdest=0x%0h while the rhs_.io_diffCommits_info_286_pdest=0x%0h",this.io_diffCommits_info_286_pdest,rhs_.io_diffCommits_info_286_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_287_ldest!=rhs_.io_diffCommits_info_287_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_287_ldest=0x%0h while the rhs_.io_diffCommits_info_287_ldest=0x%0h",this.io_diffCommits_info_287_ldest,rhs_.io_diffCommits_info_287_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_287_pdest!=rhs_.io_diffCommits_info_287_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_287_pdest=0x%0h while the rhs_.io_diffCommits_info_287_pdest=0x%0h",this.io_diffCommits_info_287_pdest,rhs_.io_diffCommits_info_287_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_288_ldest!=rhs_.io_diffCommits_info_288_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_288_ldest=0x%0h while the rhs_.io_diffCommits_info_288_ldest=0x%0h",this.io_diffCommits_info_288_ldest,rhs_.io_diffCommits_info_288_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_288_pdest!=rhs_.io_diffCommits_info_288_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_288_pdest=0x%0h while the rhs_.io_diffCommits_info_288_pdest=0x%0h",this.io_diffCommits_info_288_pdest,rhs_.io_diffCommits_info_288_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_289_ldest!=rhs_.io_diffCommits_info_289_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_289_ldest=0x%0h while the rhs_.io_diffCommits_info_289_ldest=0x%0h",this.io_diffCommits_info_289_ldest,rhs_.io_diffCommits_info_289_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_289_pdest!=rhs_.io_diffCommits_info_289_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_289_pdest=0x%0h while the rhs_.io_diffCommits_info_289_pdest=0x%0h",this.io_diffCommits_info_289_pdest,rhs_.io_diffCommits_info_289_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_290_ldest!=rhs_.io_diffCommits_info_290_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_290_ldest=0x%0h while the rhs_.io_diffCommits_info_290_ldest=0x%0h",this.io_diffCommits_info_290_ldest,rhs_.io_diffCommits_info_290_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_290_pdest!=rhs_.io_diffCommits_info_290_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_290_pdest=0x%0h while the rhs_.io_diffCommits_info_290_pdest=0x%0h",this.io_diffCommits_info_290_pdest,rhs_.io_diffCommits_info_290_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_291_ldest!=rhs_.io_diffCommits_info_291_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_291_ldest=0x%0h while the rhs_.io_diffCommits_info_291_ldest=0x%0h",this.io_diffCommits_info_291_ldest,rhs_.io_diffCommits_info_291_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_291_pdest!=rhs_.io_diffCommits_info_291_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_291_pdest=0x%0h while the rhs_.io_diffCommits_info_291_pdest=0x%0h",this.io_diffCommits_info_291_pdest,rhs_.io_diffCommits_info_291_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_292_ldest!=rhs_.io_diffCommits_info_292_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_292_ldest=0x%0h while the rhs_.io_diffCommits_info_292_ldest=0x%0h",this.io_diffCommits_info_292_ldest,rhs_.io_diffCommits_info_292_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_292_pdest!=rhs_.io_diffCommits_info_292_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_292_pdest=0x%0h while the rhs_.io_diffCommits_info_292_pdest=0x%0h",this.io_diffCommits_info_292_pdest,rhs_.io_diffCommits_info_292_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_293_ldest!=rhs_.io_diffCommits_info_293_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_293_ldest=0x%0h while the rhs_.io_diffCommits_info_293_ldest=0x%0h",this.io_diffCommits_info_293_ldest,rhs_.io_diffCommits_info_293_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_293_pdest!=rhs_.io_diffCommits_info_293_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_293_pdest=0x%0h while the rhs_.io_diffCommits_info_293_pdest=0x%0h",this.io_diffCommits_info_293_pdest,rhs_.io_diffCommits_info_293_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_294_ldest!=rhs_.io_diffCommits_info_294_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_294_ldest=0x%0h while the rhs_.io_diffCommits_info_294_ldest=0x%0h",this.io_diffCommits_info_294_ldest,rhs_.io_diffCommits_info_294_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_294_pdest!=rhs_.io_diffCommits_info_294_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_294_pdest=0x%0h while the rhs_.io_diffCommits_info_294_pdest=0x%0h",this.io_diffCommits_info_294_pdest,rhs_.io_diffCommits_info_294_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_295_ldest!=rhs_.io_diffCommits_info_295_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_295_ldest=0x%0h while the rhs_.io_diffCommits_info_295_ldest=0x%0h",this.io_diffCommits_info_295_ldest,rhs_.io_diffCommits_info_295_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_295_pdest!=rhs_.io_diffCommits_info_295_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_295_pdest=0x%0h while the rhs_.io_diffCommits_info_295_pdest=0x%0h",this.io_diffCommits_info_295_pdest,rhs_.io_diffCommits_info_295_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_296_ldest!=rhs_.io_diffCommits_info_296_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_296_ldest=0x%0h while the rhs_.io_diffCommits_info_296_ldest=0x%0h",this.io_diffCommits_info_296_ldest,rhs_.io_diffCommits_info_296_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_296_pdest!=rhs_.io_diffCommits_info_296_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_296_pdest=0x%0h while the rhs_.io_diffCommits_info_296_pdest=0x%0h",this.io_diffCommits_info_296_pdest,rhs_.io_diffCommits_info_296_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_297_ldest!=rhs_.io_diffCommits_info_297_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_297_ldest=0x%0h while the rhs_.io_diffCommits_info_297_ldest=0x%0h",this.io_diffCommits_info_297_ldest,rhs_.io_diffCommits_info_297_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_297_pdest!=rhs_.io_diffCommits_info_297_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_297_pdest=0x%0h while the rhs_.io_diffCommits_info_297_pdest=0x%0h",this.io_diffCommits_info_297_pdest,rhs_.io_diffCommits_info_297_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_298_ldest!=rhs_.io_diffCommits_info_298_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_298_ldest=0x%0h while the rhs_.io_diffCommits_info_298_ldest=0x%0h",this.io_diffCommits_info_298_ldest,rhs_.io_diffCommits_info_298_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_298_pdest!=rhs_.io_diffCommits_info_298_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_298_pdest=0x%0h while the rhs_.io_diffCommits_info_298_pdest=0x%0h",this.io_diffCommits_info_298_pdest,rhs_.io_diffCommits_info_298_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_299_ldest!=rhs_.io_diffCommits_info_299_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_299_ldest=0x%0h while the rhs_.io_diffCommits_info_299_ldest=0x%0h",this.io_diffCommits_info_299_ldest,rhs_.io_diffCommits_info_299_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_299_pdest!=rhs_.io_diffCommits_info_299_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_299_pdest=0x%0h while the rhs_.io_diffCommits_info_299_pdest=0x%0h",this.io_diffCommits_info_299_pdest,rhs_.io_diffCommits_info_299_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_300_ldest!=rhs_.io_diffCommits_info_300_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_300_ldest=0x%0h while the rhs_.io_diffCommits_info_300_ldest=0x%0h",this.io_diffCommits_info_300_ldest,rhs_.io_diffCommits_info_300_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_300_pdest!=rhs_.io_diffCommits_info_300_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_300_pdest=0x%0h while the rhs_.io_diffCommits_info_300_pdest=0x%0h",this.io_diffCommits_info_300_pdest,rhs_.io_diffCommits_info_300_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_301_ldest!=rhs_.io_diffCommits_info_301_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_301_ldest=0x%0h while the rhs_.io_diffCommits_info_301_ldest=0x%0h",this.io_diffCommits_info_301_ldest,rhs_.io_diffCommits_info_301_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_301_pdest!=rhs_.io_diffCommits_info_301_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_301_pdest=0x%0h while the rhs_.io_diffCommits_info_301_pdest=0x%0h",this.io_diffCommits_info_301_pdest,rhs_.io_diffCommits_info_301_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_302_ldest!=rhs_.io_diffCommits_info_302_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_302_ldest=0x%0h while the rhs_.io_diffCommits_info_302_ldest=0x%0h",this.io_diffCommits_info_302_ldest,rhs_.io_diffCommits_info_302_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_302_pdest!=rhs_.io_diffCommits_info_302_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_302_pdest=0x%0h while the rhs_.io_diffCommits_info_302_pdest=0x%0h",this.io_diffCommits_info_302_pdest,rhs_.io_diffCommits_info_302_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_303_ldest!=rhs_.io_diffCommits_info_303_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_303_ldest=0x%0h while the rhs_.io_diffCommits_info_303_ldest=0x%0h",this.io_diffCommits_info_303_ldest,rhs_.io_diffCommits_info_303_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_303_pdest!=rhs_.io_diffCommits_info_303_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_303_pdest=0x%0h while the rhs_.io_diffCommits_info_303_pdest=0x%0h",this.io_diffCommits_info_303_pdest,rhs_.io_diffCommits_info_303_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_304_ldest!=rhs_.io_diffCommits_info_304_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_304_ldest=0x%0h while the rhs_.io_diffCommits_info_304_ldest=0x%0h",this.io_diffCommits_info_304_ldest,rhs_.io_diffCommits_info_304_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_304_pdest!=rhs_.io_diffCommits_info_304_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_304_pdest=0x%0h while the rhs_.io_diffCommits_info_304_pdest=0x%0h",this.io_diffCommits_info_304_pdest,rhs_.io_diffCommits_info_304_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_305_ldest!=rhs_.io_diffCommits_info_305_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_305_ldest=0x%0h while the rhs_.io_diffCommits_info_305_ldest=0x%0h",this.io_diffCommits_info_305_ldest,rhs_.io_diffCommits_info_305_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_305_pdest!=rhs_.io_diffCommits_info_305_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_305_pdest=0x%0h while the rhs_.io_diffCommits_info_305_pdest=0x%0h",this.io_diffCommits_info_305_pdest,rhs_.io_diffCommits_info_305_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_306_ldest!=rhs_.io_diffCommits_info_306_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_306_ldest=0x%0h while the rhs_.io_diffCommits_info_306_ldest=0x%0h",this.io_diffCommits_info_306_ldest,rhs_.io_diffCommits_info_306_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_306_pdest!=rhs_.io_diffCommits_info_306_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_306_pdest=0x%0h while the rhs_.io_diffCommits_info_306_pdest=0x%0h",this.io_diffCommits_info_306_pdest,rhs_.io_diffCommits_info_306_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_307_ldest!=rhs_.io_diffCommits_info_307_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_307_ldest=0x%0h while the rhs_.io_diffCommits_info_307_ldest=0x%0h",this.io_diffCommits_info_307_ldest,rhs_.io_diffCommits_info_307_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_307_pdest!=rhs_.io_diffCommits_info_307_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_307_pdest=0x%0h while the rhs_.io_diffCommits_info_307_pdest=0x%0h",this.io_diffCommits_info_307_pdest,rhs_.io_diffCommits_info_307_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_308_ldest!=rhs_.io_diffCommits_info_308_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_308_ldest=0x%0h while the rhs_.io_diffCommits_info_308_ldest=0x%0h",this.io_diffCommits_info_308_ldest,rhs_.io_diffCommits_info_308_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_308_pdest!=rhs_.io_diffCommits_info_308_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_308_pdest=0x%0h while the rhs_.io_diffCommits_info_308_pdest=0x%0h",this.io_diffCommits_info_308_pdest,rhs_.io_diffCommits_info_308_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_309_ldest!=rhs_.io_diffCommits_info_309_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_309_ldest=0x%0h while the rhs_.io_diffCommits_info_309_ldest=0x%0h",this.io_diffCommits_info_309_ldest,rhs_.io_diffCommits_info_309_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_309_pdest!=rhs_.io_diffCommits_info_309_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_309_pdest=0x%0h while the rhs_.io_diffCommits_info_309_pdest=0x%0h",this.io_diffCommits_info_309_pdest,rhs_.io_diffCommits_info_309_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_310_ldest!=rhs_.io_diffCommits_info_310_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_310_ldest=0x%0h while the rhs_.io_diffCommits_info_310_ldest=0x%0h",this.io_diffCommits_info_310_ldest,rhs_.io_diffCommits_info_310_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_310_pdest!=rhs_.io_diffCommits_info_310_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_310_pdest=0x%0h while the rhs_.io_diffCommits_info_310_pdest=0x%0h",this.io_diffCommits_info_310_pdest,rhs_.io_diffCommits_info_310_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_311_ldest!=rhs_.io_diffCommits_info_311_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_311_ldest=0x%0h while the rhs_.io_diffCommits_info_311_ldest=0x%0h",this.io_diffCommits_info_311_ldest,rhs_.io_diffCommits_info_311_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_311_pdest!=rhs_.io_diffCommits_info_311_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_311_pdest=0x%0h while the rhs_.io_diffCommits_info_311_pdest=0x%0h",this.io_diffCommits_info_311_pdest,rhs_.io_diffCommits_info_311_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_312_ldest!=rhs_.io_diffCommits_info_312_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_312_ldest=0x%0h while the rhs_.io_diffCommits_info_312_ldest=0x%0h",this.io_diffCommits_info_312_ldest,rhs_.io_diffCommits_info_312_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_312_pdest!=rhs_.io_diffCommits_info_312_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_312_pdest=0x%0h while the rhs_.io_diffCommits_info_312_pdest=0x%0h",this.io_diffCommits_info_312_pdest,rhs_.io_diffCommits_info_312_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_313_ldest!=rhs_.io_diffCommits_info_313_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_313_ldest=0x%0h while the rhs_.io_diffCommits_info_313_ldest=0x%0h",this.io_diffCommits_info_313_ldest,rhs_.io_diffCommits_info_313_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_313_pdest!=rhs_.io_diffCommits_info_313_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_313_pdest=0x%0h while the rhs_.io_diffCommits_info_313_pdest=0x%0h",this.io_diffCommits_info_313_pdest,rhs_.io_diffCommits_info_313_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_314_ldest!=rhs_.io_diffCommits_info_314_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_314_ldest=0x%0h while the rhs_.io_diffCommits_info_314_ldest=0x%0h",this.io_diffCommits_info_314_ldest,rhs_.io_diffCommits_info_314_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_314_pdest!=rhs_.io_diffCommits_info_314_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_314_pdest=0x%0h while the rhs_.io_diffCommits_info_314_pdest=0x%0h",this.io_diffCommits_info_314_pdest,rhs_.io_diffCommits_info_314_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_315_ldest!=rhs_.io_diffCommits_info_315_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_315_ldest=0x%0h while the rhs_.io_diffCommits_info_315_ldest=0x%0h",this.io_diffCommits_info_315_ldest,rhs_.io_diffCommits_info_315_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_315_pdest!=rhs_.io_diffCommits_info_315_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_315_pdest=0x%0h while the rhs_.io_diffCommits_info_315_pdest=0x%0h",this.io_diffCommits_info_315_pdest,rhs_.io_diffCommits_info_315_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_316_ldest!=rhs_.io_diffCommits_info_316_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_316_ldest=0x%0h while the rhs_.io_diffCommits_info_316_ldest=0x%0h",this.io_diffCommits_info_316_ldest,rhs_.io_diffCommits_info_316_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_316_pdest!=rhs_.io_diffCommits_info_316_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_316_pdest=0x%0h while the rhs_.io_diffCommits_info_316_pdest=0x%0h",this.io_diffCommits_info_316_pdest,rhs_.io_diffCommits_info_316_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_317_ldest!=rhs_.io_diffCommits_info_317_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_317_ldest=0x%0h while the rhs_.io_diffCommits_info_317_ldest=0x%0h",this.io_diffCommits_info_317_ldest,rhs_.io_diffCommits_info_317_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_317_pdest!=rhs_.io_diffCommits_info_317_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_317_pdest=0x%0h while the rhs_.io_diffCommits_info_317_pdest=0x%0h",this.io_diffCommits_info_317_pdest,rhs_.io_diffCommits_info_317_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_318_ldest!=rhs_.io_diffCommits_info_318_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_318_ldest=0x%0h while the rhs_.io_diffCommits_info_318_ldest=0x%0h",this.io_diffCommits_info_318_ldest,rhs_.io_diffCommits_info_318_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_318_pdest!=rhs_.io_diffCommits_info_318_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_318_pdest=0x%0h while the rhs_.io_diffCommits_info_318_pdest=0x%0h",this.io_diffCommits_info_318_pdest,rhs_.io_diffCommits_info_318_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_319_ldest!=rhs_.io_diffCommits_info_319_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_319_ldest=0x%0h while the rhs_.io_diffCommits_info_319_ldest=0x%0h",this.io_diffCommits_info_319_ldest,rhs_.io_diffCommits_info_319_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_319_pdest!=rhs_.io_diffCommits_info_319_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_319_pdest=0x%0h while the rhs_.io_diffCommits_info_319_pdest=0x%0h",this.io_diffCommits_info_319_pdest,rhs_.io_diffCommits_info_319_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_320_ldest!=rhs_.io_diffCommits_info_320_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_320_ldest=0x%0h while the rhs_.io_diffCommits_info_320_ldest=0x%0h",this.io_diffCommits_info_320_ldest,rhs_.io_diffCommits_info_320_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_320_pdest!=rhs_.io_diffCommits_info_320_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_320_pdest=0x%0h while the rhs_.io_diffCommits_info_320_pdest=0x%0h",this.io_diffCommits_info_320_pdest,rhs_.io_diffCommits_info_320_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_321_ldest!=rhs_.io_diffCommits_info_321_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_321_ldest=0x%0h while the rhs_.io_diffCommits_info_321_ldest=0x%0h",this.io_diffCommits_info_321_ldest,rhs_.io_diffCommits_info_321_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_321_pdest!=rhs_.io_diffCommits_info_321_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_321_pdest=0x%0h while the rhs_.io_diffCommits_info_321_pdest=0x%0h",this.io_diffCommits_info_321_pdest,rhs_.io_diffCommits_info_321_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_322_ldest!=rhs_.io_diffCommits_info_322_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_322_ldest=0x%0h while the rhs_.io_diffCommits_info_322_ldest=0x%0h",this.io_diffCommits_info_322_ldest,rhs_.io_diffCommits_info_322_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_322_pdest!=rhs_.io_diffCommits_info_322_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_322_pdest=0x%0h while the rhs_.io_diffCommits_info_322_pdest=0x%0h",this.io_diffCommits_info_322_pdest,rhs_.io_diffCommits_info_322_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_323_ldest!=rhs_.io_diffCommits_info_323_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_323_ldest=0x%0h while the rhs_.io_diffCommits_info_323_ldest=0x%0h",this.io_diffCommits_info_323_ldest,rhs_.io_diffCommits_info_323_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_323_pdest!=rhs_.io_diffCommits_info_323_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_323_pdest=0x%0h while the rhs_.io_diffCommits_info_323_pdest=0x%0h",this.io_diffCommits_info_323_pdest,rhs_.io_diffCommits_info_323_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_324_ldest!=rhs_.io_diffCommits_info_324_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_324_ldest=0x%0h while the rhs_.io_diffCommits_info_324_ldest=0x%0h",this.io_diffCommits_info_324_ldest,rhs_.io_diffCommits_info_324_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_324_pdest!=rhs_.io_diffCommits_info_324_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_324_pdest=0x%0h while the rhs_.io_diffCommits_info_324_pdest=0x%0h",this.io_diffCommits_info_324_pdest,rhs_.io_diffCommits_info_324_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_325_ldest!=rhs_.io_diffCommits_info_325_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_325_ldest=0x%0h while the rhs_.io_diffCommits_info_325_ldest=0x%0h",this.io_diffCommits_info_325_ldest,rhs_.io_diffCommits_info_325_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_325_pdest!=rhs_.io_diffCommits_info_325_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_325_pdest=0x%0h while the rhs_.io_diffCommits_info_325_pdest=0x%0h",this.io_diffCommits_info_325_pdest,rhs_.io_diffCommits_info_325_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_326_ldest!=rhs_.io_diffCommits_info_326_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_326_ldest=0x%0h while the rhs_.io_diffCommits_info_326_ldest=0x%0h",this.io_diffCommits_info_326_ldest,rhs_.io_diffCommits_info_326_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_326_pdest!=rhs_.io_diffCommits_info_326_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_326_pdest=0x%0h while the rhs_.io_diffCommits_info_326_pdest=0x%0h",this.io_diffCommits_info_326_pdest,rhs_.io_diffCommits_info_326_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_327_ldest!=rhs_.io_diffCommits_info_327_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_327_ldest=0x%0h while the rhs_.io_diffCommits_info_327_ldest=0x%0h",this.io_diffCommits_info_327_ldest,rhs_.io_diffCommits_info_327_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_327_pdest!=rhs_.io_diffCommits_info_327_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_327_pdest=0x%0h while the rhs_.io_diffCommits_info_327_pdest=0x%0h",this.io_diffCommits_info_327_pdest,rhs_.io_diffCommits_info_327_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_328_ldest!=rhs_.io_diffCommits_info_328_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_328_ldest=0x%0h while the rhs_.io_diffCommits_info_328_ldest=0x%0h",this.io_diffCommits_info_328_ldest,rhs_.io_diffCommits_info_328_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_328_pdest!=rhs_.io_diffCommits_info_328_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_328_pdest=0x%0h while the rhs_.io_diffCommits_info_328_pdest=0x%0h",this.io_diffCommits_info_328_pdest,rhs_.io_diffCommits_info_328_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_329_ldest!=rhs_.io_diffCommits_info_329_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_329_ldest=0x%0h while the rhs_.io_diffCommits_info_329_ldest=0x%0h",this.io_diffCommits_info_329_ldest,rhs_.io_diffCommits_info_329_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_329_pdest!=rhs_.io_diffCommits_info_329_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_329_pdest=0x%0h while the rhs_.io_diffCommits_info_329_pdest=0x%0h",this.io_diffCommits_info_329_pdest,rhs_.io_diffCommits_info_329_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_330_ldest!=rhs_.io_diffCommits_info_330_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_330_ldest=0x%0h while the rhs_.io_diffCommits_info_330_ldest=0x%0h",this.io_diffCommits_info_330_ldest,rhs_.io_diffCommits_info_330_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_330_pdest!=rhs_.io_diffCommits_info_330_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_330_pdest=0x%0h while the rhs_.io_diffCommits_info_330_pdest=0x%0h",this.io_diffCommits_info_330_pdest,rhs_.io_diffCommits_info_330_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_331_ldest!=rhs_.io_diffCommits_info_331_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_331_ldest=0x%0h while the rhs_.io_diffCommits_info_331_ldest=0x%0h",this.io_diffCommits_info_331_ldest,rhs_.io_diffCommits_info_331_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_331_pdest!=rhs_.io_diffCommits_info_331_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_331_pdest=0x%0h while the rhs_.io_diffCommits_info_331_pdest=0x%0h",this.io_diffCommits_info_331_pdest,rhs_.io_diffCommits_info_331_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_332_ldest!=rhs_.io_diffCommits_info_332_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_332_ldest=0x%0h while the rhs_.io_diffCommits_info_332_ldest=0x%0h",this.io_diffCommits_info_332_ldest,rhs_.io_diffCommits_info_332_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_332_pdest!=rhs_.io_diffCommits_info_332_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_332_pdest=0x%0h while the rhs_.io_diffCommits_info_332_pdest=0x%0h",this.io_diffCommits_info_332_pdest,rhs_.io_diffCommits_info_332_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_333_ldest!=rhs_.io_diffCommits_info_333_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_333_ldest=0x%0h while the rhs_.io_diffCommits_info_333_ldest=0x%0h",this.io_diffCommits_info_333_ldest,rhs_.io_diffCommits_info_333_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_333_pdest!=rhs_.io_diffCommits_info_333_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_333_pdest=0x%0h while the rhs_.io_diffCommits_info_333_pdest=0x%0h",this.io_diffCommits_info_333_pdest,rhs_.io_diffCommits_info_333_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_334_ldest!=rhs_.io_diffCommits_info_334_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_334_ldest=0x%0h while the rhs_.io_diffCommits_info_334_ldest=0x%0h",this.io_diffCommits_info_334_ldest,rhs_.io_diffCommits_info_334_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_334_pdest!=rhs_.io_diffCommits_info_334_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_334_pdest=0x%0h while the rhs_.io_diffCommits_info_334_pdest=0x%0h",this.io_diffCommits_info_334_pdest,rhs_.io_diffCommits_info_334_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_335_ldest!=rhs_.io_diffCommits_info_335_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_335_ldest=0x%0h while the rhs_.io_diffCommits_info_335_ldest=0x%0h",this.io_diffCommits_info_335_ldest,rhs_.io_diffCommits_info_335_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_335_pdest!=rhs_.io_diffCommits_info_335_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_335_pdest=0x%0h while the rhs_.io_diffCommits_info_335_pdest=0x%0h",this.io_diffCommits_info_335_pdest,rhs_.io_diffCommits_info_335_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_336_ldest!=rhs_.io_diffCommits_info_336_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_336_ldest=0x%0h while the rhs_.io_diffCommits_info_336_ldest=0x%0h",this.io_diffCommits_info_336_ldest,rhs_.io_diffCommits_info_336_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_336_pdest!=rhs_.io_diffCommits_info_336_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_336_pdest=0x%0h while the rhs_.io_diffCommits_info_336_pdest=0x%0h",this.io_diffCommits_info_336_pdest,rhs_.io_diffCommits_info_336_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_337_ldest!=rhs_.io_diffCommits_info_337_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_337_ldest=0x%0h while the rhs_.io_diffCommits_info_337_ldest=0x%0h",this.io_diffCommits_info_337_ldest,rhs_.io_diffCommits_info_337_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_337_pdest!=rhs_.io_diffCommits_info_337_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_337_pdest=0x%0h while the rhs_.io_diffCommits_info_337_pdest=0x%0h",this.io_diffCommits_info_337_pdest,rhs_.io_diffCommits_info_337_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_338_ldest!=rhs_.io_diffCommits_info_338_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_338_ldest=0x%0h while the rhs_.io_diffCommits_info_338_ldest=0x%0h",this.io_diffCommits_info_338_ldest,rhs_.io_diffCommits_info_338_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_338_pdest!=rhs_.io_diffCommits_info_338_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_338_pdest=0x%0h while the rhs_.io_diffCommits_info_338_pdest=0x%0h",this.io_diffCommits_info_338_pdest,rhs_.io_diffCommits_info_338_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_339_ldest!=rhs_.io_diffCommits_info_339_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_339_ldest=0x%0h while the rhs_.io_diffCommits_info_339_ldest=0x%0h",this.io_diffCommits_info_339_ldest,rhs_.io_diffCommits_info_339_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_339_pdest!=rhs_.io_diffCommits_info_339_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_339_pdest=0x%0h while the rhs_.io_diffCommits_info_339_pdest=0x%0h",this.io_diffCommits_info_339_pdest,rhs_.io_diffCommits_info_339_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_340_ldest!=rhs_.io_diffCommits_info_340_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_340_ldest=0x%0h while the rhs_.io_diffCommits_info_340_ldest=0x%0h",this.io_diffCommits_info_340_ldest,rhs_.io_diffCommits_info_340_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_340_pdest!=rhs_.io_diffCommits_info_340_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_340_pdest=0x%0h while the rhs_.io_diffCommits_info_340_pdest=0x%0h",this.io_diffCommits_info_340_pdest,rhs_.io_diffCommits_info_340_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_341_ldest!=rhs_.io_diffCommits_info_341_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_341_ldest=0x%0h while the rhs_.io_diffCommits_info_341_ldest=0x%0h",this.io_diffCommits_info_341_ldest,rhs_.io_diffCommits_info_341_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_341_pdest!=rhs_.io_diffCommits_info_341_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_341_pdest=0x%0h while the rhs_.io_diffCommits_info_341_pdest=0x%0h",this.io_diffCommits_info_341_pdest,rhs_.io_diffCommits_info_341_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_342_ldest!=rhs_.io_diffCommits_info_342_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_342_ldest=0x%0h while the rhs_.io_diffCommits_info_342_ldest=0x%0h",this.io_diffCommits_info_342_ldest,rhs_.io_diffCommits_info_342_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_342_pdest!=rhs_.io_diffCommits_info_342_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_342_pdest=0x%0h while the rhs_.io_diffCommits_info_342_pdest=0x%0h",this.io_diffCommits_info_342_pdest,rhs_.io_diffCommits_info_342_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_343_ldest!=rhs_.io_diffCommits_info_343_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_343_ldest=0x%0h while the rhs_.io_diffCommits_info_343_ldest=0x%0h",this.io_diffCommits_info_343_ldest,rhs_.io_diffCommits_info_343_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_343_pdest!=rhs_.io_diffCommits_info_343_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_343_pdest=0x%0h while the rhs_.io_diffCommits_info_343_pdest=0x%0h",this.io_diffCommits_info_343_pdest,rhs_.io_diffCommits_info_343_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_344_ldest!=rhs_.io_diffCommits_info_344_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_344_ldest=0x%0h while the rhs_.io_diffCommits_info_344_ldest=0x%0h",this.io_diffCommits_info_344_ldest,rhs_.io_diffCommits_info_344_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_344_pdest!=rhs_.io_diffCommits_info_344_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_344_pdest=0x%0h while the rhs_.io_diffCommits_info_344_pdest=0x%0h",this.io_diffCommits_info_344_pdest,rhs_.io_diffCommits_info_344_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_345_ldest!=rhs_.io_diffCommits_info_345_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_345_ldest=0x%0h while the rhs_.io_diffCommits_info_345_ldest=0x%0h",this.io_diffCommits_info_345_ldest,rhs_.io_diffCommits_info_345_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_345_pdest!=rhs_.io_diffCommits_info_345_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_345_pdest=0x%0h while the rhs_.io_diffCommits_info_345_pdest=0x%0h",this.io_diffCommits_info_345_pdest,rhs_.io_diffCommits_info_345_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_346_ldest!=rhs_.io_diffCommits_info_346_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_346_ldest=0x%0h while the rhs_.io_diffCommits_info_346_ldest=0x%0h",this.io_diffCommits_info_346_ldest,rhs_.io_diffCommits_info_346_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_346_pdest!=rhs_.io_diffCommits_info_346_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_346_pdest=0x%0h while the rhs_.io_diffCommits_info_346_pdest=0x%0h",this.io_diffCommits_info_346_pdest,rhs_.io_diffCommits_info_346_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_347_ldest!=rhs_.io_diffCommits_info_347_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_347_ldest=0x%0h while the rhs_.io_diffCommits_info_347_ldest=0x%0h",this.io_diffCommits_info_347_ldest,rhs_.io_diffCommits_info_347_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_347_pdest!=rhs_.io_diffCommits_info_347_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_347_pdest=0x%0h while the rhs_.io_diffCommits_info_347_pdest=0x%0h",this.io_diffCommits_info_347_pdest,rhs_.io_diffCommits_info_347_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_348_ldest!=rhs_.io_diffCommits_info_348_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_348_ldest=0x%0h while the rhs_.io_diffCommits_info_348_ldest=0x%0h",this.io_diffCommits_info_348_ldest,rhs_.io_diffCommits_info_348_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_348_pdest!=rhs_.io_diffCommits_info_348_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_348_pdest=0x%0h while the rhs_.io_diffCommits_info_348_pdest=0x%0h",this.io_diffCommits_info_348_pdest,rhs_.io_diffCommits_info_348_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_349_ldest!=rhs_.io_diffCommits_info_349_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_349_ldest=0x%0h while the rhs_.io_diffCommits_info_349_ldest=0x%0h",this.io_diffCommits_info_349_ldest,rhs_.io_diffCommits_info_349_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_349_pdest!=rhs_.io_diffCommits_info_349_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_349_pdest=0x%0h while the rhs_.io_diffCommits_info_349_pdest=0x%0h",this.io_diffCommits_info_349_pdest,rhs_.io_diffCommits_info_349_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_350_ldest!=rhs_.io_diffCommits_info_350_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_350_ldest=0x%0h while the rhs_.io_diffCommits_info_350_ldest=0x%0h",this.io_diffCommits_info_350_ldest,rhs_.io_diffCommits_info_350_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_350_pdest!=rhs_.io_diffCommits_info_350_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_350_pdest=0x%0h while the rhs_.io_diffCommits_info_350_pdest=0x%0h",this.io_diffCommits_info_350_pdest,rhs_.io_diffCommits_info_350_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_351_ldest!=rhs_.io_diffCommits_info_351_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_351_ldest=0x%0h while the rhs_.io_diffCommits_info_351_ldest=0x%0h",this.io_diffCommits_info_351_ldest,rhs_.io_diffCommits_info_351_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_351_pdest!=rhs_.io_diffCommits_info_351_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_351_pdest=0x%0h while the rhs_.io_diffCommits_info_351_pdest=0x%0h",this.io_diffCommits_info_351_pdest,rhs_.io_diffCommits_info_351_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_352_ldest!=rhs_.io_diffCommits_info_352_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_352_ldest=0x%0h while the rhs_.io_diffCommits_info_352_ldest=0x%0h",this.io_diffCommits_info_352_ldest,rhs_.io_diffCommits_info_352_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_352_pdest!=rhs_.io_diffCommits_info_352_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_352_pdest=0x%0h while the rhs_.io_diffCommits_info_352_pdest=0x%0h",this.io_diffCommits_info_352_pdest,rhs_.io_diffCommits_info_352_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_353_ldest!=rhs_.io_diffCommits_info_353_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_353_ldest=0x%0h while the rhs_.io_diffCommits_info_353_ldest=0x%0h",this.io_diffCommits_info_353_ldest,rhs_.io_diffCommits_info_353_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_353_pdest!=rhs_.io_diffCommits_info_353_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_353_pdest=0x%0h while the rhs_.io_diffCommits_info_353_pdest=0x%0h",this.io_diffCommits_info_353_pdest,rhs_.io_diffCommits_info_353_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_354_ldest!=rhs_.io_diffCommits_info_354_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_354_ldest=0x%0h while the rhs_.io_diffCommits_info_354_ldest=0x%0h",this.io_diffCommits_info_354_ldest,rhs_.io_diffCommits_info_354_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_354_pdest!=rhs_.io_diffCommits_info_354_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_354_pdest=0x%0h while the rhs_.io_diffCommits_info_354_pdest=0x%0h",this.io_diffCommits_info_354_pdest,rhs_.io_diffCommits_info_354_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_355_ldest!=rhs_.io_diffCommits_info_355_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_355_ldest=0x%0h while the rhs_.io_diffCommits_info_355_ldest=0x%0h",this.io_diffCommits_info_355_ldest,rhs_.io_diffCommits_info_355_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_355_pdest!=rhs_.io_diffCommits_info_355_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_355_pdest=0x%0h while the rhs_.io_diffCommits_info_355_pdest=0x%0h",this.io_diffCommits_info_355_pdest,rhs_.io_diffCommits_info_355_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_356_ldest!=rhs_.io_diffCommits_info_356_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_356_ldest=0x%0h while the rhs_.io_diffCommits_info_356_ldest=0x%0h",this.io_diffCommits_info_356_ldest,rhs_.io_diffCommits_info_356_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_356_pdest!=rhs_.io_diffCommits_info_356_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_356_pdest=0x%0h while the rhs_.io_diffCommits_info_356_pdest=0x%0h",this.io_diffCommits_info_356_pdest,rhs_.io_diffCommits_info_356_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_357_ldest!=rhs_.io_diffCommits_info_357_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_357_ldest=0x%0h while the rhs_.io_diffCommits_info_357_ldest=0x%0h",this.io_diffCommits_info_357_ldest,rhs_.io_diffCommits_info_357_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_357_pdest!=rhs_.io_diffCommits_info_357_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_357_pdest=0x%0h while the rhs_.io_diffCommits_info_357_pdest=0x%0h",this.io_diffCommits_info_357_pdest,rhs_.io_diffCommits_info_357_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_358_ldest!=rhs_.io_diffCommits_info_358_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_358_ldest=0x%0h while the rhs_.io_diffCommits_info_358_ldest=0x%0h",this.io_diffCommits_info_358_ldest,rhs_.io_diffCommits_info_358_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_358_pdest!=rhs_.io_diffCommits_info_358_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_358_pdest=0x%0h while the rhs_.io_diffCommits_info_358_pdest=0x%0h",this.io_diffCommits_info_358_pdest,rhs_.io_diffCommits_info_358_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_359_ldest!=rhs_.io_diffCommits_info_359_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_359_ldest=0x%0h while the rhs_.io_diffCommits_info_359_ldest=0x%0h",this.io_diffCommits_info_359_ldest,rhs_.io_diffCommits_info_359_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_359_pdest!=rhs_.io_diffCommits_info_359_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_359_pdest=0x%0h while the rhs_.io_diffCommits_info_359_pdest=0x%0h",this.io_diffCommits_info_359_pdest,rhs_.io_diffCommits_info_359_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_360_ldest!=rhs_.io_diffCommits_info_360_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_360_ldest=0x%0h while the rhs_.io_diffCommits_info_360_ldest=0x%0h",this.io_diffCommits_info_360_ldest,rhs_.io_diffCommits_info_360_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_360_pdest!=rhs_.io_diffCommits_info_360_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_360_pdest=0x%0h while the rhs_.io_diffCommits_info_360_pdest=0x%0h",this.io_diffCommits_info_360_pdest,rhs_.io_diffCommits_info_360_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_361_ldest!=rhs_.io_diffCommits_info_361_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_361_ldest=0x%0h while the rhs_.io_diffCommits_info_361_ldest=0x%0h",this.io_diffCommits_info_361_ldest,rhs_.io_diffCommits_info_361_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_361_pdest!=rhs_.io_diffCommits_info_361_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_361_pdest=0x%0h while the rhs_.io_diffCommits_info_361_pdest=0x%0h",this.io_diffCommits_info_361_pdest,rhs_.io_diffCommits_info_361_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_362_ldest!=rhs_.io_diffCommits_info_362_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_362_ldest=0x%0h while the rhs_.io_diffCommits_info_362_ldest=0x%0h",this.io_diffCommits_info_362_ldest,rhs_.io_diffCommits_info_362_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_362_pdest!=rhs_.io_diffCommits_info_362_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_362_pdest=0x%0h while the rhs_.io_diffCommits_info_362_pdest=0x%0h",this.io_diffCommits_info_362_pdest,rhs_.io_diffCommits_info_362_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_363_ldest!=rhs_.io_diffCommits_info_363_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_363_ldest=0x%0h while the rhs_.io_diffCommits_info_363_ldest=0x%0h",this.io_diffCommits_info_363_ldest,rhs_.io_diffCommits_info_363_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_363_pdest!=rhs_.io_diffCommits_info_363_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_363_pdest=0x%0h while the rhs_.io_diffCommits_info_363_pdest=0x%0h",this.io_diffCommits_info_363_pdest,rhs_.io_diffCommits_info_363_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_364_ldest!=rhs_.io_diffCommits_info_364_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_364_ldest=0x%0h while the rhs_.io_diffCommits_info_364_ldest=0x%0h",this.io_diffCommits_info_364_ldest,rhs_.io_diffCommits_info_364_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_364_pdest!=rhs_.io_diffCommits_info_364_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_364_pdest=0x%0h while the rhs_.io_diffCommits_info_364_pdest=0x%0h",this.io_diffCommits_info_364_pdest,rhs_.io_diffCommits_info_364_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_365_ldest!=rhs_.io_diffCommits_info_365_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_365_ldest=0x%0h while the rhs_.io_diffCommits_info_365_ldest=0x%0h",this.io_diffCommits_info_365_ldest,rhs_.io_diffCommits_info_365_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_365_pdest!=rhs_.io_diffCommits_info_365_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_365_pdest=0x%0h while the rhs_.io_diffCommits_info_365_pdest=0x%0h",this.io_diffCommits_info_365_pdest,rhs_.io_diffCommits_info_365_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_366_ldest!=rhs_.io_diffCommits_info_366_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_366_ldest=0x%0h while the rhs_.io_diffCommits_info_366_ldest=0x%0h",this.io_diffCommits_info_366_ldest,rhs_.io_diffCommits_info_366_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_366_pdest!=rhs_.io_diffCommits_info_366_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_366_pdest=0x%0h while the rhs_.io_diffCommits_info_366_pdest=0x%0h",this.io_diffCommits_info_366_pdest,rhs_.io_diffCommits_info_366_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_367_ldest!=rhs_.io_diffCommits_info_367_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_367_ldest=0x%0h while the rhs_.io_diffCommits_info_367_ldest=0x%0h",this.io_diffCommits_info_367_ldest,rhs_.io_diffCommits_info_367_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_367_pdest!=rhs_.io_diffCommits_info_367_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_367_pdest=0x%0h while the rhs_.io_diffCommits_info_367_pdest=0x%0h",this.io_diffCommits_info_367_pdest,rhs_.io_diffCommits_info_367_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_368_ldest!=rhs_.io_diffCommits_info_368_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_368_ldest=0x%0h while the rhs_.io_diffCommits_info_368_ldest=0x%0h",this.io_diffCommits_info_368_ldest,rhs_.io_diffCommits_info_368_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_368_pdest!=rhs_.io_diffCommits_info_368_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_368_pdest=0x%0h while the rhs_.io_diffCommits_info_368_pdest=0x%0h",this.io_diffCommits_info_368_pdest,rhs_.io_diffCommits_info_368_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_369_ldest!=rhs_.io_diffCommits_info_369_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_369_ldest=0x%0h while the rhs_.io_diffCommits_info_369_ldest=0x%0h",this.io_diffCommits_info_369_ldest,rhs_.io_diffCommits_info_369_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_369_pdest!=rhs_.io_diffCommits_info_369_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_369_pdest=0x%0h while the rhs_.io_diffCommits_info_369_pdest=0x%0h",this.io_diffCommits_info_369_pdest,rhs_.io_diffCommits_info_369_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_370_ldest!=rhs_.io_diffCommits_info_370_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_370_ldest=0x%0h while the rhs_.io_diffCommits_info_370_ldest=0x%0h",this.io_diffCommits_info_370_ldest,rhs_.io_diffCommits_info_370_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_370_pdest!=rhs_.io_diffCommits_info_370_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_370_pdest=0x%0h while the rhs_.io_diffCommits_info_370_pdest=0x%0h",this.io_diffCommits_info_370_pdest,rhs_.io_diffCommits_info_370_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_371_ldest!=rhs_.io_diffCommits_info_371_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_371_ldest=0x%0h while the rhs_.io_diffCommits_info_371_ldest=0x%0h",this.io_diffCommits_info_371_ldest,rhs_.io_diffCommits_info_371_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_371_pdest!=rhs_.io_diffCommits_info_371_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_371_pdest=0x%0h while the rhs_.io_diffCommits_info_371_pdest=0x%0h",this.io_diffCommits_info_371_pdest,rhs_.io_diffCommits_info_371_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_372_ldest!=rhs_.io_diffCommits_info_372_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_372_ldest=0x%0h while the rhs_.io_diffCommits_info_372_ldest=0x%0h",this.io_diffCommits_info_372_ldest,rhs_.io_diffCommits_info_372_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_372_pdest!=rhs_.io_diffCommits_info_372_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_372_pdest=0x%0h while the rhs_.io_diffCommits_info_372_pdest=0x%0h",this.io_diffCommits_info_372_pdest,rhs_.io_diffCommits_info_372_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_373_ldest!=rhs_.io_diffCommits_info_373_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_373_ldest=0x%0h while the rhs_.io_diffCommits_info_373_ldest=0x%0h",this.io_diffCommits_info_373_ldest,rhs_.io_diffCommits_info_373_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_373_pdest!=rhs_.io_diffCommits_info_373_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_373_pdest=0x%0h while the rhs_.io_diffCommits_info_373_pdest=0x%0h",this.io_diffCommits_info_373_pdest,rhs_.io_diffCommits_info_373_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_374_ldest!=rhs_.io_diffCommits_info_374_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_374_ldest=0x%0h while the rhs_.io_diffCommits_info_374_ldest=0x%0h",this.io_diffCommits_info_374_ldest,rhs_.io_diffCommits_info_374_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_374_pdest!=rhs_.io_diffCommits_info_374_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_374_pdest=0x%0h while the rhs_.io_diffCommits_info_374_pdest=0x%0h",this.io_diffCommits_info_374_pdest,rhs_.io_diffCommits_info_374_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_375_ldest!=rhs_.io_diffCommits_info_375_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_375_ldest=0x%0h while the rhs_.io_diffCommits_info_375_ldest=0x%0h",this.io_diffCommits_info_375_ldest,rhs_.io_diffCommits_info_375_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_375_pdest!=rhs_.io_diffCommits_info_375_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_375_pdest=0x%0h while the rhs_.io_diffCommits_info_375_pdest=0x%0h",this.io_diffCommits_info_375_pdest,rhs_.io_diffCommits_info_375_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_376_ldest!=rhs_.io_diffCommits_info_376_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_376_ldest=0x%0h while the rhs_.io_diffCommits_info_376_ldest=0x%0h",this.io_diffCommits_info_376_ldest,rhs_.io_diffCommits_info_376_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_376_pdest!=rhs_.io_diffCommits_info_376_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_376_pdest=0x%0h while the rhs_.io_diffCommits_info_376_pdest=0x%0h",this.io_diffCommits_info_376_pdest,rhs_.io_diffCommits_info_376_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_377_ldest!=rhs_.io_diffCommits_info_377_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_377_ldest=0x%0h while the rhs_.io_diffCommits_info_377_ldest=0x%0h",this.io_diffCommits_info_377_ldest,rhs_.io_diffCommits_info_377_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_377_pdest!=rhs_.io_diffCommits_info_377_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_377_pdest=0x%0h while the rhs_.io_diffCommits_info_377_pdest=0x%0h",this.io_diffCommits_info_377_pdest,rhs_.io_diffCommits_info_377_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_378_ldest!=rhs_.io_diffCommits_info_378_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_378_ldest=0x%0h while the rhs_.io_diffCommits_info_378_ldest=0x%0h",this.io_diffCommits_info_378_ldest,rhs_.io_diffCommits_info_378_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_378_pdest!=rhs_.io_diffCommits_info_378_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_378_pdest=0x%0h while the rhs_.io_diffCommits_info_378_pdest=0x%0h",this.io_diffCommits_info_378_pdest,rhs_.io_diffCommits_info_378_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_379_ldest!=rhs_.io_diffCommits_info_379_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_379_ldest=0x%0h while the rhs_.io_diffCommits_info_379_ldest=0x%0h",this.io_diffCommits_info_379_ldest,rhs_.io_diffCommits_info_379_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_379_pdest!=rhs_.io_diffCommits_info_379_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_379_pdest=0x%0h while the rhs_.io_diffCommits_info_379_pdest=0x%0h",this.io_diffCommits_info_379_pdest,rhs_.io_diffCommits_info_379_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_380_ldest!=rhs_.io_diffCommits_info_380_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_380_ldest=0x%0h while the rhs_.io_diffCommits_info_380_ldest=0x%0h",this.io_diffCommits_info_380_ldest,rhs_.io_diffCommits_info_380_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_380_pdest!=rhs_.io_diffCommits_info_380_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_380_pdest=0x%0h while the rhs_.io_diffCommits_info_380_pdest=0x%0h",this.io_diffCommits_info_380_pdest,rhs_.io_diffCommits_info_380_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_381_ldest!=rhs_.io_diffCommits_info_381_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_381_ldest=0x%0h while the rhs_.io_diffCommits_info_381_ldest=0x%0h",this.io_diffCommits_info_381_ldest,rhs_.io_diffCommits_info_381_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_381_pdest!=rhs_.io_diffCommits_info_381_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_381_pdest=0x%0h while the rhs_.io_diffCommits_info_381_pdest=0x%0h",this.io_diffCommits_info_381_pdest,rhs_.io_diffCommits_info_381_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_382_ldest!=rhs_.io_diffCommits_info_382_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_382_ldest=0x%0h while the rhs_.io_diffCommits_info_382_ldest=0x%0h",this.io_diffCommits_info_382_ldest,rhs_.io_diffCommits_info_382_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_382_pdest!=rhs_.io_diffCommits_info_382_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_382_pdest=0x%0h while the rhs_.io_diffCommits_info_382_pdest=0x%0h",this.io_diffCommits_info_382_pdest,rhs_.io_diffCommits_info_382_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_383_ldest!=rhs_.io_diffCommits_info_383_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_383_ldest=0x%0h while the rhs_.io_diffCommits_info_383_ldest=0x%0h",this.io_diffCommits_info_383_ldest,rhs_.io_diffCommits_info_383_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_383_pdest!=rhs_.io_diffCommits_info_383_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_383_pdest=0x%0h while the rhs_.io_diffCommits_info_383_pdest=0x%0h",this.io_diffCommits_info_383_pdest,rhs_.io_diffCommits_info_383_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_384_ldest!=rhs_.io_diffCommits_info_384_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_384_ldest=0x%0h while the rhs_.io_diffCommits_info_384_ldest=0x%0h",this.io_diffCommits_info_384_ldest,rhs_.io_diffCommits_info_384_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_384_pdest!=rhs_.io_diffCommits_info_384_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_384_pdest=0x%0h while the rhs_.io_diffCommits_info_384_pdest=0x%0h",this.io_diffCommits_info_384_pdest,rhs_.io_diffCommits_info_384_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_385_ldest!=rhs_.io_diffCommits_info_385_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_385_ldest=0x%0h while the rhs_.io_diffCommits_info_385_ldest=0x%0h",this.io_diffCommits_info_385_ldest,rhs_.io_diffCommits_info_385_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_385_pdest!=rhs_.io_diffCommits_info_385_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_385_pdest=0x%0h while the rhs_.io_diffCommits_info_385_pdest=0x%0h",this.io_diffCommits_info_385_pdest,rhs_.io_diffCommits_info_385_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_386_ldest!=rhs_.io_diffCommits_info_386_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_386_ldest=0x%0h while the rhs_.io_diffCommits_info_386_ldest=0x%0h",this.io_diffCommits_info_386_ldest,rhs_.io_diffCommits_info_386_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_386_pdest!=rhs_.io_diffCommits_info_386_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_386_pdest=0x%0h while the rhs_.io_diffCommits_info_386_pdest=0x%0h",this.io_diffCommits_info_386_pdest,rhs_.io_diffCommits_info_386_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_387_ldest!=rhs_.io_diffCommits_info_387_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_387_ldest=0x%0h while the rhs_.io_diffCommits_info_387_ldest=0x%0h",this.io_diffCommits_info_387_ldest,rhs_.io_diffCommits_info_387_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_387_pdest!=rhs_.io_diffCommits_info_387_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_387_pdest=0x%0h while the rhs_.io_diffCommits_info_387_pdest=0x%0h",this.io_diffCommits_info_387_pdest,rhs_.io_diffCommits_info_387_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_388_ldest!=rhs_.io_diffCommits_info_388_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_388_ldest=0x%0h while the rhs_.io_diffCommits_info_388_ldest=0x%0h",this.io_diffCommits_info_388_ldest,rhs_.io_diffCommits_info_388_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_388_pdest!=rhs_.io_diffCommits_info_388_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_388_pdest=0x%0h while the rhs_.io_diffCommits_info_388_pdest=0x%0h",this.io_diffCommits_info_388_pdest,rhs_.io_diffCommits_info_388_pdest),UVM_NONE)
        end

        if(this.io_diffCommits_info_389_ldest!=rhs_.io_diffCommits_info_389_ldest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_389_ldest=0x%0h while the rhs_.io_diffCommits_info_389_ldest=0x%0h",this.io_diffCommits_info_389_ldest,rhs_.io_diffCommits_info_389_ldest),UVM_NONE)
        end

        if(this.io_diffCommits_info_389_pdest!=rhs_.io_diffCommits_info_389_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_diffCommits_info_389_pdest=0x%0h while the rhs_.io_diffCommits_info_389_pdest=0x%0h",this.io_diffCommits_info_389_pdest,rhs_.io_diffCommits_info_389_pdest),UVM_NONE)
        end

        if(this.io_lsq_scommit!=rhs_.io_lsq_scommit) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_lsq_scommit=0x%0h while the rhs_.io_lsq_scommit=0x%0h",this.io_lsq_scommit,rhs_.io_lsq_scommit),UVM_NONE)
        end

        if(this.io_lsq_pendingMMIOld!=rhs_.io_lsq_pendingMMIOld) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_lsq_pendingMMIOld=0x%0h while the rhs_.io_lsq_pendingMMIOld=0x%0h",this.io_lsq_pendingMMIOld,rhs_.io_lsq_pendingMMIOld),UVM_NONE)
        end

        if(this.io_lsq_pendingst!=rhs_.io_lsq_pendingst) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_lsq_pendingst=0x%0h while the rhs_.io_lsq_pendingst=0x%0h",this.io_lsq_pendingst,rhs_.io_lsq_pendingst),UVM_NONE)
        end

        if(this.io_lsq_pendingPtr_flag!=rhs_.io_lsq_pendingPtr_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_lsq_pendingPtr_flag=0x%0h while the rhs_.io_lsq_pendingPtr_flag=0x%0h",this.io_lsq_pendingPtr_flag,rhs_.io_lsq_pendingPtr_flag),UVM_NONE)
        end

        if(this.io_lsq_pendingPtr_value!=rhs_.io_lsq_pendingPtr_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_lsq_pendingPtr_value=0x%0h while the rhs_.io_lsq_pendingPtr_value=0x%0h",this.io_lsq_pendingPtr_value,rhs_.io_lsq_pendingPtr_value),UVM_NONE)
        end

        if(this.io_robDeqPtr_flag!=rhs_.io_robDeqPtr_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_robDeqPtr_flag=0x%0h while the rhs_.io_robDeqPtr_flag=0x%0h",this.io_robDeqPtr_flag,rhs_.io_robDeqPtr_flag),UVM_NONE)
        end

        if(this.io_robDeqPtr_value!=rhs_.io_robDeqPtr_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_robDeqPtr_value=0x%0h while the rhs_.io_robDeqPtr_value=0x%0h",this.io_robDeqPtr_value,rhs_.io_robDeqPtr_value),UVM_NONE)
        end

        if(this.io_csr_fflags_valid!=rhs_.io_csr_fflags_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_csr_fflags_valid=0x%0h while the rhs_.io_csr_fflags_valid=0x%0h",this.io_csr_fflags_valid,rhs_.io_csr_fflags_valid),UVM_NONE)
        end

        if(this.io_csr_fflags_bits!=rhs_.io_csr_fflags_bits) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_csr_fflags_bits=0x%0h while the rhs_.io_csr_fflags_bits=0x%0h",this.io_csr_fflags_bits,rhs_.io_csr_fflags_bits),UVM_NONE)
        end

        if(this.io_csr_vxsat_valid!=rhs_.io_csr_vxsat_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_csr_vxsat_valid=0x%0h while the rhs_.io_csr_vxsat_valid=0x%0h",this.io_csr_vxsat_valid,rhs_.io_csr_vxsat_valid),UVM_NONE)
        end

        if(this.io_csr_vxsat_bits!=rhs_.io_csr_vxsat_bits) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_csr_vxsat_bits=0x%0h while the rhs_.io_csr_vxsat_bits=0x%0h",this.io_csr_vxsat_bits,rhs_.io_csr_vxsat_bits),UVM_NONE)
        end

        if(this.io_csr_vstart_valid!=rhs_.io_csr_vstart_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_csr_vstart_valid=0x%0h while the rhs_.io_csr_vstart_valid=0x%0h",this.io_csr_vstart_valid,rhs_.io_csr_vstart_valid),UVM_NONE)
        end

        if(this.io_csr_vstart_bits!=rhs_.io_csr_vstart_bits) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_csr_vstart_bits=0x%0h while the rhs_.io_csr_vstart_bits=0x%0h",this.io_csr_vstart_bits,rhs_.io_csr_vstart_bits),UVM_NONE)
        end

        if(this.io_csr_dirty_fs!=rhs_.io_csr_dirty_fs) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_csr_dirty_fs=0x%0h while the rhs_.io_csr_dirty_fs=0x%0h",this.io_csr_dirty_fs,rhs_.io_csr_dirty_fs),UVM_NONE)
        end

        if(this.io_csr_dirty_vs!=rhs_.io_csr_dirty_vs) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_csr_dirty_vs=0x%0h while the rhs_.io_csr_dirty_vs=0x%0h",this.io_csr_dirty_vs,rhs_.io_csr_dirty_vs),UVM_NONE)
        end

        if(this.io_csr_perfinfo_retiredInstr!=rhs_.io_csr_perfinfo_retiredInstr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_csr_perfinfo_retiredInstr=0x%0h while the rhs_.io_csr_perfinfo_retiredInstr=0x%0h",this.io_csr_perfinfo_retiredInstr,rhs_.io_csr_perfinfo_retiredInstr),UVM_NONE)
        end

        if(this.io_cpu_halt!=rhs_.io_cpu_halt) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_cpu_halt=0x%0h while the rhs_.io_cpu_halt=0x%0h",this.io_cpu_halt,rhs_.io_cpu_halt),UVM_NONE)
        end

        if(this.io_wfi_wfiReq!=rhs_.io_wfi_wfiReq) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_wfi_wfiReq=0x%0h while the rhs_.io_wfi_wfiReq=0x%0h",this.io_wfi_wfiReq,rhs_.io_wfi_wfiReq),UVM_NONE)
        end

        if(this.io_toDecode_isResumeVType!=rhs_.io_toDecode_isResumeVType) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toDecode_isResumeVType=0x%0h while the rhs_.io_toDecode_isResumeVType=0x%0h",this.io_toDecode_isResumeVType,rhs_.io_toDecode_isResumeVType),UVM_NONE)
        end

        if(this.io_toDecode_walkToArchVType!=rhs_.io_toDecode_walkToArchVType) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toDecode_walkToArchVType=0x%0h while the rhs_.io_toDecode_walkToArchVType=0x%0h",this.io_toDecode_walkToArchVType,rhs_.io_toDecode_walkToArchVType),UVM_NONE)
        end

        if(this.io_toDecode_walkVType_valid!=rhs_.io_toDecode_walkVType_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toDecode_walkVType_valid=0x%0h while the rhs_.io_toDecode_walkVType_valid=0x%0h",this.io_toDecode_walkVType_valid,rhs_.io_toDecode_walkVType_valid),UVM_NONE)
        end

        if(this.io_toDecode_walkVType_bits_illegal!=rhs_.io_toDecode_walkVType_bits_illegal) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toDecode_walkVType_bits_illegal=0x%0h while the rhs_.io_toDecode_walkVType_bits_illegal=0x%0h",this.io_toDecode_walkVType_bits_illegal,rhs_.io_toDecode_walkVType_bits_illegal),UVM_NONE)
        end

        if(this.io_toDecode_walkVType_bits_vma!=rhs_.io_toDecode_walkVType_bits_vma) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toDecode_walkVType_bits_vma=0x%0h while the rhs_.io_toDecode_walkVType_bits_vma=0x%0h",this.io_toDecode_walkVType_bits_vma,rhs_.io_toDecode_walkVType_bits_vma),UVM_NONE)
        end

        if(this.io_toDecode_walkVType_bits_vta!=rhs_.io_toDecode_walkVType_bits_vta) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toDecode_walkVType_bits_vta=0x%0h while the rhs_.io_toDecode_walkVType_bits_vta=0x%0h",this.io_toDecode_walkVType_bits_vta,rhs_.io_toDecode_walkVType_bits_vta),UVM_NONE)
        end

        if(this.io_toDecode_walkVType_bits_vsew!=rhs_.io_toDecode_walkVType_bits_vsew) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toDecode_walkVType_bits_vsew=0x%0h while the rhs_.io_toDecode_walkVType_bits_vsew=0x%0h",this.io_toDecode_walkVType_bits_vsew,rhs_.io_toDecode_walkVType_bits_vsew),UVM_NONE)
        end

        if(this.io_toDecode_walkVType_bits_vlmul!=rhs_.io_toDecode_walkVType_bits_vlmul) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toDecode_walkVType_bits_vlmul=0x%0h while the rhs_.io_toDecode_walkVType_bits_vlmul=0x%0h",this.io_toDecode_walkVType_bits_vlmul,rhs_.io_toDecode_walkVType_bits_vlmul),UVM_NONE)
        end

        if(this.io_toDecode_commitVType_vtype_valid!=rhs_.io_toDecode_commitVType_vtype_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toDecode_commitVType_vtype_valid=0x%0h while the rhs_.io_toDecode_commitVType_vtype_valid=0x%0h",this.io_toDecode_commitVType_vtype_valid,rhs_.io_toDecode_commitVType_vtype_valid),UVM_NONE)
        end

        if(this.io_toDecode_commitVType_vtype_bits_illegal!=rhs_.io_toDecode_commitVType_vtype_bits_illegal) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toDecode_commitVType_vtype_bits_illegal=0x%0h while the rhs_.io_toDecode_commitVType_vtype_bits_illegal=0x%0h",this.io_toDecode_commitVType_vtype_bits_illegal,rhs_.io_toDecode_commitVType_vtype_bits_illegal),UVM_NONE)
        end

        if(this.io_toDecode_commitVType_vtype_bits_vma!=rhs_.io_toDecode_commitVType_vtype_bits_vma) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toDecode_commitVType_vtype_bits_vma=0x%0h while the rhs_.io_toDecode_commitVType_vtype_bits_vma=0x%0h",this.io_toDecode_commitVType_vtype_bits_vma,rhs_.io_toDecode_commitVType_vtype_bits_vma),UVM_NONE)
        end

        if(this.io_toDecode_commitVType_vtype_bits_vta!=rhs_.io_toDecode_commitVType_vtype_bits_vta) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toDecode_commitVType_vtype_bits_vta=0x%0h while the rhs_.io_toDecode_commitVType_vtype_bits_vta=0x%0h",this.io_toDecode_commitVType_vtype_bits_vta,rhs_.io_toDecode_commitVType_vtype_bits_vta),UVM_NONE)
        end

        if(this.io_toDecode_commitVType_vtype_bits_vsew!=rhs_.io_toDecode_commitVType_vtype_bits_vsew) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toDecode_commitVType_vtype_bits_vsew=0x%0h while the rhs_.io_toDecode_commitVType_vtype_bits_vsew=0x%0h",this.io_toDecode_commitVType_vtype_bits_vsew,rhs_.io_toDecode_commitVType_vtype_bits_vsew),UVM_NONE)
        end

        if(this.io_toDecode_commitVType_vtype_bits_vlmul!=rhs_.io_toDecode_commitVType_vtype_bits_vlmul) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toDecode_commitVType_vtype_bits_vlmul=0x%0h while the rhs_.io_toDecode_commitVType_vtype_bits_vlmul=0x%0h",this.io_toDecode_commitVType_vtype_bits_vlmul,rhs_.io_toDecode_commitVType_vtype_bits_vlmul),UVM_NONE)
        end

        if(this.io_toDecode_commitVType_hasVsetvl!=rhs_.io_toDecode_commitVType_hasVsetvl) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toDecode_commitVType_hasVsetvl=0x%0h while the rhs_.io_toDecode_commitVType_hasVsetvl=0x%0h",this.io_toDecode_commitVType_hasVsetvl,rhs_.io_toDecode_commitVType_hasVsetvl),UVM_NONE)
        end

        if(this.io_readGPAMemAddr_valid!=rhs_.io_readGPAMemAddr_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_readGPAMemAddr_valid=0x%0h while the rhs_.io_readGPAMemAddr_valid=0x%0h",this.io_readGPAMemAddr_valid,rhs_.io_readGPAMemAddr_valid),UVM_NONE)
        end

        if(this.io_readGPAMemAddr_bits_ftqPtr_value!=rhs_.io_readGPAMemAddr_bits_ftqPtr_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_readGPAMemAddr_bits_ftqPtr_value=0x%0h while the rhs_.io_readGPAMemAddr_bits_ftqPtr_value=0x%0h",this.io_readGPAMemAddr_bits_ftqPtr_value,rhs_.io_readGPAMemAddr_bits_ftqPtr_value),UVM_NONE)
        end

        if(this.io_readGPAMemAddr_bits_ftqOffset!=rhs_.io_readGPAMemAddr_bits_ftqOffset) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_readGPAMemAddr_bits_ftqOffset=0x%0h while the rhs_.io_readGPAMemAddr_bits_ftqOffset=0x%0h",this.io_readGPAMemAddr_bits_ftqOffset,rhs_.io_readGPAMemAddr_bits_ftqOffset),UVM_NONE)
        end

        if(this.io_toVecExcpMod_logicPhyRegMap_0_valid!=rhs_.io_toVecExcpMod_logicPhyRegMap_0_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toVecExcpMod_logicPhyRegMap_0_valid=0x%0h while the rhs_.io_toVecExcpMod_logicPhyRegMap_0_valid=0x%0h",this.io_toVecExcpMod_logicPhyRegMap_0_valid,rhs_.io_toVecExcpMod_logicPhyRegMap_0_valid),UVM_NONE)
        end

        if(this.io_toVecExcpMod_logicPhyRegMap_0_bits_lreg!=rhs_.io_toVecExcpMod_logicPhyRegMap_0_bits_lreg) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toVecExcpMod_logicPhyRegMap_0_bits_lreg=0x%0h while the rhs_.io_toVecExcpMod_logicPhyRegMap_0_bits_lreg=0x%0h",this.io_toVecExcpMod_logicPhyRegMap_0_bits_lreg,rhs_.io_toVecExcpMod_logicPhyRegMap_0_bits_lreg),UVM_NONE)
        end

        if(this.io_toVecExcpMod_logicPhyRegMap_0_bits_preg!=rhs_.io_toVecExcpMod_logicPhyRegMap_0_bits_preg) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toVecExcpMod_logicPhyRegMap_0_bits_preg=0x%0h while the rhs_.io_toVecExcpMod_logicPhyRegMap_0_bits_preg=0x%0h",this.io_toVecExcpMod_logicPhyRegMap_0_bits_preg,rhs_.io_toVecExcpMod_logicPhyRegMap_0_bits_preg),UVM_NONE)
        end

        if(this.io_toVecExcpMod_logicPhyRegMap_1_valid!=rhs_.io_toVecExcpMod_logicPhyRegMap_1_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toVecExcpMod_logicPhyRegMap_1_valid=0x%0h while the rhs_.io_toVecExcpMod_logicPhyRegMap_1_valid=0x%0h",this.io_toVecExcpMod_logicPhyRegMap_1_valid,rhs_.io_toVecExcpMod_logicPhyRegMap_1_valid),UVM_NONE)
        end

        if(this.io_toVecExcpMod_logicPhyRegMap_1_bits_lreg!=rhs_.io_toVecExcpMod_logicPhyRegMap_1_bits_lreg) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toVecExcpMod_logicPhyRegMap_1_bits_lreg=0x%0h while the rhs_.io_toVecExcpMod_logicPhyRegMap_1_bits_lreg=0x%0h",this.io_toVecExcpMod_logicPhyRegMap_1_bits_lreg,rhs_.io_toVecExcpMod_logicPhyRegMap_1_bits_lreg),UVM_NONE)
        end

        if(this.io_toVecExcpMod_logicPhyRegMap_1_bits_preg!=rhs_.io_toVecExcpMod_logicPhyRegMap_1_bits_preg) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toVecExcpMod_logicPhyRegMap_1_bits_preg=0x%0h while the rhs_.io_toVecExcpMod_logicPhyRegMap_1_bits_preg=0x%0h",this.io_toVecExcpMod_logicPhyRegMap_1_bits_preg,rhs_.io_toVecExcpMod_logicPhyRegMap_1_bits_preg),UVM_NONE)
        end

        if(this.io_toVecExcpMod_logicPhyRegMap_2_valid!=rhs_.io_toVecExcpMod_logicPhyRegMap_2_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toVecExcpMod_logicPhyRegMap_2_valid=0x%0h while the rhs_.io_toVecExcpMod_logicPhyRegMap_2_valid=0x%0h",this.io_toVecExcpMod_logicPhyRegMap_2_valid,rhs_.io_toVecExcpMod_logicPhyRegMap_2_valid),UVM_NONE)
        end

        if(this.io_toVecExcpMod_logicPhyRegMap_2_bits_lreg!=rhs_.io_toVecExcpMod_logicPhyRegMap_2_bits_lreg) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toVecExcpMod_logicPhyRegMap_2_bits_lreg=0x%0h while the rhs_.io_toVecExcpMod_logicPhyRegMap_2_bits_lreg=0x%0h",this.io_toVecExcpMod_logicPhyRegMap_2_bits_lreg,rhs_.io_toVecExcpMod_logicPhyRegMap_2_bits_lreg),UVM_NONE)
        end

        if(this.io_toVecExcpMod_logicPhyRegMap_2_bits_preg!=rhs_.io_toVecExcpMod_logicPhyRegMap_2_bits_preg) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toVecExcpMod_logicPhyRegMap_2_bits_preg=0x%0h while the rhs_.io_toVecExcpMod_logicPhyRegMap_2_bits_preg=0x%0h",this.io_toVecExcpMod_logicPhyRegMap_2_bits_preg,rhs_.io_toVecExcpMod_logicPhyRegMap_2_bits_preg),UVM_NONE)
        end

        if(this.io_toVecExcpMod_logicPhyRegMap_3_valid!=rhs_.io_toVecExcpMod_logicPhyRegMap_3_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toVecExcpMod_logicPhyRegMap_3_valid=0x%0h while the rhs_.io_toVecExcpMod_logicPhyRegMap_3_valid=0x%0h",this.io_toVecExcpMod_logicPhyRegMap_3_valid,rhs_.io_toVecExcpMod_logicPhyRegMap_3_valid),UVM_NONE)
        end

        if(this.io_toVecExcpMod_logicPhyRegMap_3_bits_lreg!=rhs_.io_toVecExcpMod_logicPhyRegMap_3_bits_lreg) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toVecExcpMod_logicPhyRegMap_3_bits_lreg=0x%0h while the rhs_.io_toVecExcpMod_logicPhyRegMap_3_bits_lreg=0x%0h",this.io_toVecExcpMod_logicPhyRegMap_3_bits_lreg,rhs_.io_toVecExcpMod_logicPhyRegMap_3_bits_lreg),UVM_NONE)
        end

        if(this.io_toVecExcpMod_logicPhyRegMap_3_bits_preg!=rhs_.io_toVecExcpMod_logicPhyRegMap_3_bits_preg) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toVecExcpMod_logicPhyRegMap_3_bits_preg=0x%0h while the rhs_.io_toVecExcpMod_logicPhyRegMap_3_bits_preg=0x%0h",this.io_toVecExcpMod_logicPhyRegMap_3_bits_preg,rhs_.io_toVecExcpMod_logicPhyRegMap_3_bits_preg),UVM_NONE)
        end

        if(this.io_toVecExcpMod_logicPhyRegMap_4_valid!=rhs_.io_toVecExcpMod_logicPhyRegMap_4_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toVecExcpMod_logicPhyRegMap_4_valid=0x%0h while the rhs_.io_toVecExcpMod_logicPhyRegMap_4_valid=0x%0h",this.io_toVecExcpMod_logicPhyRegMap_4_valid,rhs_.io_toVecExcpMod_logicPhyRegMap_4_valid),UVM_NONE)
        end

        if(this.io_toVecExcpMod_logicPhyRegMap_4_bits_lreg!=rhs_.io_toVecExcpMod_logicPhyRegMap_4_bits_lreg) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toVecExcpMod_logicPhyRegMap_4_bits_lreg=0x%0h while the rhs_.io_toVecExcpMod_logicPhyRegMap_4_bits_lreg=0x%0h",this.io_toVecExcpMod_logicPhyRegMap_4_bits_lreg,rhs_.io_toVecExcpMod_logicPhyRegMap_4_bits_lreg),UVM_NONE)
        end

        if(this.io_toVecExcpMod_logicPhyRegMap_4_bits_preg!=rhs_.io_toVecExcpMod_logicPhyRegMap_4_bits_preg) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toVecExcpMod_logicPhyRegMap_4_bits_preg=0x%0h while the rhs_.io_toVecExcpMod_logicPhyRegMap_4_bits_preg=0x%0h",this.io_toVecExcpMod_logicPhyRegMap_4_bits_preg,rhs_.io_toVecExcpMod_logicPhyRegMap_4_bits_preg),UVM_NONE)
        end

        if(this.io_toVecExcpMod_logicPhyRegMap_5_valid!=rhs_.io_toVecExcpMod_logicPhyRegMap_5_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toVecExcpMod_logicPhyRegMap_5_valid=0x%0h while the rhs_.io_toVecExcpMod_logicPhyRegMap_5_valid=0x%0h",this.io_toVecExcpMod_logicPhyRegMap_5_valid,rhs_.io_toVecExcpMod_logicPhyRegMap_5_valid),UVM_NONE)
        end

        if(this.io_toVecExcpMod_logicPhyRegMap_5_bits_lreg!=rhs_.io_toVecExcpMod_logicPhyRegMap_5_bits_lreg) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toVecExcpMod_logicPhyRegMap_5_bits_lreg=0x%0h while the rhs_.io_toVecExcpMod_logicPhyRegMap_5_bits_lreg=0x%0h",this.io_toVecExcpMod_logicPhyRegMap_5_bits_lreg,rhs_.io_toVecExcpMod_logicPhyRegMap_5_bits_lreg),UVM_NONE)
        end

        if(this.io_toVecExcpMod_logicPhyRegMap_5_bits_preg!=rhs_.io_toVecExcpMod_logicPhyRegMap_5_bits_preg) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toVecExcpMod_logicPhyRegMap_5_bits_preg=0x%0h while the rhs_.io_toVecExcpMod_logicPhyRegMap_5_bits_preg=0x%0h",this.io_toVecExcpMod_logicPhyRegMap_5_bits_preg,rhs_.io_toVecExcpMod_logicPhyRegMap_5_bits_preg),UVM_NONE)
        end

        if(this.io_toVecExcpMod_excpInfo_valid!=rhs_.io_toVecExcpMod_excpInfo_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toVecExcpMod_excpInfo_valid=0x%0h while the rhs_.io_toVecExcpMod_excpInfo_valid=0x%0h",this.io_toVecExcpMod_excpInfo_valid,rhs_.io_toVecExcpMod_excpInfo_valid),UVM_NONE)
        end

        if(this.io_toVecExcpMod_excpInfo_bits_vstart!=rhs_.io_toVecExcpMod_excpInfo_bits_vstart) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toVecExcpMod_excpInfo_bits_vstart=0x%0h while the rhs_.io_toVecExcpMod_excpInfo_bits_vstart=0x%0h",this.io_toVecExcpMod_excpInfo_bits_vstart,rhs_.io_toVecExcpMod_excpInfo_bits_vstart),UVM_NONE)
        end

        if(this.io_toVecExcpMod_excpInfo_bits_vsew!=rhs_.io_toVecExcpMod_excpInfo_bits_vsew) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toVecExcpMod_excpInfo_bits_vsew=0x%0h while the rhs_.io_toVecExcpMod_excpInfo_bits_vsew=0x%0h",this.io_toVecExcpMod_excpInfo_bits_vsew,rhs_.io_toVecExcpMod_excpInfo_bits_vsew),UVM_NONE)
        end

        if(this.io_toVecExcpMod_excpInfo_bits_veew!=rhs_.io_toVecExcpMod_excpInfo_bits_veew) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toVecExcpMod_excpInfo_bits_veew=0x%0h while the rhs_.io_toVecExcpMod_excpInfo_bits_veew=0x%0h",this.io_toVecExcpMod_excpInfo_bits_veew,rhs_.io_toVecExcpMod_excpInfo_bits_veew),UVM_NONE)
        end

        if(this.io_toVecExcpMod_excpInfo_bits_vlmul!=rhs_.io_toVecExcpMod_excpInfo_bits_vlmul) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toVecExcpMod_excpInfo_bits_vlmul=0x%0h while the rhs_.io_toVecExcpMod_excpInfo_bits_vlmul=0x%0h",this.io_toVecExcpMod_excpInfo_bits_vlmul,rhs_.io_toVecExcpMod_excpInfo_bits_vlmul),UVM_NONE)
        end

        if(this.io_toVecExcpMod_excpInfo_bits_nf!=rhs_.io_toVecExcpMod_excpInfo_bits_nf) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toVecExcpMod_excpInfo_bits_nf=0x%0h while the rhs_.io_toVecExcpMod_excpInfo_bits_nf=0x%0h",this.io_toVecExcpMod_excpInfo_bits_nf,rhs_.io_toVecExcpMod_excpInfo_bits_nf),UVM_NONE)
        end

        if(this.io_toVecExcpMod_excpInfo_bits_isStride!=rhs_.io_toVecExcpMod_excpInfo_bits_isStride) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toVecExcpMod_excpInfo_bits_isStride=0x%0h while the rhs_.io_toVecExcpMod_excpInfo_bits_isStride=0x%0h",this.io_toVecExcpMod_excpInfo_bits_isStride,rhs_.io_toVecExcpMod_excpInfo_bits_isStride),UVM_NONE)
        end

        if(this.io_toVecExcpMod_excpInfo_bits_isIndexed!=rhs_.io_toVecExcpMod_excpInfo_bits_isIndexed) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toVecExcpMod_excpInfo_bits_isIndexed=0x%0h while the rhs_.io_toVecExcpMod_excpInfo_bits_isIndexed=0x%0h",this.io_toVecExcpMod_excpInfo_bits_isIndexed,rhs_.io_toVecExcpMod_excpInfo_bits_isIndexed),UVM_NONE)
        end

        if(this.io_toVecExcpMod_excpInfo_bits_isWhole!=rhs_.io_toVecExcpMod_excpInfo_bits_isWhole) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toVecExcpMod_excpInfo_bits_isWhole=0x%0h while the rhs_.io_toVecExcpMod_excpInfo_bits_isWhole=0x%0h",this.io_toVecExcpMod_excpInfo_bits_isWhole,rhs_.io_toVecExcpMod_excpInfo_bits_isWhole),UVM_NONE)
        end

        if(this.io_toVecExcpMod_excpInfo_bits_isVlm!=rhs_.io_toVecExcpMod_excpInfo_bits_isVlm) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_toVecExcpMod_excpInfo_bits_isVlm=0x%0h while the rhs_.io_toVecExcpMod_excpInfo_bits_isVlm=0x%0h",this.io_toVecExcpMod_excpInfo_bits_isVlm,rhs_.io_toVecExcpMod_excpInfo_bits_isVlm),UVM_NONE)
        end

        if(this.io_storeDebugInfo_1_pc!=rhs_.io_storeDebugInfo_1_pc) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_storeDebugInfo_1_pc=0x%0h while the rhs_.io_storeDebugInfo_1_pc=0x%0h",this.io_storeDebugInfo_1_pc,rhs_.io_storeDebugInfo_1_pc),UVM_NONE)
        end

        if(this.io_perf_0_value!=rhs_.io_perf_0_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_perf_0_value=0x%0h while the rhs_.io_perf_0_value=0x%0h",this.io_perf_0_value,rhs_.io_perf_0_value),UVM_NONE)
        end

        if(this.io_perf_1_value!=rhs_.io_perf_1_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_perf_1_value=0x%0h while the rhs_.io_perf_1_value=0x%0h",this.io_perf_1_value,rhs_.io_perf_1_value),UVM_NONE)
        end

        if(this.io_perf_2_value!=rhs_.io_perf_2_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_perf_2_value=0x%0h while the rhs_.io_perf_2_value=0x%0h",this.io_perf_2_value,rhs_.io_perf_2_value),UVM_NONE)
        end

        if(this.io_perf_3_value!=rhs_.io_perf_3_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_perf_3_value=0x%0h while the rhs_.io_perf_3_value=0x%0h",this.io_perf_3_value,rhs_.io_perf_3_value),UVM_NONE)
        end

        if(this.io_perf_4_value!=rhs_.io_perf_4_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_perf_4_value=0x%0h while the rhs_.io_perf_4_value=0x%0h",this.io_perf_4_value,rhs_.io_perf_4_value),UVM_NONE)
        end

        if(this.io_perf_5_value!=rhs_.io_perf_5_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_perf_5_value=0x%0h while the rhs_.io_perf_5_value=0x%0h",this.io_perf_5_value,rhs_.io_perf_5_value),UVM_NONE)
        end

        if(this.io_perf_6_value!=rhs_.io_perf_6_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_perf_6_value=0x%0h while the rhs_.io_perf_6_value=0x%0h",this.io_perf_6_value,rhs_.io_perf_6_value),UVM_NONE)
        end

        if(this.io_perf_7_value!=rhs_.io_perf_7_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_perf_7_value=0x%0h while the rhs_.io_perf_7_value=0x%0h",this.io_perf_7_value,rhs_.io_perf_7_value),UVM_NONE)
        end

        if(this.io_perf_8_value!=rhs_.io_perf_8_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_perf_8_value=0x%0h while the rhs_.io_perf_8_value=0x%0h",this.io_perf_8_value,rhs_.io_perf_8_value),UVM_NONE)
        end

        if(this.io_perf_9_value!=rhs_.io_perf_9_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_perf_9_value=0x%0h while the rhs_.io_perf_9_value=0x%0h",this.io_perf_9_value,rhs_.io_perf_9_value),UVM_NONE)
        end

        if(this.io_perf_10_value!=rhs_.io_perf_10_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_perf_10_value=0x%0h while the rhs_.io_perf_10_value=0x%0h",this.io_perf_10_value,rhs_.io_perf_10_value),UVM_NONE)
        end

        if(this.io_perf_11_value!=rhs_.io_perf_11_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_perf_11_value=0x%0h while the rhs_.io_perf_11_value=0x%0h",this.io_perf_11_value,rhs_.io_perf_11_value),UVM_NONE)
        end

        if(this.io_perf_12_value!=rhs_.io_perf_12_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_perf_12_value=0x%0h while the rhs_.io_perf_12_value=0x%0h",this.io_perf_12_value,rhs_.io_perf_12_value),UVM_NONE)
        end

        if(this.io_perf_13_value!=rhs_.io_perf_13_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_perf_13_value=0x%0h while the rhs_.io_perf_13_value=0x%0h",this.io_perf_13_value,rhs_.io_perf_13_value),UVM_NONE)
        end

        if(this.io_perf_14_value!=rhs_.io_perf_14_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_perf_14_value=0x%0h while the rhs_.io_perf_14_value=0x%0h",this.io_perf_14_value,rhs_.io_perf_14_value),UVM_NONE)
        end

        if(this.io_perf_15_value!=rhs_.io_perf_15_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_perf_15_value=0x%0h while the rhs_.io_perf_15_value=0x%0h",this.io_perf_15_value,rhs_.io_perf_15_value),UVM_NONE)
        end

        if(this.io_perf_16_value!=rhs_.io_perf_16_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_perf_16_value=0x%0h while the rhs_.io_perf_16_value=0x%0h",this.io_perf_16_value,rhs_.io_perf_16_value),UVM_NONE)
        end

        if(this.io_perf_17_value!=rhs_.io_perf_17_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_perf_17_value=0x%0h while the rhs_.io_perf_17_value=0x%0h",this.io_perf_17_value,rhs_.io_perf_17_value),UVM_NONE)
        end

        if(this.io_error_0!=rhs_.io_error_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_error_0=0x%0h while the rhs_.io_error_0=0x%0h",this.io_error_0,rhs_.io_error_0),UVM_NONE)
        end

    end
    return super_result;
endfunction:compare

`endif


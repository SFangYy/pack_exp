//=========================================================
//File name    : Redirect_in_agent_dec.sv
//Author       : nanyunhao
//Module name  : Redirect_in_agent_dec
//Discribution : Redirect_in_agent_dec : parameter
//Date         : 2026-01-22
//=========================================================
`ifndef REDIRECT_IN_AGENT_DEC__SV
`define REDIRECT_IN_AGENT_DEC__SV

package Redirect_in_agent_dec;

endpackage:Redirect_in_agent_dec

import Redirect_in_agent_dec::*;

`endif


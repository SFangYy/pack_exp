//=========================================================
//File name    : WriteBack_in_agent_interface.sv
//Author       : nanyunhao
//Module name  : WriteBack_in_agent_interface
//Discribution : WriteBack_in_agent_interface : signal interface
//Date         : 2026-01-22
//=========================================================
`ifndef WRITEBACK_IN_AGENT_INTERFACE__SV
`define WRITEBACK_IN_AGENT_INTERFACE__SV

`ifndef DEF_SETUP_TIME
    `define DEF_SETUP_TIME 1
`endif
`ifndef DEF_HOLD_TIME
    `define DEF_HOLD_TIME 1
`endif

interface WriteBack_in_agent_interface  (input bit clk,input bit rst_n);

    logic         io_writeback_24_valid;
    logic [127:0] io_writeback_24_bits_data_0;
    logic [6:0]   io_writeback_24_bits_pdest;
    logic         io_writeback_24_bits_robIdx_flag;
    logic [7:0]   io_writeback_24_bits_robIdx_value;
    logic         io_writeback_24_bits_vecWen;
    logic         io_writeback_24_bits_v0Wen;
    logic         io_writeback_24_bits_vlWen;
    logic         io_writeback_24_bits_exceptionVec_0;
    logic         io_writeback_24_bits_exceptionVec_1;
    logic         io_writeback_24_bits_exceptionVec_2;
    logic         io_writeback_24_bits_exceptionVec_3;
    logic         io_writeback_24_bits_exceptionVec_4;
    logic         io_writeback_24_bits_exceptionVec_5;
    logic         io_writeback_24_bits_exceptionVec_6;
    logic         io_writeback_24_bits_exceptionVec_7;
    logic         io_writeback_24_bits_exceptionVec_8;
    logic         io_writeback_24_bits_exceptionVec_9;
    logic         io_writeback_24_bits_exceptionVec_10;
    logic         io_writeback_24_bits_exceptionVec_11;
    logic         io_writeback_24_bits_exceptionVec_12;
    logic         io_writeback_24_bits_exceptionVec_13;
    logic         io_writeback_24_bits_exceptionVec_14;
    logic         io_writeback_24_bits_exceptionVec_15;
    logic         io_writeback_24_bits_exceptionVec_16;
    logic         io_writeback_24_bits_exceptionVec_17;
    logic         io_writeback_24_bits_exceptionVec_18;
    logic         io_writeback_24_bits_exceptionVec_19;
    logic         io_writeback_24_bits_exceptionVec_20;
    logic         io_writeback_24_bits_exceptionVec_21;
    logic         io_writeback_24_bits_exceptionVec_22;
    logic         io_writeback_24_bits_exceptionVec_23;
    logic         io_writeback_24_bits_flushPipe;
    logic         io_writeback_24_bits_replay;
    logic [3:0]   io_writeback_24_bits_trigger;
    logic         io_writeback_24_bits_vls_vpu_vill;
    logic         io_writeback_24_bits_vls_vpu_vma;
    logic         io_writeback_24_bits_vls_vpu_vta;
    logic [1:0]   io_writeback_24_bits_vls_vpu_vsew;
    logic [2:0]   io_writeback_24_bits_vls_vpu_vlmul;
    logic         io_writeback_24_bits_vls_vpu_specVill;
    logic         io_writeback_24_bits_vls_vpu_specVma;
    logic         io_writeback_24_bits_vls_vpu_specVta;
    logic [1:0]   io_writeback_24_bits_vls_vpu_specVsew;
    logic [2:0]   io_writeback_24_bits_vls_vpu_specVlmul;
    logic         io_writeback_24_bits_vls_vpu_vm;
    logic [7:0]   io_writeback_24_bits_vls_vpu_vstart;
    logic [2:0]   io_writeback_24_bits_vls_vpu_frm;
    logic         io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst;
    logic         io_writeback_24_bits_vls_vpu_fpu_isFP32Instr;
    logic         io_writeback_24_bits_vls_vpu_fpu_isFP64Instr;
    logic         io_writeback_24_bits_vls_vpu_fpu_isReduction;
    logic         io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2;
    logic         io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4;
    logic         io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8;
    logic [1:0]   io_writeback_24_bits_vls_vpu_vxrm;
    logic [6:0]   io_writeback_24_bits_vls_vpu_vuopIdx;
    logic         io_writeback_24_bits_vls_vpu_lastUop;
    logic [127:0] io_writeback_24_bits_vls_vpu_vmask;
    logic [7:0]   io_writeback_24_bits_vls_vpu_vl;
    logic [2:0]   io_writeback_24_bits_vls_vpu_nf;
    logic [1:0]   io_writeback_24_bits_vls_vpu_veew;
    logic         io_writeback_24_bits_vls_vpu_isReverse;
    logic         io_writeback_24_bits_vls_vpu_isExt;
    logic         io_writeback_24_bits_vls_vpu_isNarrow;
    logic         io_writeback_24_bits_vls_vpu_isDstMask;
    logic         io_writeback_24_bits_vls_vpu_isOpMask;
    logic         io_writeback_24_bits_vls_vpu_isMove;
    logic         io_writeback_24_bits_vls_vpu_isDependOldVd;
    logic         io_writeback_24_bits_vls_vpu_isWritePartVd;
    logic         io_writeback_24_bits_vls_vpu_isVleff;
    logic [7:0]   io_writeback_24_bits_vls_oldVdPsrc;
    logic [2:0]   io_writeback_24_bits_vls_vdIdx;
    logic [2:0]   io_writeback_24_bits_vls_vdIdxInField;
    logic         io_writeback_24_bits_vls_isIndexed;
    logic         io_writeback_24_bits_vls_isMasked;
    logic         io_writeback_24_bits_vls_isStrided;
    logic         io_writeback_24_bits_vls_isWhole;
    logic         io_writeback_24_bits_vls_isVecLoad;
    logic         io_writeback_24_bits_vls_isVlm;
    logic         io_writeback_24_bits_debug_isMMIO;
    logic         io_writeback_24_bits_debug_isNCIO;
    logic         io_writeback_24_bits_debug_isPerfCnt;
    logic [47:0]  io_writeback_24_bits_debug_paddr;
    logic [49:0]  io_writeback_24_bits_debug_vaddr;
    logic         io_writeback_24_bits_debugInfo_eliminatedMove;
    logic [63:0]  io_writeback_24_bits_debugInfo_renameTime;
    logic [63:0]  io_writeback_24_bits_debugInfo_dispatchTime;
    logic [63:0]  io_writeback_24_bits_debugInfo_enqRsTime;
    logic [63:0]  io_writeback_24_bits_debugInfo_selectTime;
    logic [63:0]  io_writeback_24_bits_debugInfo_issueTime;
    logic [63:0]  io_writeback_24_bits_debugInfo_writebackTime;
    logic [63:0]  io_writeback_24_bits_debugInfo_runahead_checkpoint_id;
    logic [63:0]  io_writeback_24_bits_debugInfo_tlbFirstReqTime;
    logic [63:0]  io_writeback_24_bits_debugInfo_tlbRespTime;
    logic [63:0]  io_writeback_24_bits_debug_seqNum;
    logic         io_writeback_23_valid;
    logic [127:0] io_writeback_23_bits_data_0;
    logic [6:0]   io_writeback_23_bits_pdest;
    logic         io_writeback_23_bits_robIdx_flag;
    logic [7:0]   io_writeback_23_bits_robIdx_value;
    logic         io_writeback_23_bits_vecWen;
    logic         io_writeback_23_bits_v0Wen;
    logic         io_writeback_23_bits_vlWen;
    logic         io_writeback_23_bits_exceptionVec_0;
    logic         io_writeback_23_bits_exceptionVec_1;
    logic         io_writeback_23_bits_exceptionVec_2;
    logic         io_writeback_23_bits_exceptionVec_3;
    logic         io_writeback_23_bits_exceptionVec_4;
    logic         io_writeback_23_bits_exceptionVec_5;
    logic         io_writeback_23_bits_exceptionVec_6;
    logic         io_writeback_23_bits_exceptionVec_7;
    logic         io_writeback_23_bits_exceptionVec_8;
    logic         io_writeback_23_bits_exceptionVec_9;
    logic         io_writeback_23_bits_exceptionVec_10;
    logic         io_writeback_23_bits_exceptionVec_11;
    logic         io_writeback_23_bits_exceptionVec_12;
    logic         io_writeback_23_bits_exceptionVec_13;
    logic         io_writeback_23_bits_exceptionVec_14;
    logic         io_writeback_23_bits_exceptionVec_15;
    logic         io_writeback_23_bits_exceptionVec_16;
    logic         io_writeback_23_bits_exceptionVec_17;
    logic         io_writeback_23_bits_exceptionVec_18;
    logic         io_writeback_23_bits_exceptionVec_19;
    logic         io_writeback_23_bits_exceptionVec_20;
    logic         io_writeback_23_bits_exceptionVec_21;
    logic         io_writeback_23_bits_exceptionVec_22;
    logic         io_writeback_23_bits_exceptionVec_23;
    logic         io_writeback_23_bits_flushPipe;
    logic         io_writeback_23_bits_replay;
    logic [3:0]   io_writeback_23_bits_trigger;
    logic         io_writeback_23_bits_vls_vpu_vill;
    logic         io_writeback_23_bits_vls_vpu_vma;
    logic         io_writeback_23_bits_vls_vpu_vta;
    logic [1:0]   io_writeback_23_bits_vls_vpu_vsew;
    logic [2:0]   io_writeback_23_bits_vls_vpu_vlmul;
    logic         io_writeback_23_bits_vls_vpu_specVill;
    logic         io_writeback_23_bits_vls_vpu_specVma;
    logic         io_writeback_23_bits_vls_vpu_specVta;
    logic [1:0]   io_writeback_23_bits_vls_vpu_specVsew;
    logic [2:0]   io_writeback_23_bits_vls_vpu_specVlmul;
    logic         io_writeback_23_bits_vls_vpu_vm;
    logic [7:0]   io_writeback_23_bits_vls_vpu_vstart;
    logic [2:0]   io_writeback_23_bits_vls_vpu_frm;
    logic         io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst;
    logic         io_writeback_23_bits_vls_vpu_fpu_isFP32Instr;
    logic         io_writeback_23_bits_vls_vpu_fpu_isFP64Instr;
    logic         io_writeback_23_bits_vls_vpu_fpu_isReduction;
    logic         io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2;
    logic         io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4;
    logic         io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8;
    logic [1:0]   io_writeback_23_bits_vls_vpu_vxrm;
    logic [6:0]   io_writeback_23_bits_vls_vpu_vuopIdx;
    logic         io_writeback_23_bits_vls_vpu_lastUop;
    logic [127:0] io_writeback_23_bits_vls_vpu_vmask;
    logic [7:0]   io_writeback_23_bits_vls_vpu_vl;
    logic [2:0]   io_writeback_23_bits_vls_vpu_nf;
    logic [1:0]   io_writeback_23_bits_vls_vpu_veew;
    logic         io_writeback_23_bits_vls_vpu_isReverse;
    logic         io_writeback_23_bits_vls_vpu_isExt;
    logic         io_writeback_23_bits_vls_vpu_isNarrow;
    logic         io_writeback_23_bits_vls_vpu_isDstMask;
    logic         io_writeback_23_bits_vls_vpu_isOpMask;
    logic         io_writeback_23_bits_vls_vpu_isMove;
    logic         io_writeback_23_bits_vls_vpu_isDependOldVd;
    logic         io_writeback_23_bits_vls_vpu_isWritePartVd;
    logic         io_writeback_23_bits_vls_vpu_isVleff;
    logic [7:0]   io_writeback_23_bits_vls_oldVdPsrc;
    logic [2:0]   io_writeback_23_bits_vls_vdIdx;
    logic [2:0]   io_writeback_23_bits_vls_vdIdxInField;
    logic         io_writeback_23_bits_vls_isIndexed;
    logic         io_writeback_23_bits_vls_isMasked;
    logic         io_writeback_23_bits_vls_isStrided;
    logic         io_writeback_23_bits_vls_isWhole;
    logic         io_writeback_23_bits_vls_isVecLoad;
    logic         io_writeback_23_bits_vls_isVlm;
    logic         io_writeback_23_bits_debug_isMMIO;
    logic         io_writeback_23_bits_debug_isNCIO;
    logic         io_writeback_23_bits_debug_isPerfCnt;
    logic [47:0]  io_writeback_23_bits_debug_paddr;
    logic [49:0]  io_writeback_23_bits_debug_vaddr;
    logic         io_writeback_23_bits_debugInfo_eliminatedMove;
    logic [63:0]  io_writeback_23_bits_debugInfo_renameTime;
    logic [63:0]  io_writeback_23_bits_debugInfo_dispatchTime;
    logic [63:0]  io_writeback_23_bits_debugInfo_enqRsTime;
    logic [63:0]  io_writeback_23_bits_debugInfo_selectTime;
    logic [63:0]  io_writeback_23_bits_debugInfo_issueTime;
    logic [63:0]  io_writeback_23_bits_debugInfo_writebackTime;
    logic [63:0]  io_writeback_23_bits_debugInfo_runahead_checkpoint_id;
    logic [63:0]  io_writeback_23_bits_debugInfo_tlbFirstReqTime;
    logic [63:0]  io_writeback_23_bits_debugInfo_tlbRespTime;
    logic [63:0]  io_writeback_23_bits_debug_seqNum;
    logic         io_writeback_22_valid;
    logic [63:0]  io_writeback_22_bits_data_0;
    logic [7:0]   io_writeback_22_bits_pdest;
    logic         io_writeback_22_bits_robIdx_flag;
    logic [7:0]   io_writeback_22_bits_robIdx_value;
    logic         io_writeback_22_bits_intWen;
    logic         io_writeback_22_bits_fpWen;
    logic         io_writeback_22_bits_exceptionVec_0;
    logic         io_writeback_22_bits_exceptionVec_1;
    logic         io_writeback_22_bits_exceptionVec_2;
    logic         io_writeback_22_bits_exceptionVec_3;
    logic         io_writeback_22_bits_exceptionVec_4;
    logic         io_writeback_22_bits_exceptionVec_5;
    logic         io_writeback_22_bits_exceptionVec_6;
    logic         io_writeback_22_bits_exceptionVec_7;
    logic         io_writeback_22_bits_exceptionVec_8;
    logic         io_writeback_22_bits_exceptionVec_9;
    logic         io_writeback_22_bits_exceptionVec_10;
    logic         io_writeback_22_bits_exceptionVec_11;
    logic         io_writeback_22_bits_exceptionVec_12;
    logic         io_writeback_22_bits_exceptionVec_13;
    logic         io_writeback_22_bits_exceptionVec_14;
    logic         io_writeback_22_bits_exceptionVec_15;
    logic         io_writeback_22_bits_exceptionVec_16;
    logic         io_writeback_22_bits_exceptionVec_17;
    logic         io_writeback_22_bits_exceptionVec_18;
    logic         io_writeback_22_bits_exceptionVec_19;
    logic         io_writeback_22_bits_exceptionVec_20;
    logic         io_writeback_22_bits_exceptionVec_21;
    logic         io_writeback_22_bits_exceptionVec_22;
    logic         io_writeback_22_bits_exceptionVec_23;
    logic         io_writeback_22_bits_flushPipe;
    logic         io_writeback_22_bits_replay;
    logic         io_writeback_22_bits_lqIdx_flag;
    logic [6:0]   io_writeback_22_bits_lqIdx_value;
    logic [3:0]   io_writeback_22_bits_trigger;
    logic         io_writeback_22_bits_predecodeInfo_valid;
    logic         io_writeback_22_bits_predecodeInfo_isRVC;
    logic [1:0]   io_writeback_22_bits_predecodeInfo_brType;
    logic         io_writeback_22_bits_predecodeInfo_isCall;
    logic         io_writeback_22_bits_predecodeInfo_isRet;
    logic         io_writeback_22_bits_debug_isMMIO;
    logic         io_writeback_22_bits_debug_isNCIO;
    logic         io_writeback_22_bits_debug_isPerfCnt;
    logic [47:0]  io_writeback_22_bits_debug_paddr;
    logic [49:0]  io_writeback_22_bits_debug_vaddr;
    logic         io_writeback_22_bits_debugInfo_eliminatedMove;
    logic [63:0]  io_writeback_22_bits_debugInfo_renameTime;
    logic [63:0]  io_writeback_22_bits_debugInfo_dispatchTime;
    logic [63:0]  io_writeback_22_bits_debugInfo_enqRsTime;
    logic [63:0]  io_writeback_22_bits_debugInfo_selectTime;
    logic [63:0]  io_writeback_22_bits_debugInfo_issueTime;
    logic [63:0]  io_writeback_22_bits_debugInfo_writebackTime;
    logic [63:0]  io_writeback_22_bits_debugInfo_runahead_checkpoint_id;
    logic [63:0]  io_writeback_22_bits_debugInfo_tlbFirstReqTime;
    logic [63:0]  io_writeback_22_bits_debugInfo_tlbRespTime;
    logic [63:0]  io_writeback_22_bits_debug_seqNum;
    logic         io_writeback_21_valid;
    logic [63:0]  io_writeback_21_bits_data_0;
    logic [7:0]   io_writeback_21_bits_pdest;
    logic         io_writeback_21_bits_robIdx_flag;
    logic [7:0]   io_writeback_21_bits_robIdx_value;
    logic         io_writeback_21_bits_intWen;
    logic         io_writeback_21_bits_fpWen;
    logic         io_writeback_21_bits_exceptionVec_0;
    logic         io_writeback_21_bits_exceptionVec_1;
    logic         io_writeback_21_bits_exceptionVec_2;
    logic         io_writeback_21_bits_exceptionVec_3;
    logic         io_writeback_21_bits_exceptionVec_4;
    logic         io_writeback_21_bits_exceptionVec_5;
    logic         io_writeback_21_bits_exceptionVec_6;
    logic         io_writeback_21_bits_exceptionVec_7;
    logic         io_writeback_21_bits_exceptionVec_8;
    logic         io_writeback_21_bits_exceptionVec_9;
    logic         io_writeback_21_bits_exceptionVec_10;
    logic         io_writeback_21_bits_exceptionVec_11;
    logic         io_writeback_21_bits_exceptionVec_12;
    logic         io_writeback_21_bits_exceptionVec_13;
    logic         io_writeback_21_bits_exceptionVec_14;
    logic         io_writeback_21_bits_exceptionVec_15;
    logic         io_writeback_21_bits_exceptionVec_16;
    logic         io_writeback_21_bits_exceptionVec_17;
    logic         io_writeback_21_bits_exceptionVec_18;
    logic         io_writeback_21_bits_exceptionVec_19;
    logic         io_writeback_21_bits_exceptionVec_20;
    logic         io_writeback_21_bits_exceptionVec_21;
    logic         io_writeback_21_bits_exceptionVec_22;
    logic         io_writeback_21_bits_exceptionVec_23;
    logic         io_writeback_21_bits_flushPipe;
    logic         io_writeback_21_bits_replay;
    logic         io_writeback_21_bits_lqIdx_flag;
    logic [6:0]   io_writeback_21_bits_lqIdx_value;
    logic [3:0]   io_writeback_21_bits_trigger;
    logic         io_writeback_21_bits_predecodeInfo_valid;
    logic         io_writeback_21_bits_predecodeInfo_isRVC;
    logic [1:0]   io_writeback_21_bits_predecodeInfo_brType;
    logic         io_writeback_21_bits_predecodeInfo_isCall;
    logic         io_writeback_21_bits_predecodeInfo_isRet;
    logic         io_writeback_21_bits_debug_isMMIO;
    logic         io_writeback_21_bits_debug_isNCIO;
    logic         io_writeback_21_bits_debug_isPerfCnt;
    logic [47:0]  io_writeback_21_bits_debug_paddr;
    logic [49:0]  io_writeback_21_bits_debug_vaddr;
    logic         io_writeback_21_bits_debugInfo_eliminatedMove;
    logic [63:0]  io_writeback_21_bits_debugInfo_renameTime;
    logic [63:0]  io_writeback_21_bits_debugInfo_dispatchTime;
    logic [63:0]  io_writeback_21_bits_debugInfo_enqRsTime;
    logic [63:0]  io_writeback_21_bits_debugInfo_selectTime;
    logic [63:0]  io_writeback_21_bits_debugInfo_issueTime;
    logic [63:0]  io_writeback_21_bits_debugInfo_writebackTime;
    logic [63:0]  io_writeback_21_bits_debugInfo_runahead_checkpoint_id;
    logic [63:0]  io_writeback_21_bits_debugInfo_tlbFirstReqTime;
    logic [63:0]  io_writeback_21_bits_debugInfo_tlbRespTime;
    logic [63:0]  io_writeback_21_bits_debug_seqNum;
    logic         io_writeback_20_valid;
    logic [63:0]  io_writeback_20_bits_data_0;
    logic [7:0]   io_writeback_20_bits_pdest;
    logic         io_writeback_20_bits_robIdx_flag;
    logic [7:0]   io_writeback_20_bits_robIdx_value;
    logic         io_writeback_20_bits_intWen;
    logic         io_writeback_20_bits_fpWen;
    logic         io_writeback_20_bits_exceptionVec_0;
    logic         io_writeback_20_bits_exceptionVec_1;
    logic         io_writeback_20_bits_exceptionVec_2;
    logic         io_writeback_20_bits_exceptionVec_3;
    logic         io_writeback_20_bits_exceptionVec_4;
    logic         io_writeback_20_bits_exceptionVec_5;
    logic         io_writeback_20_bits_exceptionVec_6;
    logic         io_writeback_20_bits_exceptionVec_7;
    logic         io_writeback_20_bits_exceptionVec_8;
    logic         io_writeback_20_bits_exceptionVec_9;
    logic         io_writeback_20_bits_exceptionVec_10;
    logic         io_writeback_20_bits_exceptionVec_11;
    logic         io_writeback_20_bits_exceptionVec_12;
    logic         io_writeback_20_bits_exceptionVec_13;
    logic         io_writeback_20_bits_exceptionVec_14;
    logic         io_writeback_20_bits_exceptionVec_15;
    logic         io_writeback_20_bits_exceptionVec_16;
    logic         io_writeback_20_bits_exceptionVec_17;
    logic         io_writeback_20_bits_exceptionVec_18;
    logic         io_writeback_20_bits_exceptionVec_19;
    logic         io_writeback_20_bits_exceptionVec_20;
    logic         io_writeback_20_bits_exceptionVec_21;
    logic         io_writeback_20_bits_exceptionVec_22;
    logic         io_writeback_20_bits_exceptionVec_23;
    logic         io_writeback_20_bits_flushPipe;
    logic         io_writeback_20_bits_replay;
    logic         io_writeback_20_bits_lqIdx_flag;
    logic [6:0]   io_writeback_20_bits_lqIdx_value;
    logic [3:0]   io_writeback_20_bits_trigger;
    logic         io_writeback_20_bits_predecodeInfo_valid;
    logic         io_writeback_20_bits_predecodeInfo_isRVC;
    logic [1:0]   io_writeback_20_bits_predecodeInfo_brType;
    logic         io_writeback_20_bits_predecodeInfo_isCall;
    logic         io_writeback_20_bits_predecodeInfo_isRet;
    logic         io_writeback_20_bits_debug_isMMIO;
    logic         io_writeback_20_bits_debug_isNCIO;
    logic         io_writeback_20_bits_debug_isPerfCnt;
    logic [47:0]  io_writeback_20_bits_debug_paddr;
    logic [49:0]  io_writeback_20_bits_debug_vaddr;
    logic         io_writeback_20_bits_debugInfo_eliminatedMove;
    logic [63:0]  io_writeback_20_bits_debugInfo_renameTime;
    logic [63:0]  io_writeback_20_bits_debugInfo_dispatchTime;
    logic [63:0]  io_writeback_20_bits_debugInfo_enqRsTime;
    logic [63:0]  io_writeback_20_bits_debugInfo_selectTime;
    logic [63:0]  io_writeback_20_bits_debugInfo_issueTime;
    logic [63:0]  io_writeback_20_bits_debugInfo_writebackTime;
    logic [63:0]  io_writeback_20_bits_debugInfo_runahead_checkpoint_id;
    logic [63:0]  io_writeback_20_bits_debugInfo_tlbFirstReqTime;
    logic [63:0]  io_writeback_20_bits_debugInfo_tlbRespTime;
    logic [63:0]  io_writeback_20_bits_debug_seqNum;
    logic         io_writeback_19_valid;
    logic [63:0]  io_writeback_19_bits_data_0;
    logic [7:0]   io_writeback_19_bits_pdest;
    logic         io_writeback_19_bits_robIdx_flag;
    logic [7:0]   io_writeback_19_bits_robIdx_value;
    logic         io_writeback_19_bits_intWen;
    logic         io_writeback_19_bits_exceptionVec_0;
    logic         io_writeback_19_bits_exceptionVec_1;
    logic         io_writeback_19_bits_exceptionVec_2;
    logic         io_writeback_19_bits_exceptionVec_3;
    logic         io_writeback_19_bits_exceptionVec_4;
    logic         io_writeback_19_bits_exceptionVec_5;
    logic         io_writeback_19_bits_exceptionVec_6;
    logic         io_writeback_19_bits_exceptionVec_7;
    logic         io_writeback_19_bits_exceptionVec_8;
    logic         io_writeback_19_bits_exceptionVec_9;
    logic         io_writeback_19_bits_exceptionVec_10;
    logic         io_writeback_19_bits_exceptionVec_11;
    logic         io_writeback_19_bits_exceptionVec_12;
    logic         io_writeback_19_bits_exceptionVec_13;
    logic         io_writeback_19_bits_exceptionVec_14;
    logic         io_writeback_19_bits_exceptionVec_15;
    logic         io_writeback_19_bits_exceptionVec_16;
    logic         io_writeback_19_bits_exceptionVec_17;
    logic         io_writeback_19_bits_exceptionVec_18;
    logic         io_writeback_19_bits_exceptionVec_19;
    logic         io_writeback_19_bits_exceptionVec_20;
    logic         io_writeback_19_bits_exceptionVec_21;
    logic         io_writeback_19_bits_exceptionVec_22;
    logic         io_writeback_19_bits_exceptionVec_23;
    logic         io_writeback_19_bits_flushPipe;
    logic         io_writeback_19_bits_sqIdx_flag;
    logic [5:0]   io_writeback_19_bits_sqIdx_value;
    logic [3:0]   io_writeback_19_bits_trigger;
    logic         io_writeback_19_bits_debug_isMMIO;
    logic         io_writeback_19_bits_debug_isNCIO;
    logic         io_writeback_19_bits_debug_isPerfCnt;
    logic [47:0]  io_writeback_19_bits_debug_paddr;
    logic [49:0]  io_writeback_19_bits_debug_vaddr;
    logic         io_writeback_19_bits_debugInfo_eliminatedMove;
    logic [63:0]  io_writeback_19_bits_debugInfo_renameTime;
    logic [63:0]  io_writeback_19_bits_debugInfo_dispatchTime;
    logic [63:0]  io_writeback_19_bits_debugInfo_enqRsTime;
    logic [63:0]  io_writeback_19_bits_debugInfo_selectTime;
    logic [63:0]  io_writeback_19_bits_debugInfo_issueTime;
    logic [63:0]  io_writeback_19_bits_debugInfo_writebackTime;
    logic [63:0]  io_writeback_19_bits_debugInfo_runahead_checkpoint_id;
    logic [63:0]  io_writeback_19_bits_debugInfo_tlbFirstReqTime;
    logic [63:0]  io_writeback_19_bits_debugInfo_tlbRespTime;
    logic [63:0]  io_writeback_19_bits_debug_seqNum;
    logic         io_writeback_18_valid;
    logic [63:0]  io_writeback_18_bits_data_0;
    logic [7:0]   io_writeback_18_bits_pdest;
    logic         io_writeback_18_bits_robIdx_flag;
    logic [7:0]   io_writeback_18_bits_robIdx_value;
    logic         io_writeback_18_bits_intWen;
    logic         io_writeback_18_bits_exceptionVec_0;
    logic         io_writeback_18_bits_exceptionVec_1;
    logic         io_writeback_18_bits_exceptionVec_2;
    logic         io_writeback_18_bits_exceptionVec_3;
    logic         io_writeback_18_bits_exceptionVec_4;
    logic         io_writeback_18_bits_exceptionVec_5;
    logic         io_writeback_18_bits_exceptionVec_6;
    logic         io_writeback_18_bits_exceptionVec_7;
    logic         io_writeback_18_bits_exceptionVec_8;
    logic         io_writeback_18_bits_exceptionVec_9;
    logic         io_writeback_18_bits_exceptionVec_10;
    logic         io_writeback_18_bits_exceptionVec_11;
    logic         io_writeback_18_bits_exceptionVec_12;
    logic         io_writeback_18_bits_exceptionVec_13;
    logic         io_writeback_18_bits_exceptionVec_14;
    logic         io_writeback_18_bits_exceptionVec_15;
    logic         io_writeback_18_bits_exceptionVec_16;
    logic         io_writeback_18_bits_exceptionVec_17;
    logic         io_writeback_18_bits_exceptionVec_18;
    logic         io_writeback_18_bits_exceptionVec_19;
    logic         io_writeback_18_bits_exceptionVec_20;
    logic         io_writeback_18_bits_exceptionVec_21;
    logic         io_writeback_18_bits_exceptionVec_22;
    logic         io_writeback_18_bits_exceptionVec_23;
    logic         io_writeback_18_bits_flushPipe;
    logic         io_writeback_18_bits_sqIdx_flag;
    logic [5:0]   io_writeback_18_bits_sqIdx_value;
    logic [3:0]   io_writeback_18_bits_trigger;
    logic         io_writeback_18_bits_debug_isMMIO;
    logic         io_writeback_18_bits_debug_isNCIO;
    logic         io_writeback_18_bits_debug_isPerfCnt;
    logic [47:0]  io_writeback_18_bits_debug_paddr;
    logic [49:0]  io_writeback_18_bits_debug_vaddr;
    logic         io_writeback_18_bits_debugInfo_eliminatedMove;
    logic [63:0]  io_writeback_18_bits_debugInfo_renameTime;
    logic [63:0]  io_writeback_18_bits_debugInfo_dispatchTime;
    logic [63:0]  io_writeback_18_bits_debugInfo_enqRsTime;
    logic [63:0]  io_writeback_18_bits_debugInfo_selectTime;
    logic [63:0]  io_writeback_18_bits_debugInfo_issueTime;
    logic [63:0]  io_writeback_18_bits_debugInfo_writebackTime;
    logic [63:0]  io_writeback_18_bits_debugInfo_runahead_checkpoint_id;
    logic [63:0]  io_writeback_18_bits_debugInfo_tlbFirstReqTime;
    logic [63:0]  io_writeback_18_bits_debugInfo_tlbRespTime;
    logic [63:0]  io_writeback_18_bits_debug_seqNum;
    logic         io_writeback_17_valid;
    logic [127:0] io_writeback_17_bits_data_0;
    logic [127:0] io_writeback_17_bits_data_1;
    logic [127:0] io_writeback_17_bits_data_2;
    logic [6:0]   io_writeback_17_bits_pdest;
    logic         io_writeback_17_bits_robIdx_flag;
    logic [7:0]   io_writeback_17_bits_robIdx_value;
    logic         io_writeback_17_bits_vecWen;
    logic         io_writeback_17_bits_v0Wen;
    logic [4:0]   io_writeback_17_bits_fflags;
    logic         io_writeback_17_bits_wflags;
    logic         io_writeback_17_bits_debugInfo_eliminatedMove;
    logic [63:0]  io_writeback_17_bits_debugInfo_renameTime;
    logic [63:0]  io_writeback_17_bits_debugInfo_dispatchTime;
    logic [63:0]  io_writeback_17_bits_debugInfo_enqRsTime;
    logic [63:0]  io_writeback_17_bits_debugInfo_selectTime;
    logic [63:0]  io_writeback_17_bits_debugInfo_issueTime;
    logic [63:0]  io_writeback_17_bits_debugInfo_writebackTime;
    logic [63:0]  io_writeback_17_bits_debugInfo_runahead_checkpoint_id;
    logic [63:0]  io_writeback_17_bits_debugInfo_tlbFirstReqTime;
    logic [63:0]  io_writeback_17_bits_debugInfo_tlbRespTime;
    logic [63:0]  io_writeback_17_bits_debug_seqNum;
    logic         io_writeback_16_valid;
    logic [127:0] io_writeback_16_bits_data_0;
    logic [127:0] io_writeback_16_bits_data_1;
    logic [127:0] io_writeback_16_bits_data_2;
    logic [127:0] io_writeback_16_bits_data_3;
    logic [7:0]   io_writeback_16_bits_pdest;
    logic         io_writeback_16_bits_robIdx_flag;
    logic [7:0]   io_writeback_16_bits_robIdx_value;
    logic         io_writeback_16_bits_fpWen;
    logic         io_writeback_16_bits_vecWen;
    logic         io_writeback_16_bits_v0Wen;
    logic [4:0]   io_writeback_16_bits_fflags;
    logic         io_writeback_16_bits_wflags;
    logic         io_writeback_16_bits_debugInfo_eliminatedMove;
    logic [63:0]  io_writeback_16_bits_debugInfo_renameTime;
    logic [63:0]  io_writeback_16_bits_debugInfo_dispatchTime;
    logic [63:0]  io_writeback_16_bits_debugInfo_enqRsTime;
    logic [63:0]  io_writeback_16_bits_debugInfo_selectTime;
    logic [63:0]  io_writeback_16_bits_debugInfo_issueTime;
    logic [63:0]  io_writeback_16_bits_debugInfo_writebackTime;
    logic [63:0]  io_writeback_16_bits_debugInfo_runahead_checkpoint_id;
    logic [63:0]  io_writeback_16_bits_debugInfo_tlbFirstReqTime;
    logic [63:0]  io_writeback_16_bits_debugInfo_tlbRespTime;
    logic [63:0]  io_writeback_16_bits_debug_seqNum;
    logic         io_writeback_15_valid;
    logic [127:0] io_writeback_15_bits_data_0;
    logic [127:0] io_writeback_15_bits_data_1;
    logic [127:0] io_writeback_15_bits_data_2;
    logic [6:0]   io_writeback_15_bits_pdest;
    logic         io_writeback_15_bits_robIdx_flag;
    logic [7:0]   io_writeback_15_bits_robIdx_value;
    logic         io_writeback_15_bits_vecWen;
    logic         io_writeback_15_bits_v0Wen;
    logic [4:0]   io_writeback_15_bits_fflags;
    logic         io_writeback_15_bits_wflags;
    logic         io_writeback_15_bits_vxsat;
    logic         io_writeback_15_bits_debugInfo_eliminatedMove;
    logic [63:0]  io_writeback_15_bits_debugInfo_renameTime;
    logic [63:0]  io_writeback_15_bits_debugInfo_dispatchTime;
    logic [63:0]  io_writeback_15_bits_debugInfo_enqRsTime;
    logic [63:0]  io_writeback_15_bits_debugInfo_selectTime;
    logic [63:0]  io_writeback_15_bits_debugInfo_issueTime;
    logic [63:0]  io_writeback_15_bits_debugInfo_writebackTime;
    logic [63:0]  io_writeback_15_bits_debugInfo_runahead_checkpoint_id;
    logic [63:0]  io_writeback_15_bits_debugInfo_tlbFirstReqTime;
    logic [63:0]  io_writeback_15_bits_debugInfo_tlbRespTime;
    logic [63:0]  io_writeback_15_bits_debug_seqNum;
    logic         io_writeback_14_valid;
    logic [127:0] io_writeback_14_bits_data_0;
    logic [127:0] io_writeback_14_bits_data_1;
    logic [127:0] io_writeback_14_bits_data_2;
    logic [127:0] io_writeback_14_bits_data_3;
    logic [127:0] io_writeback_14_bits_data_4;
    logic [127:0] io_writeback_14_bits_data_5;
    logic [7:0]   io_writeback_14_bits_pdest;
    logic         io_writeback_14_bits_robIdx_flag;
    logic [7:0]   io_writeback_14_bits_robIdx_value;
    logic         io_writeback_14_bits_intWen;
    logic         io_writeback_14_bits_fpWen;
    logic         io_writeback_14_bits_vecWen;
    logic         io_writeback_14_bits_v0Wen;
    logic         io_writeback_14_bits_vlWen;
    logic [4:0]   io_writeback_14_bits_fflags;
    logic         io_writeback_14_bits_wflags;
    logic         io_writeback_14_bits_exceptionVec_2;
    logic         io_writeback_14_bits_debugInfo_eliminatedMove;
    logic [63:0]  io_writeback_14_bits_debugInfo_renameTime;
    logic [63:0]  io_writeback_14_bits_debugInfo_dispatchTime;
    logic [63:0]  io_writeback_14_bits_debugInfo_enqRsTime;
    logic [63:0]  io_writeback_14_bits_debugInfo_selectTime;
    logic [63:0]  io_writeback_14_bits_debugInfo_issueTime;
    logic [63:0]  io_writeback_14_bits_debugInfo_writebackTime;
    logic [63:0]  io_writeback_14_bits_debugInfo_runahead_checkpoint_id;
    logic [63:0]  io_writeback_14_bits_debugInfo_tlbFirstReqTime;
    logic [63:0]  io_writeback_14_bits_debugInfo_tlbRespTime;
    logic [63:0]  io_writeback_14_bits_debug_seqNum;
    logic         io_writeback_13_valid;
    logic [127:0] io_writeback_13_bits_data_0;
    logic [127:0] io_writeback_13_bits_data_1;
    logic [127:0] io_writeback_13_bits_data_2;
    logic [6:0]   io_writeback_13_bits_pdest;
    logic         io_writeback_13_bits_robIdx_flag;
    logic [7:0]   io_writeback_13_bits_robIdx_value;
    logic         io_writeback_13_bits_vecWen;
    logic         io_writeback_13_bits_v0Wen;
    logic [4:0]   io_writeback_13_bits_fflags;
    logic         io_writeback_13_bits_wflags;
    logic         io_writeback_13_bits_vxsat;
    logic         io_writeback_13_bits_exceptionVec_2;
    logic         io_writeback_13_bits_debugInfo_eliminatedMove;
    logic [63:0]  io_writeback_13_bits_debugInfo_renameTime;
    logic [63:0]  io_writeback_13_bits_debugInfo_dispatchTime;
    logic [63:0]  io_writeback_13_bits_debugInfo_enqRsTime;
    logic [63:0]  io_writeback_13_bits_debugInfo_selectTime;
    logic [63:0]  io_writeback_13_bits_debugInfo_issueTime;
    logic [63:0]  io_writeback_13_bits_debugInfo_writebackTime;
    logic [63:0]  io_writeback_13_bits_debugInfo_runahead_checkpoint_id;
    logic [63:0]  io_writeback_13_bits_debugInfo_tlbFirstReqTime;
    logic [63:0]  io_writeback_13_bits_debugInfo_tlbRespTime;
    logic [63:0]  io_writeback_13_bits_debug_seqNum;
    logic         io_writeback_7_valid ;
    logic [63:0]  io_writeback_7_bits_data_0;
    logic [63:0]  io_writeback_7_bits_data_1;
    logic [7:0]   io_writeback_7_bits_pdest;
    logic         io_writeback_7_bits_robIdx_flag;
    logic [7:0]   io_writeback_7_bits_robIdx_value;
    logic         io_writeback_7_bits_intWen;
    logic         io_writeback_7_bits_redirect_valid;
    logic         io_writeback_7_bits_redirect_bits_isRVC;
    logic         io_writeback_7_bits_redirect_bits_robIdx_flag;
    logic [7:0]   io_writeback_7_bits_redirect_bits_robIdx_value;
    logic         io_writeback_7_bits_redirect_bits_ftqIdx_flag;
    logic [5:0]   io_writeback_7_bits_redirect_bits_ftqIdx_value;
    logic [3:0]   io_writeback_7_bits_redirect_bits_ftqOffset;
    logic         io_writeback_7_bits_redirect_bits_level;
    logic         io_writeback_7_bits_redirect_bits_interrupt;
    logic [49:0]  io_writeback_7_bits_redirect_bits_cfiUpdate_pc;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC;
    logic [1:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet;
    logic [3:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_ssp;
    logic [2:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_sctr;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag;
    logic [4:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag;
    logic [4:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag;
    logic [4:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value;
    logic [49:0]  io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr;
    logic [10:0]  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist;
    logic [10:0]  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist;
    logic [6:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist;
    logic [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist;
    logic [8:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist;
    logic [3:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist;
    logic [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist;
    logic [8:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist;
    logic [6:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist;
    logic [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist;
    logic [6:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist;
    logic [8:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist;
    logic [6:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist;
    logic [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist;
    logic [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist;
    logic [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist;
    logic [10:0]  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist;
    logic [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3;
    logic [2:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH;
    logic [3:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_ghr;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag;
    logic [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value;
    logic [9:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0;
    logic [9:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken;
    logic [49:0]  io_writeback_7_bits_redirect_bits_cfiUpdate_target;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_taken;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred;
    logic [1:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_shift;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF;
    logic         io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF;
    logic [63:0]  io_writeback_7_bits_redirect_bits_fullTarget;
    logic         io_writeback_7_bits_redirect_bits_stFtqIdx_flag;
    logic [5:0]   io_writeback_7_bits_redirect_bits_stFtqIdx_value;
    logic [3:0]   io_writeback_7_bits_redirect_bits_stFtqOffset;
    logic [63:0]  io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id;
    logic         io_writeback_7_bits_redirect_bits_debugIsCtrl;
    logic         io_writeback_7_bits_redirect_bits_debugIsMemVio;
    logic         io_writeback_7_bits_exceptionVec_2;
    logic         io_writeback_7_bits_exceptionVec_3;
    logic         io_writeback_7_bits_exceptionVec_8;
    logic         io_writeback_7_bits_exceptionVec_9;
    logic         io_writeback_7_bits_exceptionVec_10;
    logic         io_writeback_7_bits_exceptionVec_11;
    logic         io_writeback_7_bits_exceptionVec_22;
    logic         io_writeback_7_bits_flushPipe;
    logic         io_writeback_7_bits_predecodeInfo_valid;
    logic         io_writeback_7_bits_predecodeInfo_isRVC;
    logic [1:0]   io_writeback_7_bits_predecodeInfo_brType;
    logic         io_writeback_7_bits_predecodeInfo_isCall;
    logic         io_writeback_7_bits_predecodeInfo_isRet;
    logic         io_writeback_7_bits_debug_isPerfCnt;
    logic         io_writeback_7_bits_debugInfo_eliminatedMove;
    logic [63:0]  io_writeback_7_bits_debugInfo_renameTime;
    logic [63:0]  io_writeback_7_bits_debugInfo_dispatchTime;
    logic [63:0]  io_writeback_7_bits_debugInfo_enqRsTime;
    logic [63:0]  io_writeback_7_bits_debugInfo_selectTime;
    logic [63:0]  io_writeback_7_bits_debugInfo_issueTime;
    logic [63:0]  io_writeback_7_bits_debugInfo_writebackTime;
    logic [63:0]  io_writeback_7_bits_debugInfo_runahead_checkpoint_id;
    logic [63:0]  io_writeback_7_bits_debugInfo_tlbFirstReqTime;
    logic [63:0]  io_writeback_7_bits_debugInfo_tlbRespTime;
    logic [63:0]  io_writeback_7_bits_debug_seqNum;
    logic         io_writeback_5_valid ;
    logic         io_writeback_5_bits_redirect_valid;
    logic         io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred;
    logic         io_writeback_3_valid ;
    logic         io_writeback_3_bits_redirect_valid;
    logic         io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred;
    logic         io_writeback_1_valid ;
    logic         io_writeback_1_bits_redirect_valid;
    logic         io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred;
    logic         io_exuWriteback_26_valid;
    logic [7:0]   io_exuWriteback_26_bits_robIdx_value;
    logic         io_exuWriteback_25_valid;
    logic [7:0]   io_exuWriteback_25_bits_robIdx_value;
    logic         io_exuWriteback_24_valid;
    logic [127:0] io_exuWriteback_24_bits_data_0;
    logic [6:0]   io_exuWriteback_24_bits_pdest;
    logic [7:0]   io_exuWriteback_24_bits_robIdx_value;
    logic         io_exuWriteback_24_bits_vecWen;
    logic         io_exuWriteback_24_bits_v0Wen;
    logic [2:0]   io_exuWriteback_24_bits_vls_vdIdx;
    logic         io_exuWriteback_24_bits_debug_isMMIO;
    logic         io_exuWriteback_24_bits_debug_isNCIO;
    logic         io_exuWriteback_24_bits_debug_isPerfCnt;
    logic [47:0]  io_exuWriteback_24_bits_debug_paddr;
    logic         io_exuWriteback_23_valid;
    logic [127:0] io_exuWriteback_23_bits_data_0;
    logic [6:0]   io_exuWriteback_23_bits_pdest;
    logic [7:0]   io_exuWriteback_23_bits_robIdx_value;
    logic         io_exuWriteback_23_bits_vecWen;
    logic         io_exuWriteback_23_bits_v0Wen;
    logic [2:0]   io_exuWriteback_23_bits_vls_vdIdx;
    logic         io_exuWriteback_23_bits_debug_isMMIO;
    logic         io_exuWriteback_23_bits_debug_isNCIO;
    logic         io_exuWriteback_23_bits_debug_isPerfCnt;
    logic [47:0]  io_exuWriteback_23_bits_debug_paddr;
    logic         io_exuWriteback_22_valid;
    logic [63:0]  io_exuWriteback_22_bits_data_0;
    logic [7:0]   io_exuWriteback_22_bits_robIdx_value;
    logic [6:0]   io_exuWriteback_22_bits_lqIdx_value;
    logic         io_exuWriteback_22_bits_debug_isMMIO;
    logic         io_exuWriteback_22_bits_debug_isNCIO;
    logic         io_exuWriteback_22_bits_debug_isPerfCnt;
    logic [47:0]  io_exuWriteback_22_bits_debug_paddr;
    logic         io_exuWriteback_21_valid;
    logic [63:0]  io_exuWriteback_21_bits_data_0;
    logic [7:0]   io_exuWriteback_21_bits_robIdx_value;
    logic [6:0]   io_exuWriteback_21_bits_lqIdx_value;
    logic         io_exuWriteback_21_bits_debug_isMMIO;
    logic         io_exuWriteback_21_bits_debug_isNCIO;
    logic         io_exuWriteback_21_bits_debug_isPerfCnt;
    logic [47:0]  io_exuWriteback_21_bits_debug_paddr;
    logic         io_exuWriteback_20_valid;
    logic [63:0]  io_exuWriteback_20_bits_data_0;
    logic [7:0]   io_exuWriteback_20_bits_robIdx_value;
    logic [6:0]   io_exuWriteback_20_bits_lqIdx_value;
    logic         io_exuWriteback_20_bits_debug_isMMIO;
    logic         io_exuWriteback_20_bits_debug_isNCIO;
    logic         io_exuWriteback_20_bits_debug_isPerfCnt;
    logic [47:0]  io_exuWriteback_20_bits_debug_paddr;
    logic         io_exuWriteback_19_valid;
    logic [63:0]  io_exuWriteback_19_bits_data_0;
    logic [7:0]   io_exuWriteback_19_bits_robIdx_value;
    logic [5:0]   io_exuWriteback_19_bits_sqIdx_value;
    logic         io_exuWriteback_19_bits_debug_isMMIO;
    logic         io_exuWriteback_19_bits_debug_isNCIO;
    logic         io_exuWriteback_19_bits_debug_isPerfCnt;
    logic [47:0]  io_exuWriteback_19_bits_debug_paddr;
    logic         io_exuWriteback_18_valid;
    logic [63:0]  io_exuWriteback_18_bits_data_0;
    logic [7:0]   io_exuWriteback_18_bits_robIdx_value;
    logic [5:0]   io_exuWriteback_18_bits_sqIdx_value;
    logic         io_exuWriteback_18_bits_debug_isMMIO;
    logic         io_exuWriteback_18_bits_debug_isNCIO;
    logic         io_exuWriteback_18_bits_debug_isPerfCnt;
    logic [47:0]  io_exuWriteback_18_bits_debug_paddr;
    logic         io_exuWriteback_17_valid;
    logic [127:0] io_exuWriteback_17_bits_data_0;
    logic [7:0]   io_exuWriteback_17_bits_robIdx_value;
    logic [4:0]   io_exuWriteback_17_bits_fflags;
    logic         io_exuWriteback_17_bits_wflags;
    logic         io_exuWriteback_16_valid;
    logic [127:0] io_exuWriteback_16_bits_data_0;
    logic [7:0]   io_exuWriteback_16_bits_robIdx_value;
    logic [4:0]   io_exuWriteback_16_bits_fflags;
    logic         io_exuWriteback_16_bits_wflags;
    logic         io_exuWriteback_15_valid;
    logic [127:0] io_exuWriteback_15_bits_data_0;
    logic [7:0]   io_exuWriteback_15_bits_robIdx_value;
    logic [4:0]   io_exuWriteback_15_bits_fflags;
    logic         io_exuWriteback_15_bits_wflags;
    logic         io_exuWriteback_15_bits_vxsat;
    logic         io_exuWriteback_14_valid;
    logic [127:0] io_exuWriteback_14_bits_data_0;
    logic [7:0]   io_exuWriteback_14_bits_robIdx_value;
    logic [4:0]   io_exuWriteback_14_bits_fflags;
    logic         io_exuWriteback_14_bits_wflags;
    logic         io_exuWriteback_13_valid;
    logic [127:0] io_exuWriteback_13_bits_data_0;
    logic [7:0]   io_exuWriteback_13_bits_robIdx_value;
    logic [4:0]   io_exuWriteback_13_bits_fflags;
    logic         io_exuWriteback_13_bits_wflags;
    logic         io_exuWriteback_13_bits_vxsat;
    logic         io_exuWriteback_12_valid;
    logic [63:0]  io_exuWriteback_12_bits_data_0;
    logic [7:0]   io_exuWriteback_12_bits_robIdx_value;
    logic [4:0]   io_exuWriteback_12_bits_fflags;
    logic         io_exuWriteback_12_bits_wflags;
    logic         io_exuWriteback_11_valid;
    logic [63:0]  io_exuWriteback_11_bits_data_0;
    logic [7:0]   io_exuWriteback_11_bits_robIdx_value;
    logic [4:0]   io_exuWriteback_11_bits_fflags;
    logic         io_exuWriteback_11_bits_wflags;
    logic         io_exuWriteback_10_valid;
    logic [63:0]  io_exuWriteback_10_bits_data_0;
    logic [7:0]   io_exuWriteback_10_bits_robIdx_value;
    logic [4:0]   io_exuWriteback_10_bits_fflags;
    logic         io_exuWriteback_10_bits_wflags;
    logic         io_exuWriteback_9_valid;
    logic [63:0]  io_exuWriteback_9_bits_data_0;
    logic [7:0]   io_exuWriteback_9_bits_robIdx_value;
    logic [4:0]   io_exuWriteback_9_bits_fflags;
    logic         io_exuWriteback_9_bits_wflags;
    logic         io_exuWriteback_8_valid;
    logic [127:0] io_exuWriteback_8_bits_data_0;
    logic [7:0]   io_exuWriteback_8_bits_robIdx_value;
    logic [4:0]   io_exuWriteback_8_bits_fflags;
    logic         io_exuWriteback_8_bits_wflags;
    logic         io_exuWriteback_7_valid;
    logic [63:0]  io_exuWriteback_7_bits_data_0;
    logic [7:0]   io_exuWriteback_7_bits_robIdx_value;
    logic         io_exuWriteback_7_bits_debug_isPerfCnt;
    logic         io_exuWriteback_6_valid;
    logic [63:0]  io_exuWriteback_6_bits_data_0;
    logic [7:0]   io_exuWriteback_6_bits_robIdx_value;
    logic         io_exuWriteback_5_valid;
    logic [127:0] io_exuWriteback_5_bits_data_0;
    logic [7:0]   io_exuWriteback_5_bits_robIdx_value;
    logic         io_exuWriteback_5_bits_redirect_valid;
    logic         io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken;
    logic [4:0]   io_exuWriteback_5_bits_fflags;
    logic         io_exuWriteback_5_bits_wflags;
    logic         io_exuWriteback_4_valid;
    logic [63:0]  io_exuWriteback_4_bits_data_0;
    logic [7:0]   io_exuWriteback_4_bits_robIdx_value;
    logic         io_exuWriteback_3_valid;
    logic [63:0]  io_exuWriteback_3_bits_data_0;
    logic [7:0]   io_exuWriteback_3_bits_robIdx_value;
    logic         io_exuWriteback_3_bits_redirect_valid;
    logic         io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken;
    logic         io_exuWriteback_2_valid;
    logic [63:0]  io_exuWriteback_2_bits_data_0;
    logic [7:0]   io_exuWriteback_2_bits_robIdx_value;
    logic         io_exuWriteback_1_valid;
    logic [63:0]  io_exuWriteback_1_bits_data_0;
    logic [7:0]   io_exuWriteback_1_bits_robIdx_value;
    logic         io_exuWriteback_1_bits_redirect_valid;
    logic         io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken;
    logic         io_exuWriteback_0_valid;
    logic [63:0]  io_exuWriteback_0_bits_data_0;
    logic [7:0]   io_exuWriteback_0_bits_robIdx_value;
    logic [4:0]   io_writebackNums_0_bits;
    logic [4:0]   io_writebackNums_1_bits;
    logic [4:0]   io_writebackNums_2_bits;
    logic [4:0]   io_writebackNums_3_bits;
    logic [4:0]   io_writebackNums_4_bits;
    logic [4:0]   io_writebackNums_5_bits;
    logic [4:0]   io_writebackNums_6_bits;
    logic [4:0]   io_writebackNums_7_bits;
    logic [4:0]   io_writebackNums_8_bits;
    logic [4:0]   io_writebackNums_9_bits;
    logic [4:0]   io_writebackNums_10_bits;
    logic [4:0]   io_writebackNums_11_bits;
    logic [4:0]   io_writebackNums_12_bits;
    logic [4:0]   io_writebackNums_13_bits;
    logic [4:0]   io_writebackNums_14_bits;
    logic [4:0]   io_writebackNums_15_bits;
    logic [4:0]   io_writebackNums_16_bits;
    logic [4:0]   io_writebackNums_17_bits;
    logic [4:0]   io_writebackNums_18_bits;
    logic [4:0]   io_writebackNums_19_bits;
    logic [4:0]   io_writebackNums_20_bits;
    logic [4:0]   io_writebackNums_21_bits;
    logic [4:0]   io_writebackNums_22_bits;
    logic [4:0]   io_writebackNums_23_bits;
    logic [4:0]   io_writebackNums_24_bits;
    logic         io_writebackNeedFlush_0;
    logic         io_writebackNeedFlush_1;
    logic         io_writebackNeedFlush_2;
    logic         io_writebackNeedFlush_6;
    logic         io_writebackNeedFlush_7;
    logic         io_writebackNeedFlush_8;
    logic         io_writebackNeedFlush_9;
    logic         io_writebackNeedFlush_10;
    logic         io_writebackNeedFlush_11;
    logic         io_writebackNeedFlush_12;

    clocking drv_cb @(posedge clk);
        `ifdef INTERFACE_ADD_DELAY
            default input #`DEF_SETUP_TIME output #`DEF_HOLD_TIME;
        `endif
        output io_writeback_24_valid;
        output io_writeback_24_bits_data_0;
        output io_writeback_24_bits_pdest;
        output io_writeback_24_bits_robIdx_flag;
        output io_writeback_24_bits_robIdx_value;
        output io_writeback_24_bits_vecWen;
        output io_writeback_24_bits_v0Wen;
        output io_writeback_24_bits_vlWen;
        output io_writeback_24_bits_exceptionVec_0;
        output io_writeback_24_bits_exceptionVec_1;
        output io_writeback_24_bits_exceptionVec_2;
        output io_writeback_24_bits_exceptionVec_3;
        output io_writeback_24_bits_exceptionVec_4;
        output io_writeback_24_bits_exceptionVec_5;
        output io_writeback_24_bits_exceptionVec_6;
        output io_writeback_24_bits_exceptionVec_7;
        output io_writeback_24_bits_exceptionVec_8;
        output io_writeback_24_bits_exceptionVec_9;
        output io_writeback_24_bits_exceptionVec_10;
        output io_writeback_24_bits_exceptionVec_11;
        output io_writeback_24_bits_exceptionVec_12;
        output io_writeback_24_bits_exceptionVec_13;
        output io_writeback_24_bits_exceptionVec_14;
        output io_writeback_24_bits_exceptionVec_15;
        output io_writeback_24_bits_exceptionVec_16;
        output io_writeback_24_bits_exceptionVec_17;
        output io_writeback_24_bits_exceptionVec_18;
        output io_writeback_24_bits_exceptionVec_19;
        output io_writeback_24_bits_exceptionVec_20;
        output io_writeback_24_bits_exceptionVec_21;
        output io_writeback_24_bits_exceptionVec_22;
        output io_writeback_24_bits_exceptionVec_23;
        output io_writeback_24_bits_flushPipe;
        output io_writeback_24_bits_replay;
        output io_writeback_24_bits_trigger;
        output io_writeback_24_bits_vls_vpu_vill;
        output io_writeback_24_bits_vls_vpu_vma;
        output io_writeback_24_bits_vls_vpu_vta;
        output io_writeback_24_bits_vls_vpu_vsew;
        output io_writeback_24_bits_vls_vpu_vlmul;
        output io_writeback_24_bits_vls_vpu_specVill;
        output io_writeback_24_bits_vls_vpu_specVma;
        output io_writeback_24_bits_vls_vpu_specVta;
        output io_writeback_24_bits_vls_vpu_specVsew;
        output io_writeback_24_bits_vls_vpu_specVlmul;
        output io_writeback_24_bits_vls_vpu_vm;
        output io_writeback_24_bits_vls_vpu_vstart;
        output io_writeback_24_bits_vls_vpu_frm;
        output io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst;
        output io_writeback_24_bits_vls_vpu_fpu_isFP32Instr;
        output io_writeback_24_bits_vls_vpu_fpu_isFP64Instr;
        output io_writeback_24_bits_vls_vpu_fpu_isReduction;
        output io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2;
        output io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4;
        output io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8;
        output io_writeback_24_bits_vls_vpu_vxrm;
        output io_writeback_24_bits_vls_vpu_vuopIdx;
        output io_writeback_24_bits_vls_vpu_lastUop;
        output io_writeback_24_bits_vls_vpu_vmask;
        output io_writeback_24_bits_vls_vpu_vl;
        output io_writeback_24_bits_vls_vpu_nf;
        output io_writeback_24_bits_vls_vpu_veew;
        output io_writeback_24_bits_vls_vpu_isReverse;
        output io_writeback_24_bits_vls_vpu_isExt;
        output io_writeback_24_bits_vls_vpu_isNarrow;
        output io_writeback_24_bits_vls_vpu_isDstMask;
        output io_writeback_24_bits_vls_vpu_isOpMask;
        output io_writeback_24_bits_vls_vpu_isMove;
        output io_writeback_24_bits_vls_vpu_isDependOldVd;
        output io_writeback_24_bits_vls_vpu_isWritePartVd;
        output io_writeback_24_bits_vls_vpu_isVleff;
        output io_writeback_24_bits_vls_oldVdPsrc;
        output io_writeback_24_bits_vls_vdIdx;
        output io_writeback_24_bits_vls_vdIdxInField;
        output io_writeback_24_bits_vls_isIndexed;
        output io_writeback_24_bits_vls_isMasked;
        output io_writeback_24_bits_vls_isStrided;
        output io_writeback_24_bits_vls_isWhole;
        output io_writeback_24_bits_vls_isVecLoad;
        output io_writeback_24_bits_vls_isVlm;
        output io_writeback_24_bits_debug_isMMIO;
        output io_writeback_24_bits_debug_isNCIO;
        output io_writeback_24_bits_debug_isPerfCnt;
        output io_writeback_24_bits_debug_paddr;
        output io_writeback_24_bits_debug_vaddr;
        output io_writeback_24_bits_debugInfo_eliminatedMove;
        output io_writeback_24_bits_debugInfo_renameTime;
        output io_writeback_24_bits_debugInfo_dispatchTime;
        output io_writeback_24_bits_debugInfo_enqRsTime;
        output io_writeback_24_bits_debugInfo_selectTime;
        output io_writeback_24_bits_debugInfo_issueTime;
        output io_writeback_24_bits_debugInfo_writebackTime;
        output io_writeback_24_bits_debugInfo_runahead_checkpoint_id;
        output io_writeback_24_bits_debugInfo_tlbFirstReqTime;
        output io_writeback_24_bits_debugInfo_tlbRespTime;
        output io_writeback_24_bits_debug_seqNum;
        output io_writeback_23_valid;
        output io_writeback_23_bits_data_0;
        output io_writeback_23_bits_pdest;
        output io_writeback_23_bits_robIdx_flag;
        output io_writeback_23_bits_robIdx_value;
        output io_writeback_23_bits_vecWen;
        output io_writeback_23_bits_v0Wen;
        output io_writeback_23_bits_vlWen;
        output io_writeback_23_bits_exceptionVec_0;
        output io_writeback_23_bits_exceptionVec_1;
        output io_writeback_23_bits_exceptionVec_2;
        output io_writeback_23_bits_exceptionVec_3;
        output io_writeback_23_bits_exceptionVec_4;
        output io_writeback_23_bits_exceptionVec_5;
        output io_writeback_23_bits_exceptionVec_6;
        output io_writeback_23_bits_exceptionVec_7;
        output io_writeback_23_bits_exceptionVec_8;
        output io_writeback_23_bits_exceptionVec_9;
        output io_writeback_23_bits_exceptionVec_10;
        output io_writeback_23_bits_exceptionVec_11;
        output io_writeback_23_bits_exceptionVec_12;
        output io_writeback_23_bits_exceptionVec_13;
        output io_writeback_23_bits_exceptionVec_14;
        output io_writeback_23_bits_exceptionVec_15;
        output io_writeback_23_bits_exceptionVec_16;
        output io_writeback_23_bits_exceptionVec_17;
        output io_writeback_23_bits_exceptionVec_18;
        output io_writeback_23_bits_exceptionVec_19;
        output io_writeback_23_bits_exceptionVec_20;
        output io_writeback_23_bits_exceptionVec_21;
        output io_writeback_23_bits_exceptionVec_22;
        output io_writeback_23_bits_exceptionVec_23;
        output io_writeback_23_bits_flushPipe;
        output io_writeback_23_bits_replay;
        output io_writeback_23_bits_trigger;
        output io_writeback_23_bits_vls_vpu_vill;
        output io_writeback_23_bits_vls_vpu_vma;
        output io_writeback_23_bits_vls_vpu_vta;
        output io_writeback_23_bits_vls_vpu_vsew;
        output io_writeback_23_bits_vls_vpu_vlmul;
        output io_writeback_23_bits_vls_vpu_specVill;
        output io_writeback_23_bits_vls_vpu_specVma;
        output io_writeback_23_bits_vls_vpu_specVta;
        output io_writeback_23_bits_vls_vpu_specVsew;
        output io_writeback_23_bits_vls_vpu_specVlmul;
        output io_writeback_23_bits_vls_vpu_vm;
        output io_writeback_23_bits_vls_vpu_vstart;
        output io_writeback_23_bits_vls_vpu_frm;
        output io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst;
        output io_writeback_23_bits_vls_vpu_fpu_isFP32Instr;
        output io_writeback_23_bits_vls_vpu_fpu_isFP64Instr;
        output io_writeback_23_bits_vls_vpu_fpu_isReduction;
        output io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2;
        output io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4;
        output io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8;
        output io_writeback_23_bits_vls_vpu_vxrm;
        output io_writeback_23_bits_vls_vpu_vuopIdx;
        output io_writeback_23_bits_vls_vpu_lastUop;
        output io_writeback_23_bits_vls_vpu_vmask;
        output io_writeback_23_bits_vls_vpu_vl;
        output io_writeback_23_bits_vls_vpu_nf;
        output io_writeback_23_bits_vls_vpu_veew;
        output io_writeback_23_bits_vls_vpu_isReverse;
        output io_writeback_23_bits_vls_vpu_isExt;
        output io_writeback_23_bits_vls_vpu_isNarrow;
        output io_writeback_23_bits_vls_vpu_isDstMask;
        output io_writeback_23_bits_vls_vpu_isOpMask;
        output io_writeback_23_bits_vls_vpu_isMove;
        output io_writeback_23_bits_vls_vpu_isDependOldVd;
        output io_writeback_23_bits_vls_vpu_isWritePartVd;
        output io_writeback_23_bits_vls_vpu_isVleff;
        output io_writeback_23_bits_vls_oldVdPsrc;
        output io_writeback_23_bits_vls_vdIdx;
        output io_writeback_23_bits_vls_vdIdxInField;
        output io_writeback_23_bits_vls_isIndexed;
        output io_writeback_23_bits_vls_isMasked;
        output io_writeback_23_bits_vls_isStrided;
        output io_writeback_23_bits_vls_isWhole;
        output io_writeback_23_bits_vls_isVecLoad;
        output io_writeback_23_bits_vls_isVlm;
        output io_writeback_23_bits_debug_isMMIO;
        output io_writeback_23_bits_debug_isNCIO;
        output io_writeback_23_bits_debug_isPerfCnt;
        output io_writeback_23_bits_debug_paddr;
        output io_writeback_23_bits_debug_vaddr;
        output io_writeback_23_bits_debugInfo_eliminatedMove;
        output io_writeback_23_bits_debugInfo_renameTime;
        output io_writeback_23_bits_debugInfo_dispatchTime;
        output io_writeback_23_bits_debugInfo_enqRsTime;
        output io_writeback_23_bits_debugInfo_selectTime;
        output io_writeback_23_bits_debugInfo_issueTime;
        output io_writeback_23_bits_debugInfo_writebackTime;
        output io_writeback_23_bits_debugInfo_runahead_checkpoint_id;
        output io_writeback_23_bits_debugInfo_tlbFirstReqTime;
        output io_writeback_23_bits_debugInfo_tlbRespTime;
        output io_writeback_23_bits_debug_seqNum;
        output io_writeback_22_valid;
        output io_writeback_22_bits_data_0;
        output io_writeback_22_bits_pdest;
        output io_writeback_22_bits_robIdx_flag;
        output io_writeback_22_bits_robIdx_value;
        output io_writeback_22_bits_intWen;
        output io_writeback_22_bits_fpWen;
        output io_writeback_22_bits_exceptionVec_0;
        output io_writeback_22_bits_exceptionVec_1;
        output io_writeback_22_bits_exceptionVec_2;
        output io_writeback_22_bits_exceptionVec_3;
        output io_writeback_22_bits_exceptionVec_4;
        output io_writeback_22_bits_exceptionVec_5;
        output io_writeback_22_bits_exceptionVec_6;
        output io_writeback_22_bits_exceptionVec_7;
        output io_writeback_22_bits_exceptionVec_8;
        output io_writeback_22_bits_exceptionVec_9;
        output io_writeback_22_bits_exceptionVec_10;
        output io_writeback_22_bits_exceptionVec_11;
        output io_writeback_22_bits_exceptionVec_12;
        output io_writeback_22_bits_exceptionVec_13;
        output io_writeback_22_bits_exceptionVec_14;
        output io_writeback_22_bits_exceptionVec_15;
        output io_writeback_22_bits_exceptionVec_16;
        output io_writeback_22_bits_exceptionVec_17;
        output io_writeback_22_bits_exceptionVec_18;
        output io_writeback_22_bits_exceptionVec_19;
        output io_writeback_22_bits_exceptionVec_20;
        output io_writeback_22_bits_exceptionVec_21;
        output io_writeback_22_bits_exceptionVec_22;
        output io_writeback_22_bits_exceptionVec_23;
        output io_writeback_22_bits_flushPipe;
        output io_writeback_22_bits_replay;
        output io_writeback_22_bits_lqIdx_flag;
        output io_writeback_22_bits_lqIdx_value;
        output io_writeback_22_bits_trigger;
        output io_writeback_22_bits_predecodeInfo_valid;
        output io_writeback_22_bits_predecodeInfo_isRVC;
        output io_writeback_22_bits_predecodeInfo_brType;
        output io_writeback_22_bits_predecodeInfo_isCall;
        output io_writeback_22_bits_predecodeInfo_isRet;
        output io_writeback_22_bits_debug_isMMIO;
        output io_writeback_22_bits_debug_isNCIO;
        output io_writeback_22_bits_debug_isPerfCnt;
        output io_writeback_22_bits_debug_paddr;
        output io_writeback_22_bits_debug_vaddr;
        output io_writeback_22_bits_debugInfo_eliminatedMove;
        output io_writeback_22_bits_debugInfo_renameTime;
        output io_writeback_22_bits_debugInfo_dispatchTime;
        output io_writeback_22_bits_debugInfo_enqRsTime;
        output io_writeback_22_bits_debugInfo_selectTime;
        output io_writeback_22_bits_debugInfo_issueTime;
        output io_writeback_22_bits_debugInfo_writebackTime;
        output io_writeback_22_bits_debugInfo_runahead_checkpoint_id;
        output io_writeback_22_bits_debugInfo_tlbFirstReqTime;
        output io_writeback_22_bits_debugInfo_tlbRespTime;
        output io_writeback_22_bits_debug_seqNum;
        output io_writeback_21_valid;
        output io_writeback_21_bits_data_0;
        output io_writeback_21_bits_pdest;
        output io_writeback_21_bits_robIdx_flag;
        output io_writeback_21_bits_robIdx_value;
        output io_writeback_21_bits_intWen;
        output io_writeback_21_bits_fpWen;
        output io_writeback_21_bits_exceptionVec_0;
        output io_writeback_21_bits_exceptionVec_1;
        output io_writeback_21_bits_exceptionVec_2;
        output io_writeback_21_bits_exceptionVec_3;
        output io_writeback_21_bits_exceptionVec_4;
        output io_writeback_21_bits_exceptionVec_5;
        output io_writeback_21_bits_exceptionVec_6;
        output io_writeback_21_bits_exceptionVec_7;
        output io_writeback_21_bits_exceptionVec_8;
        output io_writeback_21_bits_exceptionVec_9;
        output io_writeback_21_bits_exceptionVec_10;
        output io_writeback_21_bits_exceptionVec_11;
        output io_writeback_21_bits_exceptionVec_12;
        output io_writeback_21_bits_exceptionVec_13;
        output io_writeback_21_bits_exceptionVec_14;
        output io_writeback_21_bits_exceptionVec_15;
        output io_writeback_21_bits_exceptionVec_16;
        output io_writeback_21_bits_exceptionVec_17;
        output io_writeback_21_bits_exceptionVec_18;
        output io_writeback_21_bits_exceptionVec_19;
        output io_writeback_21_bits_exceptionVec_20;
        output io_writeback_21_bits_exceptionVec_21;
        output io_writeback_21_bits_exceptionVec_22;
        output io_writeback_21_bits_exceptionVec_23;
        output io_writeback_21_bits_flushPipe;
        output io_writeback_21_bits_replay;
        output io_writeback_21_bits_lqIdx_flag;
        output io_writeback_21_bits_lqIdx_value;
        output io_writeback_21_bits_trigger;
        output io_writeback_21_bits_predecodeInfo_valid;
        output io_writeback_21_bits_predecodeInfo_isRVC;
        output io_writeback_21_bits_predecodeInfo_brType;
        output io_writeback_21_bits_predecodeInfo_isCall;
        output io_writeback_21_bits_predecodeInfo_isRet;
        output io_writeback_21_bits_debug_isMMIO;
        output io_writeback_21_bits_debug_isNCIO;
        output io_writeback_21_bits_debug_isPerfCnt;
        output io_writeback_21_bits_debug_paddr;
        output io_writeback_21_bits_debug_vaddr;
        output io_writeback_21_bits_debugInfo_eliminatedMove;
        output io_writeback_21_bits_debugInfo_renameTime;
        output io_writeback_21_bits_debugInfo_dispatchTime;
        output io_writeback_21_bits_debugInfo_enqRsTime;
        output io_writeback_21_bits_debugInfo_selectTime;
        output io_writeback_21_bits_debugInfo_issueTime;
        output io_writeback_21_bits_debugInfo_writebackTime;
        output io_writeback_21_bits_debugInfo_runahead_checkpoint_id;
        output io_writeback_21_bits_debugInfo_tlbFirstReqTime;
        output io_writeback_21_bits_debugInfo_tlbRespTime;
        output io_writeback_21_bits_debug_seqNum;
        output io_writeback_20_valid;
        output io_writeback_20_bits_data_0;
        output io_writeback_20_bits_pdest;
        output io_writeback_20_bits_robIdx_flag;
        output io_writeback_20_bits_robIdx_value;
        output io_writeback_20_bits_intWen;
        output io_writeback_20_bits_fpWen;
        output io_writeback_20_bits_exceptionVec_0;
        output io_writeback_20_bits_exceptionVec_1;
        output io_writeback_20_bits_exceptionVec_2;
        output io_writeback_20_bits_exceptionVec_3;
        output io_writeback_20_bits_exceptionVec_4;
        output io_writeback_20_bits_exceptionVec_5;
        output io_writeback_20_bits_exceptionVec_6;
        output io_writeback_20_bits_exceptionVec_7;
        output io_writeback_20_bits_exceptionVec_8;
        output io_writeback_20_bits_exceptionVec_9;
        output io_writeback_20_bits_exceptionVec_10;
        output io_writeback_20_bits_exceptionVec_11;
        output io_writeback_20_bits_exceptionVec_12;
        output io_writeback_20_bits_exceptionVec_13;
        output io_writeback_20_bits_exceptionVec_14;
        output io_writeback_20_bits_exceptionVec_15;
        output io_writeback_20_bits_exceptionVec_16;
        output io_writeback_20_bits_exceptionVec_17;
        output io_writeback_20_bits_exceptionVec_18;
        output io_writeback_20_bits_exceptionVec_19;
        output io_writeback_20_bits_exceptionVec_20;
        output io_writeback_20_bits_exceptionVec_21;
        output io_writeback_20_bits_exceptionVec_22;
        output io_writeback_20_bits_exceptionVec_23;
        output io_writeback_20_bits_flushPipe;
        output io_writeback_20_bits_replay;
        output io_writeback_20_bits_lqIdx_flag;
        output io_writeback_20_bits_lqIdx_value;
        output io_writeback_20_bits_trigger;
        output io_writeback_20_bits_predecodeInfo_valid;
        output io_writeback_20_bits_predecodeInfo_isRVC;
        output io_writeback_20_bits_predecodeInfo_brType;
        output io_writeback_20_bits_predecodeInfo_isCall;
        output io_writeback_20_bits_predecodeInfo_isRet;
        output io_writeback_20_bits_debug_isMMIO;
        output io_writeback_20_bits_debug_isNCIO;
        output io_writeback_20_bits_debug_isPerfCnt;
        output io_writeback_20_bits_debug_paddr;
        output io_writeback_20_bits_debug_vaddr;
        output io_writeback_20_bits_debugInfo_eliminatedMove;
        output io_writeback_20_bits_debugInfo_renameTime;
        output io_writeback_20_bits_debugInfo_dispatchTime;
        output io_writeback_20_bits_debugInfo_enqRsTime;
        output io_writeback_20_bits_debugInfo_selectTime;
        output io_writeback_20_bits_debugInfo_issueTime;
        output io_writeback_20_bits_debugInfo_writebackTime;
        output io_writeback_20_bits_debugInfo_runahead_checkpoint_id;
        output io_writeback_20_bits_debugInfo_tlbFirstReqTime;
        output io_writeback_20_bits_debugInfo_tlbRespTime;
        output io_writeback_20_bits_debug_seqNum;
        output io_writeback_19_valid;
        output io_writeback_19_bits_data_0;
        output io_writeback_19_bits_pdest;
        output io_writeback_19_bits_robIdx_flag;
        output io_writeback_19_bits_robIdx_value;
        output io_writeback_19_bits_intWen;
        output io_writeback_19_bits_exceptionVec_0;
        output io_writeback_19_bits_exceptionVec_1;
        output io_writeback_19_bits_exceptionVec_2;
        output io_writeback_19_bits_exceptionVec_3;
        output io_writeback_19_bits_exceptionVec_4;
        output io_writeback_19_bits_exceptionVec_5;
        output io_writeback_19_bits_exceptionVec_6;
        output io_writeback_19_bits_exceptionVec_7;
        output io_writeback_19_bits_exceptionVec_8;
        output io_writeback_19_bits_exceptionVec_9;
        output io_writeback_19_bits_exceptionVec_10;
        output io_writeback_19_bits_exceptionVec_11;
        output io_writeback_19_bits_exceptionVec_12;
        output io_writeback_19_bits_exceptionVec_13;
        output io_writeback_19_bits_exceptionVec_14;
        output io_writeback_19_bits_exceptionVec_15;
        output io_writeback_19_bits_exceptionVec_16;
        output io_writeback_19_bits_exceptionVec_17;
        output io_writeback_19_bits_exceptionVec_18;
        output io_writeback_19_bits_exceptionVec_19;
        output io_writeback_19_bits_exceptionVec_20;
        output io_writeback_19_bits_exceptionVec_21;
        output io_writeback_19_bits_exceptionVec_22;
        output io_writeback_19_bits_exceptionVec_23;
        output io_writeback_19_bits_flushPipe;
        output io_writeback_19_bits_sqIdx_flag;
        output io_writeback_19_bits_sqIdx_value;
        output io_writeback_19_bits_trigger;
        output io_writeback_19_bits_debug_isMMIO;
        output io_writeback_19_bits_debug_isNCIO;
        output io_writeback_19_bits_debug_isPerfCnt;
        output io_writeback_19_bits_debug_paddr;
        output io_writeback_19_bits_debug_vaddr;
        output io_writeback_19_bits_debugInfo_eliminatedMove;
        output io_writeback_19_bits_debugInfo_renameTime;
        output io_writeback_19_bits_debugInfo_dispatchTime;
        output io_writeback_19_bits_debugInfo_enqRsTime;
        output io_writeback_19_bits_debugInfo_selectTime;
        output io_writeback_19_bits_debugInfo_issueTime;
        output io_writeback_19_bits_debugInfo_writebackTime;
        output io_writeback_19_bits_debugInfo_runahead_checkpoint_id;
        output io_writeback_19_bits_debugInfo_tlbFirstReqTime;
        output io_writeback_19_bits_debugInfo_tlbRespTime;
        output io_writeback_19_bits_debug_seqNum;
        output io_writeback_18_valid;
        output io_writeback_18_bits_data_0;
        output io_writeback_18_bits_pdest;
        output io_writeback_18_bits_robIdx_flag;
        output io_writeback_18_bits_robIdx_value;
        output io_writeback_18_bits_intWen;
        output io_writeback_18_bits_exceptionVec_0;
        output io_writeback_18_bits_exceptionVec_1;
        output io_writeback_18_bits_exceptionVec_2;
        output io_writeback_18_bits_exceptionVec_3;
        output io_writeback_18_bits_exceptionVec_4;
        output io_writeback_18_bits_exceptionVec_5;
        output io_writeback_18_bits_exceptionVec_6;
        output io_writeback_18_bits_exceptionVec_7;
        output io_writeback_18_bits_exceptionVec_8;
        output io_writeback_18_bits_exceptionVec_9;
        output io_writeback_18_bits_exceptionVec_10;
        output io_writeback_18_bits_exceptionVec_11;
        output io_writeback_18_bits_exceptionVec_12;
        output io_writeback_18_bits_exceptionVec_13;
        output io_writeback_18_bits_exceptionVec_14;
        output io_writeback_18_bits_exceptionVec_15;
        output io_writeback_18_bits_exceptionVec_16;
        output io_writeback_18_bits_exceptionVec_17;
        output io_writeback_18_bits_exceptionVec_18;
        output io_writeback_18_bits_exceptionVec_19;
        output io_writeback_18_bits_exceptionVec_20;
        output io_writeback_18_bits_exceptionVec_21;
        output io_writeback_18_bits_exceptionVec_22;
        output io_writeback_18_bits_exceptionVec_23;
        output io_writeback_18_bits_flushPipe;
        output io_writeback_18_bits_sqIdx_flag;
        output io_writeback_18_bits_sqIdx_value;
        output io_writeback_18_bits_trigger;
        output io_writeback_18_bits_debug_isMMIO;
        output io_writeback_18_bits_debug_isNCIO;
        output io_writeback_18_bits_debug_isPerfCnt;
        output io_writeback_18_bits_debug_paddr;
        output io_writeback_18_bits_debug_vaddr;
        output io_writeback_18_bits_debugInfo_eliminatedMove;
        output io_writeback_18_bits_debugInfo_renameTime;
        output io_writeback_18_bits_debugInfo_dispatchTime;
        output io_writeback_18_bits_debugInfo_enqRsTime;
        output io_writeback_18_bits_debugInfo_selectTime;
        output io_writeback_18_bits_debugInfo_issueTime;
        output io_writeback_18_bits_debugInfo_writebackTime;
        output io_writeback_18_bits_debugInfo_runahead_checkpoint_id;
        output io_writeback_18_bits_debugInfo_tlbFirstReqTime;
        output io_writeback_18_bits_debugInfo_tlbRespTime;
        output io_writeback_18_bits_debug_seqNum;
        output io_writeback_17_valid;
        output io_writeback_17_bits_data_0;
        output io_writeback_17_bits_data_1;
        output io_writeback_17_bits_data_2;
        output io_writeback_17_bits_pdest;
        output io_writeback_17_bits_robIdx_flag;
        output io_writeback_17_bits_robIdx_value;
        output io_writeback_17_bits_vecWen;
        output io_writeback_17_bits_v0Wen;
        output io_writeback_17_bits_fflags;
        output io_writeback_17_bits_wflags;
        output io_writeback_17_bits_debugInfo_eliminatedMove;
        output io_writeback_17_bits_debugInfo_renameTime;
        output io_writeback_17_bits_debugInfo_dispatchTime;
        output io_writeback_17_bits_debugInfo_enqRsTime;
        output io_writeback_17_bits_debugInfo_selectTime;
        output io_writeback_17_bits_debugInfo_issueTime;
        output io_writeback_17_bits_debugInfo_writebackTime;
        output io_writeback_17_bits_debugInfo_runahead_checkpoint_id;
        output io_writeback_17_bits_debugInfo_tlbFirstReqTime;
        output io_writeback_17_bits_debugInfo_tlbRespTime;
        output io_writeback_17_bits_debug_seqNum;
        output io_writeback_16_valid;
        output io_writeback_16_bits_data_0;
        output io_writeback_16_bits_data_1;
        output io_writeback_16_bits_data_2;
        output io_writeback_16_bits_data_3;
        output io_writeback_16_bits_pdest;
        output io_writeback_16_bits_robIdx_flag;
        output io_writeback_16_bits_robIdx_value;
        output io_writeback_16_bits_fpWen;
        output io_writeback_16_bits_vecWen;
        output io_writeback_16_bits_v0Wen;
        output io_writeback_16_bits_fflags;
        output io_writeback_16_bits_wflags;
        output io_writeback_16_bits_debugInfo_eliminatedMove;
        output io_writeback_16_bits_debugInfo_renameTime;
        output io_writeback_16_bits_debugInfo_dispatchTime;
        output io_writeback_16_bits_debugInfo_enqRsTime;
        output io_writeback_16_bits_debugInfo_selectTime;
        output io_writeback_16_bits_debugInfo_issueTime;
        output io_writeback_16_bits_debugInfo_writebackTime;
        output io_writeback_16_bits_debugInfo_runahead_checkpoint_id;
        output io_writeback_16_bits_debugInfo_tlbFirstReqTime;
        output io_writeback_16_bits_debugInfo_tlbRespTime;
        output io_writeback_16_bits_debug_seqNum;
        output io_writeback_15_valid;
        output io_writeback_15_bits_data_0;
        output io_writeback_15_bits_data_1;
        output io_writeback_15_bits_data_2;
        output io_writeback_15_bits_pdest;
        output io_writeback_15_bits_robIdx_flag;
        output io_writeback_15_bits_robIdx_value;
        output io_writeback_15_bits_vecWen;
        output io_writeback_15_bits_v0Wen;
        output io_writeback_15_bits_fflags;
        output io_writeback_15_bits_wflags;
        output io_writeback_15_bits_vxsat;
        output io_writeback_15_bits_debugInfo_eliminatedMove;
        output io_writeback_15_bits_debugInfo_renameTime;
        output io_writeback_15_bits_debugInfo_dispatchTime;
        output io_writeback_15_bits_debugInfo_enqRsTime;
        output io_writeback_15_bits_debugInfo_selectTime;
        output io_writeback_15_bits_debugInfo_issueTime;
        output io_writeback_15_bits_debugInfo_writebackTime;
        output io_writeback_15_bits_debugInfo_runahead_checkpoint_id;
        output io_writeback_15_bits_debugInfo_tlbFirstReqTime;
        output io_writeback_15_bits_debugInfo_tlbRespTime;
        output io_writeback_15_bits_debug_seqNum;
        output io_writeback_14_valid;
        output io_writeback_14_bits_data_0;
        output io_writeback_14_bits_data_1;
        output io_writeback_14_bits_data_2;
        output io_writeback_14_bits_data_3;
        output io_writeback_14_bits_data_4;
        output io_writeback_14_bits_data_5;
        output io_writeback_14_bits_pdest;
        output io_writeback_14_bits_robIdx_flag;
        output io_writeback_14_bits_robIdx_value;
        output io_writeback_14_bits_intWen;
        output io_writeback_14_bits_fpWen;
        output io_writeback_14_bits_vecWen;
        output io_writeback_14_bits_v0Wen;
        output io_writeback_14_bits_vlWen;
        output io_writeback_14_bits_fflags;
        output io_writeback_14_bits_wflags;
        output io_writeback_14_bits_exceptionVec_2;
        output io_writeback_14_bits_debugInfo_eliminatedMove;
        output io_writeback_14_bits_debugInfo_renameTime;
        output io_writeback_14_bits_debugInfo_dispatchTime;
        output io_writeback_14_bits_debugInfo_enqRsTime;
        output io_writeback_14_bits_debugInfo_selectTime;
        output io_writeback_14_bits_debugInfo_issueTime;
        output io_writeback_14_bits_debugInfo_writebackTime;
        output io_writeback_14_bits_debugInfo_runahead_checkpoint_id;
        output io_writeback_14_bits_debugInfo_tlbFirstReqTime;
        output io_writeback_14_bits_debugInfo_tlbRespTime;
        output io_writeback_14_bits_debug_seqNum;
        output io_writeback_13_valid;
        output io_writeback_13_bits_data_0;
        output io_writeback_13_bits_data_1;
        output io_writeback_13_bits_data_2;
        output io_writeback_13_bits_pdest;
        output io_writeback_13_bits_robIdx_flag;
        output io_writeback_13_bits_robIdx_value;
        output io_writeback_13_bits_vecWen;
        output io_writeback_13_bits_v0Wen;
        output io_writeback_13_bits_fflags;
        output io_writeback_13_bits_wflags;
        output io_writeback_13_bits_vxsat;
        output io_writeback_13_bits_exceptionVec_2;
        output io_writeback_13_bits_debugInfo_eliminatedMove;
        output io_writeback_13_bits_debugInfo_renameTime;
        output io_writeback_13_bits_debugInfo_dispatchTime;
        output io_writeback_13_bits_debugInfo_enqRsTime;
        output io_writeback_13_bits_debugInfo_selectTime;
        output io_writeback_13_bits_debugInfo_issueTime;
        output io_writeback_13_bits_debugInfo_writebackTime;
        output io_writeback_13_bits_debugInfo_runahead_checkpoint_id;
        output io_writeback_13_bits_debugInfo_tlbFirstReqTime;
        output io_writeback_13_bits_debugInfo_tlbRespTime;
        output io_writeback_13_bits_debug_seqNum;
        output io_writeback_7_valid;
        output io_writeback_7_bits_data_0;
        output io_writeback_7_bits_data_1;
        output io_writeback_7_bits_pdest;
        output io_writeback_7_bits_robIdx_flag;
        output io_writeback_7_bits_robIdx_value;
        output io_writeback_7_bits_intWen;
        output io_writeback_7_bits_redirect_valid;
        output io_writeback_7_bits_redirect_bits_isRVC;
        output io_writeback_7_bits_redirect_bits_robIdx_flag;
        output io_writeback_7_bits_redirect_bits_robIdx_value;
        output io_writeback_7_bits_redirect_bits_ftqIdx_flag;
        output io_writeback_7_bits_redirect_bits_ftqIdx_value;
        output io_writeback_7_bits_redirect_bits_ftqOffset;
        output io_writeback_7_bits_redirect_bits_level;
        output io_writeback_7_bits_redirect_bits_interrupt;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_pc;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_ssp;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_sctr;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_ghr;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_target;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_taken;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_shift;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF;
        output io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF;
        output io_writeback_7_bits_redirect_bits_fullTarget;
        output io_writeback_7_bits_redirect_bits_stFtqIdx_flag;
        output io_writeback_7_bits_redirect_bits_stFtqIdx_value;
        output io_writeback_7_bits_redirect_bits_stFtqOffset;
        output io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id;
        output io_writeback_7_bits_redirect_bits_debugIsCtrl;
        output io_writeback_7_bits_redirect_bits_debugIsMemVio;
        output io_writeback_7_bits_exceptionVec_2;
        output io_writeback_7_bits_exceptionVec_3;
        output io_writeback_7_bits_exceptionVec_8;
        output io_writeback_7_bits_exceptionVec_9;
        output io_writeback_7_bits_exceptionVec_10;
        output io_writeback_7_bits_exceptionVec_11;
        output io_writeback_7_bits_exceptionVec_22;
        output io_writeback_7_bits_flushPipe;
        output io_writeback_7_bits_predecodeInfo_valid;
        output io_writeback_7_bits_predecodeInfo_isRVC;
        output io_writeback_7_bits_predecodeInfo_brType;
        output io_writeback_7_bits_predecodeInfo_isCall;
        output io_writeback_7_bits_predecodeInfo_isRet;
        output io_writeback_7_bits_debug_isPerfCnt;
        output io_writeback_7_bits_debugInfo_eliminatedMove;
        output io_writeback_7_bits_debugInfo_renameTime;
        output io_writeback_7_bits_debugInfo_dispatchTime;
        output io_writeback_7_bits_debugInfo_enqRsTime;
        output io_writeback_7_bits_debugInfo_selectTime;
        output io_writeback_7_bits_debugInfo_issueTime;
        output io_writeback_7_bits_debugInfo_writebackTime;
        output io_writeback_7_bits_debugInfo_runahead_checkpoint_id;
        output io_writeback_7_bits_debugInfo_tlbFirstReqTime;
        output io_writeback_7_bits_debugInfo_tlbRespTime;
        output io_writeback_7_bits_debug_seqNum;
        output io_writeback_5_valid;
        output io_writeback_5_bits_redirect_valid;
        output io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred;
        output io_writeback_3_valid;
        output io_writeback_3_bits_redirect_valid;
        output io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred;
        output io_writeback_1_valid;
        output io_writeback_1_bits_redirect_valid;
        output io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred;
        output io_exuWriteback_26_valid;
        output io_exuWriteback_26_bits_robIdx_value;
        output io_exuWriteback_25_valid;
        output io_exuWriteback_25_bits_robIdx_value;
        output io_exuWriteback_24_valid;
        output io_exuWriteback_24_bits_data_0;
        output io_exuWriteback_24_bits_pdest;
        output io_exuWriteback_24_bits_robIdx_value;
        output io_exuWriteback_24_bits_vecWen;
        output io_exuWriteback_24_bits_v0Wen;
        output io_exuWriteback_24_bits_vls_vdIdx;
        output io_exuWriteback_24_bits_debug_isMMIO;
        output io_exuWriteback_24_bits_debug_isNCIO;
        output io_exuWriteback_24_bits_debug_isPerfCnt;
        output io_exuWriteback_24_bits_debug_paddr;
        output io_exuWriteback_23_valid;
        output io_exuWriteback_23_bits_data_0;
        output io_exuWriteback_23_bits_pdest;
        output io_exuWriteback_23_bits_robIdx_value;
        output io_exuWriteback_23_bits_vecWen;
        output io_exuWriteback_23_bits_v0Wen;
        output io_exuWriteback_23_bits_vls_vdIdx;
        output io_exuWriteback_23_bits_debug_isMMIO;
        output io_exuWriteback_23_bits_debug_isNCIO;
        output io_exuWriteback_23_bits_debug_isPerfCnt;
        output io_exuWriteback_23_bits_debug_paddr;
        output io_exuWriteback_22_valid;
        output io_exuWriteback_22_bits_data_0;
        output io_exuWriteback_22_bits_robIdx_value;
        output io_exuWriteback_22_bits_lqIdx_value;
        output io_exuWriteback_22_bits_debug_isMMIO;
        output io_exuWriteback_22_bits_debug_isNCIO;
        output io_exuWriteback_22_bits_debug_isPerfCnt;
        output io_exuWriteback_22_bits_debug_paddr;
        output io_exuWriteback_21_valid;
        output io_exuWriteback_21_bits_data_0;
        output io_exuWriteback_21_bits_robIdx_value;
        output io_exuWriteback_21_bits_lqIdx_value;
        output io_exuWriteback_21_bits_debug_isMMIO;
        output io_exuWriteback_21_bits_debug_isNCIO;
        output io_exuWriteback_21_bits_debug_isPerfCnt;
        output io_exuWriteback_21_bits_debug_paddr;
        output io_exuWriteback_20_valid;
        output io_exuWriteback_20_bits_data_0;
        output io_exuWriteback_20_bits_robIdx_value;
        output io_exuWriteback_20_bits_lqIdx_value;
        output io_exuWriteback_20_bits_debug_isMMIO;
        output io_exuWriteback_20_bits_debug_isNCIO;
        output io_exuWriteback_20_bits_debug_isPerfCnt;
        output io_exuWriteback_20_bits_debug_paddr;
        output io_exuWriteback_19_valid;
        output io_exuWriteback_19_bits_data_0;
        output io_exuWriteback_19_bits_robIdx_value;
        output io_exuWriteback_19_bits_sqIdx_value;
        output io_exuWriteback_19_bits_debug_isMMIO;
        output io_exuWriteback_19_bits_debug_isNCIO;
        output io_exuWriteback_19_bits_debug_isPerfCnt;
        output io_exuWriteback_19_bits_debug_paddr;
        output io_exuWriteback_18_valid;
        output io_exuWriteback_18_bits_data_0;
        output io_exuWriteback_18_bits_robIdx_value;
        output io_exuWriteback_18_bits_sqIdx_value;
        output io_exuWriteback_18_bits_debug_isMMIO;
        output io_exuWriteback_18_bits_debug_isNCIO;
        output io_exuWriteback_18_bits_debug_isPerfCnt;
        output io_exuWriteback_18_bits_debug_paddr;
        output io_exuWriteback_17_valid;
        output io_exuWriteback_17_bits_data_0;
        output io_exuWriteback_17_bits_robIdx_value;
        output io_exuWriteback_17_bits_fflags;
        output io_exuWriteback_17_bits_wflags;
        output io_exuWriteback_16_valid;
        output io_exuWriteback_16_bits_data_0;
        output io_exuWriteback_16_bits_robIdx_value;
        output io_exuWriteback_16_bits_fflags;
        output io_exuWriteback_16_bits_wflags;
        output io_exuWriteback_15_valid;
        output io_exuWriteback_15_bits_data_0;
        output io_exuWriteback_15_bits_robIdx_value;
        output io_exuWriteback_15_bits_fflags;
        output io_exuWriteback_15_bits_wflags;
        output io_exuWriteback_15_bits_vxsat;
        output io_exuWriteback_14_valid;
        output io_exuWriteback_14_bits_data_0;
        output io_exuWriteback_14_bits_robIdx_value;
        output io_exuWriteback_14_bits_fflags;
        output io_exuWriteback_14_bits_wflags;
        output io_exuWriteback_13_valid;
        output io_exuWriteback_13_bits_data_0;
        output io_exuWriteback_13_bits_robIdx_value;
        output io_exuWriteback_13_bits_fflags;
        output io_exuWriteback_13_bits_wflags;
        output io_exuWriteback_13_bits_vxsat;
        output io_exuWriteback_12_valid;
        output io_exuWriteback_12_bits_data_0;
        output io_exuWriteback_12_bits_robIdx_value;
        output io_exuWriteback_12_bits_fflags;
        output io_exuWriteback_12_bits_wflags;
        output io_exuWriteback_11_valid;
        output io_exuWriteback_11_bits_data_0;
        output io_exuWriteback_11_bits_robIdx_value;
        output io_exuWriteback_11_bits_fflags;
        output io_exuWriteback_11_bits_wflags;
        output io_exuWriteback_10_valid;
        output io_exuWriteback_10_bits_data_0;
        output io_exuWriteback_10_bits_robIdx_value;
        output io_exuWriteback_10_bits_fflags;
        output io_exuWriteback_10_bits_wflags;
        output io_exuWriteback_9_valid;
        output io_exuWriteback_9_bits_data_0;
        output io_exuWriteback_9_bits_robIdx_value;
        output io_exuWriteback_9_bits_fflags;
        output io_exuWriteback_9_bits_wflags;
        output io_exuWriteback_8_valid;
        output io_exuWriteback_8_bits_data_0;
        output io_exuWriteback_8_bits_robIdx_value;
        output io_exuWriteback_8_bits_fflags;
        output io_exuWriteback_8_bits_wflags;
        output io_exuWriteback_7_valid;
        output io_exuWriteback_7_bits_data_0;
        output io_exuWriteback_7_bits_robIdx_value;
        output io_exuWriteback_7_bits_debug_isPerfCnt;
        output io_exuWriteback_6_valid;
        output io_exuWriteback_6_bits_data_0;
        output io_exuWriteback_6_bits_robIdx_value;
        output io_exuWriteback_5_valid;
        output io_exuWriteback_5_bits_data_0;
        output io_exuWriteback_5_bits_robIdx_value;
        output io_exuWriteback_5_bits_redirect_valid;
        output io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken;
        output io_exuWriteback_5_bits_fflags;
        output io_exuWriteback_5_bits_wflags;
        output io_exuWriteback_4_valid;
        output io_exuWriteback_4_bits_data_0;
        output io_exuWriteback_4_bits_robIdx_value;
        output io_exuWriteback_3_valid;
        output io_exuWriteback_3_bits_data_0;
        output io_exuWriteback_3_bits_robIdx_value;
        output io_exuWriteback_3_bits_redirect_valid;
        output io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken;
        output io_exuWriteback_2_valid;
        output io_exuWriteback_2_bits_data_0;
        output io_exuWriteback_2_bits_robIdx_value;
        output io_exuWriteback_1_valid;
        output io_exuWriteback_1_bits_data_0;
        output io_exuWriteback_1_bits_robIdx_value;
        output io_exuWriteback_1_bits_redirect_valid;
        output io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken;
        output io_exuWriteback_0_valid;
        output io_exuWriteback_0_bits_data_0;
        output io_exuWriteback_0_bits_robIdx_value;
        output io_writebackNums_0_bits;
        output io_writebackNums_1_bits;
        output io_writebackNums_2_bits;
        output io_writebackNums_3_bits;
        output io_writebackNums_4_bits;
        output io_writebackNums_5_bits;
        output io_writebackNums_6_bits;
        output io_writebackNums_7_bits;
        output io_writebackNums_8_bits;
        output io_writebackNums_9_bits;
        output io_writebackNums_10_bits;
        output io_writebackNums_11_bits;
        output io_writebackNums_12_bits;
        output io_writebackNums_13_bits;
        output io_writebackNums_14_bits;
        output io_writebackNums_15_bits;
        output io_writebackNums_16_bits;
        output io_writebackNums_17_bits;
        output io_writebackNums_18_bits;
        output io_writebackNums_19_bits;
        output io_writebackNums_20_bits;
        output io_writebackNums_21_bits;
        output io_writebackNums_22_bits;
        output io_writebackNums_23_bits;
        output io_writebackNums_24_bits;
        output io_writebackNeedFlush_0;
        output io_writebackNeedFlush_1;
        output io_writebackNeedFlush_2;
        output io_writebackNeedFlush_6;
        output io_writebackNeedFlush_7;
        output io_writebackNeedFlush_8;
        output io_writebackNeedFlush_9;
        output io_writebackNeedFlush_10;
        output io_writebackNeedFlush_11;
        output io_writebackNeedFlush_12;

    endclocking:drv_cb

    clocking mon_cb @(posedge clk);
        `ifdef INTERFACE_ADD_DELAY
            default input #`DEF_SETUP_TIME output #`DEF_HOLD_TIME;
        `endif
        input  io_writeback_24_valid;
        input  io_writeback_24_bits_data_0;
        input  io_writeback_24_bits_pdest;
        input  io_writeback_24_bits_robIdx_flag;
        input  io_writeback_24_bits_robIdx_value;
        input  io_writeback_24_bits_vecWen;
        input  io_writeback_24_bits_v0Wen;
        input  io_writeback_24_bits_vlWen;
        input  io_writeback_24_bits_exceptionVec_0;
        input  io_writeback_24_bits_exceptionVec_1;
        input  io_writeback_24_bits_exceptionVec_2;
        input  io_writeback_24_bits_exceptionVec_3;
        input  io_writeback_24_bits_exceptionVec_4;
        input  io_writeback_24_bits_exceptionVec_5;
        input  io_writeback_24_bits_exceptionVec_6;
        input  io_writeback_24_bits_exceptionVec_7;
        input  io_writeback_24_bits_exceptionVec_8;
        input  io_writeback_24_bits_exceptionVec_9;
        input  io_writeback_24_bits_exceptionVec_10;
        input  io_writeback_24_bits_exceptionVec_11;
        input  io_writeback_24_bits_exceptionVec_12;
        input  io_writeback_24_bits_exceptionVec_13;
        input  io_writeback_24_bits_exceptionVec_14;
        input  io_writeback_24_bits_exceptionVec_15;
        input  io_writeback_24_bits_exceptionVec_16;
        input  io_writeback_24_bits_exceptionVec_17;
        input  io_writeback_24_bits_exceptionVec_18;
        input  io_writeback_24_bits_exceptionVec_19;
        input  io_writeback_24_bits_exceptionVec_20;
        input  io_writeback_24_bits_exceptionVec_21;
        input  io_writeback_24_bits_exceptionVec_22;
        input  io_writeback_24_bits_exceptionVec_23;
        input  io_writeback_24_bits_flushPipe;
        input  io_writeback_24_bits_replay;
        input  io_writeback_24_bits_trigger;
        input  io_writeback_24_bits_vls_vpu_vill;
        input  io_writeback_24_bits_vls_vpu_vma;
        input  io_writeback_24_bits_vls_vpu_vta;
        input  io_writeback_24_bits_vls_vpu_vsew;
        input  io_writeback_24_bits_vls_vpu_vlmul;
        input  io_writeback_24_bits_vls_vpu_specVill;
        input  io_writeback_24_bits_vls_vpu_specVma;
        input  io_writeback_24_bits_vls_vpu_specVta;
        input  io_writeback_24_bits_vls_vpu_specVsew;
        input  io_writeback_24_bits_vls_vpu_specVlmul;
        input  io_writeback_24_bits_vls_vpu_vm;
        input  io_writeback_24_bits_vls_vpu_vstart;
        input  io_writeback_24_bits_vls_vpu_frm;
        input  io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst;
        input  io_writeback_24_bits_vls_vpu_fpu_isFP32Instr;
        input  io_writeback_24_bits_vls_vpu_fpu_isFP64Instr;
        input  io_writeback_24_bits_vls_vpu_fpu_isReduction;
        input  io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2;
        input  io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4;
        input  io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8;
        input  io_writeback_24_bits_vls_vpu_vxrm;
        input  io_writeback_24_bits_vls_vpu_vuopIdx;
        input  io_writeback_24_bits_vls_vpu_lastUop;
        input  io_writeback_24_bits_vls_vpu_vmask;
        input  io_writeback_24_bits_vls_vpu_vl;
        input  io_writeback_24_bits_vls_vpu_nf;
        input  io_writeback_24_bits_vls_vpu_veew;
        input  io_writeback_24_bits_vls_vpu_isReverse;
        input  io_writeback_24_bits_vls_vpu_isExt;
        input  io_writeback_24_bits_vls_vpu_isNarrow;
        input  io_writeback_24_bits_vls_vpu_isDstMask;
        input  io_writeback_24_bits_vls_vpu_isOpMask;
        input  io_writeback_24_bits_vls_vpu_isMove;
        input  io_writeback_24_bits_vls_vpu_isDependOldVd;
        input  io_writeback_24_bits_vls_vpu_isWritePartVd;
        input  io_writeback_24_bits_vls_vpu_isVleff;
        input  io_writeback_24_bits_vls_oldVdPsrc;
        input  io_writeback_24_bits_vls_vdIdx;
        input  io_writeback_24_bits_vls_vdIdxInField;
        input  io_writeback_24_bits_vls_isIndexed;
        input  io_writeback_24_bits_vls_isMasked;
        input  io_writeback_24_bits_vls_isStrided;
        input  io_writeback_24_bits_vls_isWhole;
        input  io_writeback_24_bits_vls_isVecLoad;
        input  io_writeback_24_bits_vls_isVlm;
        input  io_writeback_24_bits_debug_isMMIO;
        input  io_writeback_24_bits_debug_isNCIO;
        input  io_writeback_24_bits_debug_isPerfCnt;
        input  io_writeback_24_bits_debug_paddr;
        input  io_writeback_24_bits_debug_vaddr;
        input  io_writeback_24_bits_debugInfo_eliminatedMove;
        input  io_writeback_24_bits_debugInfo_renameTime;
        input  io_writeback_24_bits_debugInfo_dispatchTime;
        input  io_writeback_24_bits_debugInfo_enqRsTime;
        input  io_writeback_24_bits_debugInfo_selectTime;
        input  io_writeback_24_bits_debugInfo_issueTime;
        input  io_writeback_24_bits_debugInfo_writebackTime;
        input  io_writeback_24_bits_debugInfo_runahead_checkpoint_id;
        input  io_writeback_24_bits_debugInfo_tlbFirstReqTime;
        input  io_writeback_24_bits_debugInfo_tlbRespTime;
        input  io_writeback_24_bits_debug_seqNum;
        input  io_writeback_23_valid;
        input  io_writeback_23_bits_data_0;
        input  io_writeback_23_bits_pdest;
        input  io_writeback_23_bits_robIdx_flag;
        input  io_writeback_23_bits_robIdx_value;
        input  io_writeback_23_bits_vecWen;
        input  io_writeback_23_bits_v0Wen;
        input  io_writeback_23_bits_vlWen;
        input  io_writeback_23_bits_exceptionVec_0;
        input  io_writeback_23_bits_exceptionVec_1;
        input  io_writeback_23_bits_exceptionVec_2;
        input  io_writeback_23_bits_exceptionVec_3;
        input  io_writeback_23_bits_exceptionVec_4;
        input  io_writeback_23_bits_exceptionVec_5;
        input  io_writeback_23_bits_exceptionVec_6;
        input  io_writeback_23_bits_exceptionVec_7;
        input  io_writeback_23_bits_exceptionVec_8;
        input  io_writeback_23_bits_exceptionVec_9;
        input  io_writeback_23_bits_exceptionVec_10;
        input  io_writeback_23_bits_exceptionVec_11;
        input  io_writeback_23_bits_exceptionVec_12;
        input  io_writeback_23_bits_exceptionVec_13;
        input  io_writeback_23_bits_exceptionVec_14;
        input  io_writeback_23_bits_exceptionVec_15;
        input  io_writeback_23_bits_exceptionVec_16;
        input  io_writeback_23_bits_exceptionVec_17;
        input  io_writeback_23_bits_exceptionVec_18;
        input  io_writeback_23_bits_exceptionVec_19;
        input  io_writeback_23_bits_exceptionVec_20;
        input  io_writeback_23_bits_exceptionVec_21;
        input  io_writeback_23_bits_exceptionVec_22;
        input  io_writeback_23_bits_exceptionVec_23;
        input  io_writeback_23_bits_flushPipe;
        input  io_writeback_23_bits_replay;
        input  io_writeback_23_bits_trigger;
        input  io_writeback_23_bits_vls_vpu_vill;
        input  io_writeback_23_bits_vls_vpu_vma;
        input  io_writeback_23_bits_vls_vpu_vta;
        input  io_writeback_23_bits_vls_vpu_vsew;
        input  io_writeback_23_bits_vls_vpu_vlmul;
        input  io_writeback_23_bits_vls_vpu_specVill;
        input  io_writeback_23_bits_vls_vpu_specVma;
        input  io_writeback_23_bits_vls_vpu_specVta;
        input  io_writeback_23_bits_vls_vpu_specVsew;
        input  io_writeback_23_bits_vls_vpu_specVlmul;
        input  io_writeback_23_bits_vls_vpu_vm;
        input  io_writeback_23_bits_vls_vpu_vstart;
        input  io_writeback_23_bits_vls_vpu_frm;
        input  io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst;
        input  io_writeback_23_bits_vls_vpu_fpu_isFP32Instr;
        input  io_writeback_23_bits_vls_vpu_fpu_isFP64Instr;
        input  io_writeback_23_bits_vls_vpu_fpu_isReduction;
        input  io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2;
        input  io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4;
        input  io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8;
        input  io_writeback_23_bits_vls_vpu_vxrm;
        input  io_writeback_23_bits_vls_vpu_vuopIdx;
        input  io_writeback_23_bits_vls_vpu_lastUop;
        input  io_writeback_23_bits_vls_vpu_vmask;
        input  io_writeback_23_bits_vls_vpu_vl;
        input  io_writeback_23_bits_vls_vpu_nf;
        input  io_writeback_23_bits_vls_vpu_veew;
        input  io_writeback_23_bits_vls_vpu_isReverse;
        input  io_writeback_23_bits_vls_vpu_isExt;
        input  io_writeback_23_bits_vls_vpu_isNarrow;
        input  io_writeback_23_bits_vls_vpu_isDstMask;
        input  io_writeback_23_bits_vls_vpu_isOpMask;
        input  io_writeback_23_bits_vls_vpu_isMove;
        input  io_writeback_23_bits_vls_vpu_isDependOldVd;
        input  io_writeback_23_bits_vls_vpu_isWritePartVd;
        input  io_writeback_23_bits_vls_vpu_isVleff;
        input  io_writeback_23_bits_vls_oldVdPsrc;
        input  io_writeback_23_bits_vls_vdIdx;
        input  io_writeback_23_bits_vls_vdIdxInField;
        input  io_writeback_23_bits_vls_isIndexed;
        input  io_writeback_23_bits_vls_isMasked;
        input  io_writeback_23_bits_vls_isStrided;
        input  io_writeback_23_bits_vls_isWhole;
        input  io_writeback_23_bits_vls_isVecLoad;
        input  io_writeback_23_bits_vls_isVlm;
        input  io_writeback_23_bits_debug_isMMIO;
        input  io_writeback_23_bits_debug_isNCIO;
        input  io_writeback_23_bits_debug_isPerfCnt;
        input  io_writeback_23_bits_debug_paddr;
        input  io_writeback_23_bits_debug_vaddr;
        input  io_writeback_23_bits_debugInfo_eliminatedMove;
        input  io_writeback_23_bits_debugInfo_renameTime;
        input  io_writeback_23_bits_debugInfo_dispatchTime;
        input  io_writeback_23_bits_debugInfo_enqRsTime;
        input  io_writeback_23_bits_debugInfo_selectTime;
        input  io_writeback_23_bits_debugInfo_issueTime;
        input  io_writeback_23_bits_debugInfo_writebackTime;
        input  io_writeback_23_bits_debugInfo_runahead_checkpoint_id;
        input  io_writeback_23_bits_debugInfo_tlbFirstReqTime;
        input  io_writeback_23_bits_debugInfo_tlbRespTime;
        input  io_writeback_23_bits_debug_seqNum;
        input  io_writeback_22_valid;
        input  io_writeback_22_bits_data_0;
        input  io_writeback_22_bits_pdest;
        input  io_writeback_22_bits_robIdx_flag;
        input  io_writeback_22_bits_robIdx_value;
        input  io_writeback_22_bits_intWen;
        input  io_writeback_22_bits_fpWen;
        input  io_writeback_22_bits_exceptionVec_0;
        input  io_writeback_22_bits_exceptionVec_1;
        input  io_writeback_22_bits_exceptionVec_2;
        input  io_writeback_22_bits_exceptionVec_3;
        input  io_writeback_22_bits_exceptionVec_4;
        input  io_writeback_22_bits_exceptionVec_5;
        input  io_writeback_22_bits_exceptionVec_6;
        input  io_writeback_22_bits_exceptionVec_7;
        input  io_writeback_22_bits_exceptionVec_8;
        input  io_writeback_22_bits_exceptionVec_9;
        input  io_writeback_22_bits_exceptionVec_10;
        input  io_writeback_22_bits_exceptionVec_11;
        input  io_writeback_22_bits_exceptionVec_12;
        input  io_writeback_22_bits_exceptionVec_13;
        input  io_writeback_22_bits_exceptionVec_14;
        input  io_writeback_22_bits_exceptionVec_15;
        input  io_writeback_22_bits_exceptionVec_16;
        input  io_writeback_22_bits_exceptionVec_17;
        input  io_writeback_22_bits_exceptionVec_18;
        input  io_writeback_22_bits_exceptionVec_19;
        input  io_writeback_22_bits_exceptionVec_20;
        input  io_writeback_22_bits_exceptionVec_21;
        input  io_writeback_22_bits_exceptionVec_22;
        input  io_writeback_22_bits_exceptionVec_23;
        input  io_writeback_22_bits_flushPipe;
        input  io_writeback_22_bits_replay;
        input  io_writeback_22_bits_lqIdx_flag;
        input  io_writeback_22_bits_lqIdx_value;
        input  io_writeback_22_bits_trigger;
        input  io_writeback_22_bits_predecodeInfo_valid;
        input  io_writeback_22_bits_predecodeInfo_isRVC;
        input  io_writeback_22_bits_predecodeInfo_brType;
        input  io_writeback_22_bits_predecodeInfo_isCall;
        input  io_writeback_22_bits_predecodeInfo_isRet;
        input  io_writeback_22_bits_debug_isMMIO;
        input  io_writeback_22_bits_debug_isNCIO;
        input  io_writeback_22_bits_debug_isPerfCnt;
        input  io_writeback_22_bits_debug_paddr;
        input  io_writeback_22_bits_debug_vaddr;
        input  io_writeback_22_bits_debugInfo_eliminatedMove;
        input  io_writeback_22_bits_debugInfo_renameTime;
        input  io_writeback_22_bits_debugInfo_dispatchTime;
        input  io_writeback_22_bits_debugInfo_enqRsTime;
        input  io_writeback_22_bits_debugInfo_selectTime;
        input  io_writeback_22_bits_debugInfo_issueTime;
        input  io_writeback_22_bits_debugInfo_writebackTime;
        input  io_writeback_22_bits_debugInfo_runahead_checkpoint_id;
        input  io_writeback_22_bits_debugInfo_tlbFirstReqTime;
        input  io_writeback_22_bits_debugInfo_tlbRespTime;
        input  io_writeback_22_bits_debug_seqNum;
        input  io_writeback_21_valid;
        input  io_writeback_21_bits_data_0;
        input  io_writeback_21_bits_pdest;
        input  io_writeback_21_bits_robIdx_flag;
        input  io_writeback_21_bits_robIdx_value;
        input  io_writeback_21_bits_intWen;
        input  io_writeback_21_bits_fpWen;
        input  io_writeback_21_bits_exceptionVec_0;
        input  io_writeback_21_bits_exceptionVec_1;
        input  io_writeback_21_bits_exceptionVec_2;
        input  io_writeback_21_bits_exceptionVec_3;
        input  io_writeback_21_bits_exceptionVec_4;
        input  io_writeback_21_bits_exceptionVec_5;
        input  io_writeback_21_bits_exceptionVec_6;
        input  io_writeback_21_bits_exceptionVec_7;
        input  io_writeback_21_bits_exceptionVec_8;
        input  io_writeback_21_bits_exceptionVec_9;
        input  io_writeback_21_bits_exceptionVec_10;
        input  io_writeback_21_bits_exceptionVec_11;
        input  io_writeback_21_bits_exceptionVec_12;
        input  io_writeback_21_bits_exceptionVec_13;
        input  io_writeback_21_bits_exceptionVec_14;
        input  io_writeback_21_bits_exceptionVec_15;
        input  io_writeback_21_bits_exceptionVec_16;
        input  io_writeback_21_bits_exceptionVec_17;
        input  io_writeback_21_bits_exceptionVec_18;
        input  io_writeback_21_bits_exceptionVec_19;
        input  io_writeback_21_bits_exceptionVec_20;
        input  io_writeback_21_bits_exceptionVec_21;
        input  io_writeback_21_bits_exceptionVec_22;
        input  io_writeback_21_bits_exceptionVec_23;
        input  io_writeback_21_bits_flushPipe;
        input  io_writeback_21_bits_replay;
        input  io_writeback_21_bits_lqIdx_flag;
        input  io_writeback_21_bits_lqIdx_value;
        input  io_writeback_21_bits_trigger;
        input  io_writeback_21_bits_predecodeInfo_valid;
        input  io_writeback_21_bits_predecodeInfo_isRVC;
        input  io_writeback_21_bits_predecodeInfo_brType;
        input  io_writeback_21_bits_predecodeInfo_isCall;
        input  io_writeback_21_bits_predecodeInfo_isRet;
        input  io_writeback_21_bits_debug_isMMIO;
        input  io_writeback_21_bits_debug_isNCIO;
        input  io_writeback_21_bits_debug_isPerfCnt;
        input  io_writeback_21_bits_debug_paddr;
        input  io_writeback_21_bits_debug_vaddr;
        input  io_writeback_21_bits_debugInfo_eliminatedMove;
        input  io_writeback_21_bits_debugInfo_renameTime;
        input  io_writeback_21_bits_debugInfo_dispatchTime;
        input  io_writeback_21_bits_debugInfo_enqRsTime;
        input  io_writeback_21_bits_debugInfo_selectTime;
        input  io_writeback_21_bits_debugInfo_issueTime;
        input  io_writeback_21_bits_debugInfo_writebackTime;
        input  io_writeback_21_bits_debugInfo_runahead_checkpoint_id;
        input  io_writeback_21_bits_debugInfo_tlbFirstReqTime;
        input  io_writeback_21_bits_debugInfo_tlbRespTime;
        input  io_writeback_21_bits_debug_seqNum;
        input  io_writeback_20_valid;
        input  io_writeback_20_bits_data_0;
        input  io_writeback_20_bits_pdest;
        input  io_writeback_20_bits_robIdx_flag;
        input  io_writeback_20_bits_robIdx_value;
        input  io_writeback_20_bits_intWen;
        input  io_writeback_20_bits_fpWen;
        input  io_writeback_20_bits_exceptionVec_0;
        input  io_writeback_20_bits_exceptionVec_1;
        input  io_writeback_20_bits_exceptionVec_2;
        input  io_writeback_20_bits_exceptionVec_3;
        input  io_writeback_20_bits_exceptionVec_4;
        input  io_writeback_20_bits_exceptionVec_5;
        input  io_writeback_20_bits_exceptionVec_6;
        input  io_writeback_20_bits_exceptionVec_7;
        input  io_writeback_20_bits_exceptionVec_8;
        input  io_writeback_20_bits_exceptionVec_9;
        input  io_writeback_20_bits_exceptionVec_10;
        input  io_writeback_20_bits_exceptionVec_11;
        input  io_writeback_20_bits_exceptionVec_12;
        input  io_writeback_20_bits_exceptionVec_13;
        input  io_writeback_20_bits_exceptionVec_14;
        input  io_writeback_20_bits_exceptionVec_15;
        input  io_writeback_20_bits_exceptionVec_16;
        input  io_writeback_20_bits_exceptionVec_17;
        input  io_writeback_20_bits_exceptionVec_18;
        input  io_writeback_20_bits_exceptionVec_19;
        input  io_writeback_20_bits_exceptionVec_20;
        input  io_writeback_20_bits_exceptionVec_21;
        input  io_writeback_20_bits_exceptionVec_22;
        input  io_writeback_20_bits_exceptionVec_23;
        input  io_writeback_20_bits_flushPipe;
        input  io_writeback_20_bits_replay;
        input  io_writeback_20_bits_lqIdx_flag;
        input  io_writeback_20_bits_lqIdx_value;
        input  io_writeback_20_bits_trigger;
        input  io_writeback_20_bits_predecodeInfo_valid;
        input  io_writeback_20_bits_predecodeInfo_isRVC;
        input  io_writeback_20_bits_predecodeInfo_brType;
        input  io_writeback_20_bits_predecodeInfo_isCall;
        input  io_writeback_20_bits_predecodeInfo_isRet;
        input  io_writeback_20_bits_debug_isMMIO;
        input  io_writeback_20_bits_debug_isNCIO;
        input  io_writeback_20_bits_debug_isPerfCnt;
        input  io_writeback_20_bits_debug_paddr;
        input  io_writeback_20_bits_debug_vaddr;
        input  io_writeback_20_bits_debugInfo_eliminatedMove;
        input  io_writeback_20_bits_debugInfo_renameTime;
        input  io_writeback_20_bits_debugInfo_dispatchTime;
        input  io_writeback_20_bits_debugInfo_enqRsTime;
        input  io_writeback_20_bits_debugInfo_selectTime;
        input  io_writeback_20_bits_debugInfo_issueTime;
        input  io_writeback_20_bits_debugInfo_writebackTime;
        input  io_writeback_20_bits_debugInfo_runahead_checkpoint_id;
        input  io_writeback_20_bits_debugInfo_tlbFirstReqTime;
        input  io_writeback_20_bits_debugInfo_tlbRespTime;
        input  io_writeback_20_bits_debug_seqNum;
        input  io_writeback_19_valid;
        input  io_writeback_19_bits_data_0;
        input  io_writeback_19_bits_pdest;
        input  io_writeback_19_bits_robIdx_flag;
        input  io_writeback_19_bits_robIdx_value;
        input  io_writeback_19_bits_intWen;
        input  io_writeback_19_bits_exceptionVec_0;
        input  io_writeback_19_bits_exceptionVec_1;
        input  io_writeback_19_bits_exceptionVec_2;
        input  io_writeback_19_bits_exceptionVec_3;
        input  io_writeback_19_bits_exceptionVec_4;
        input  io_writeback_19_bits_exceptionVec_5;
        input  io_writeback_19_bits_exceptionVec_6;
        input  io_writeback_19_bits_exceptionVec_7;
        input  io_writeback_19_bits_exceptionVec_8;
        input  io_writeback_19_bits_exceptionVec_9;
        input  io_writeback_19_bits_exceptionVec_10;
        input  io_writeback_19_bits_exceptionVec_11;
        input  io_writeback_19_bits_exceptionVec_12;
        input  io_writeback_19_bits_exceptionVec_13;
        input  io_writeback_19_bits_exceptionVec_14;
        input  io_writeback_19_bits_exceptionVec_15;
        input  io_writeback_19_bits_exceptionVec_16;
        input  io_writeback_19_bits_exceptionVec_17;
        input  io_writeback_19_bits_exceptionVec_18;
        input  io_writeback_19_bits_exceptionVec_19;
        input  io_writeback_19_bits_exceptionVec_20;
        input  io_writeback_19_bits_exceptionVec_21;
        input  io_writeback_19_bits_exceptionVec_22;
        input  io_writeback_19_bits_exceptionVec_23;
        input  io_writeback_19_bits_flushPipe;
        input  io_writeback_19_bits_sqIdx_flag;
        input  io_writeback_19_bits_sqIdx_value;
        input  io_writeback_19_bits_trigger;
        input  io_writeback_19_bits_debug_isMMIO;
        input  io_writeback_19_bits_debug_isNCIO;
        input  io_writeback_19_bits_debug_isPerfCnt;
        input  io_writeback_19_bits_debug_paddr;
        input  io_writeback_19_bits_debug_vaddr;
        input  io_writeback_19_bits_debugInfo_eliminatedMove;
        input  io_writeback_19_bits_debugInfo_renameTime;
        input  io_writeback_19_bits_debugInfo_dispatchTime;
        input  io_writeback_19_bits_debugInfo_enqRsTime;
        input  io_writeback_19_bits_debugInfo_selectTime;
        input  io_writeback_19_bits_debugInfo_issueTime;
        input  io_writeback_19_bits_debugInfo_writebackTime;
        input  io_writeback_19_bits_debugInfo_runahead_checkpoint_id;
        input  io_writeback_19_bits_debugInfo_tlbFirstReqTime;
        input  io_writeback_19_bits_debugInfo_tlbRespTime;
        input  io_writeback_19_bits_debug_seqNum;
        input  io_writeback_18_valid;
        input  io_writeback_18_bits_data_0;
        input  io_writeback_18_bits_pdest;
        input  io_writeback_18_bits_robIdx_flag;
        input  io_writeback_18_bits_robIdx_value;
        input  io_writeback_18_bits_intWen;
        input  io_writeback_18_bits_exceptionVec_0;
        input  io_writeback_18_bits_exceptionVec_1;
        input  io_writeback_18_bits_exceptionVec_2;
        input  io_writeback_18_bits_exceptionVec_3;
        input  io_writeback_18_bits_exceptionVec_4;
        input  io_writeback_18_bits_exceptionVec_5;
        input  io_writeback_18_bits_exceptionVec_6;
        input  io_writeback_18_bits_exceptionVec_7;
        input  io_writeback_18_bits_exceptionVec_8;
        input  io_writeback_18_bits_exceptionVec_9;
        input  io_writeback_18_bits_exceptionVec_10;
        input  io_writeback_18_bits_exceptionVec_11;
        input  io_writeback_18_bits_exceptionVec_12;
        input  io_writeback_18_bits_exceptionVec_13;
        input  io_writeback_18_bits_exceptionVec_14;
        input  io_writeback_18_bits_exceptionVec_15;
        input  io_writeback_18_bits_exceptionVec_16;
        input  io_writeback_18_bits_exceptionVec_17;
        input  io_writeback_18_bits_exceptionVec_18;
        input  io_writeback_18_bits_exceptionVec_19;
        input  io_writeback_18_bits_exceptionVec_20;
        input  io_writeback_18_bits_exceptionVec_21;
        input  io_writeback_18_bits_exceptionVec_22;
        input  io_writeback_18_bits_exceptionVec_23;
        input  io_writeback_18_bits_flushPipe;
        input  io_writeback_18_bits_sqIdx_flag;
        input  io_writeback_18_bits_sqIdx_value;
        input  io_writeback_18_bits_trigger;
        input  io_writeback_18_bits_debug_isMMIO;
        input  io_writeback_18_bits_debug_isNCIO;
        input  io_writeback_18_bits_debug_isPerfCnt;
        input  io_writeback_18_bits_debug_paddr;
        input  io_writeback_18_bits_debug_vaddr;
        input  io_writeback_18_bits_debugInfo_eliminatedMove;
        input  io_writeback_18_bits_debugInfo_renameTime;
        input  io_writeback_18_bits_debugInfo_dispatchTime;
        input  io_writeback_18_bits_debugInfo_enqRsTime;
        input  io_writeback_18_bits_debugInfo_selectTime;
        input  io_writeback_18_bits_debugInfo_issueTime;
        input  io_writeback_18_bits_debugInfo_writebackTime;
        input  io_writeback_18_bits_debugInfo_runahead_checkpoint_id;
        input  io_writeback_18_bits_debugInfo_tlbFirstReqTime;
        input  io_writeback_18_bits_debugInfo_tlbRespTime;
        input  io_writeback_18_bits_debug_seqNum;
        input  io_writeback_17_valid;
        input  io_writeback_17_bits_data_0;
        input  io_writeback_17_bits_data_1;
        input  io_writeback_17_bits_data_2;
        input  io_writeback_17_bits_pdest;
        input  io_writeback_17_bits_robIdx_flag;
        input  io_writeback_17_bits_robIdx_value;
        input  io_writeback_17_bits_vecWen;
        input  io_writeback_17_bits_v0Wen;
        input  io_writeback_17_bits_fflags;
        input  io_writeback_17_bits_wflags;
        input  io_writeback_17_bits_debugInfo_eliminatedMove;
        input  io_writeback_17_bits_debugInfo_renameTime;
        input  io_writeback_17_bits_debugInfo_dispatchTime;
        input  io_writeback_17_bits_debugInfo_enqRsTime;
        input  io_writeback_17_bits_debugInfo_selectTime;
        input  io_writeback_17_bits_debugInfo_issueTime;
        input  io_writeback_17_bits_debugInfo_writebackTime;
        input  io_writeback_17_bits_debugInfo_runahead_checkpoint_id;
        input  io_writeback_17_bits_debugInfo_tlbFirstReqTime;
        input  io_writeback_17_bits_debugInfo_tlbRespTime;
        input  io_writeback_17_bits_debug_seqNum;
        input  io_writeback_16_valid;
        input  io_writeback_16_bits_data_0;
        input  io_writeback_16_bits_data_1;
        input  io_writeback_16_bits_data_2;
        input  io_writeback_16_bits_data_3;
        input  io_writeback_16_bits_pdest;
        input  io_writeback_16_bits_robIdx_flag;
        input  io_writeback_16_bits_robIdx_value;
        input  io_writeback_16_bits_fpWen;
        input  io_writeback_16_bits_vecWen;
        input  io_writeback_16_bits_v0Wen;
        input  io_writeback_16_bits_fflags;
        input  io_writeback_16_bits_wflags;
        input  io_writeback_16_bits_debugInfo_eliminatedMove;
        input  io_writeback_16_bits_debugInfo_renameTime;
        input  io_writeback_16_bits_debugInfo_dispatchTime;
        input  io_writeback_16_bits_debugInfo_enqRsTime;
        input  io_writeback_16_bits_debugInfo_selectTime;
        input  io_writeback_16_bits_debugInfo_issueTime;
        input  io_writeback_16_bits_debugInfo_writebackTime;
        input  io_writeback_16_bits_debugInfo_runahead_checkpoint_id;
        input  io_writeback_16_bits_debugInfo_tlbFirstReqTime;
        input  io_writeback_16_bits_debugInfo_tlbRespTime;
        input  io_writeback_16_bits_debug_seqNum;
        input  io_writeback_15_valid;
        input  io_writeback_15_bits_data_0;
        input  io_writeback_15_bits_data_1;
        input  io_writeback_15_bits_data_2;
        input  io_writeback_15_bits_pdest;
        input  io_writeback_15_bits_robIdx_flag;
        input  io_writeback_15_bits_robIdx_value;
        input  io_writeback_15_bits_vecWen;
        input  io_writeback_15_bits_v0Wen;
        input  io_writeback_15_bits_fflags;
        input  io_writeback_15_bits_wflags;
        input  io_writeback_15_bits_vxsat;
        input  io_writeback_15_bits_debugInfo_eliminatedMove;
        input  io_writeback_15_bits_debugInfo_renameTime;
        input  io_writeback_15_bits_debugInfo_dispatchTime;
        input  io_writeback_15_bits_debugInfo_enqRsTime;
        input  io_writeback_15_bits_debugInfo_selectTime;
        input  io_writeback_15_bits_debugInfo_issueTime;
        input  io_writeback_15_bits_debugInfo_writebackTime;
        input  io_writeback_15_bits_debugInfo_runahead_checkpoint_id;
        input  io_writeback_15_bits_debugInfo_tlbFirstReqTime;
        input  io_writeback_15_bits_debugInfo_tlbRespTime;
        input  io_writeback_15_bits_debug_seqNum;
        input  io_writeback_14_valid;
        input  io_writeback_14_bits_data_0;
        input  io_writeback_14_bits_data_1;
        input  io_writeback_14_bits_data_2;
        input  io_writeback_14_bits_data_3;
        input  io_writeback_14_bits_data_4;
        input  io_writeback_14_bits_data_5;
        input  io_writeback_14_bits_pdest;
        input  io_writeback_14_bits_robIdx_flag;
        input  io_writeback_14_bits_robIdx_value;
        input  io_writeback_14_bits_intWen;
        input  io_writeback_14_bits_fpWen;
        input  io_writeback_14_bits_vecWen;
        input  io_writeback_14_bits_v0Wen;
        input  io_writeback_14_bits_vlWen;
        input  io_writeback_14_bits_fflags;
        input  io_writeback_14_bits_wflags;
        input  io_writeback_14_bits_exceptionVec_2;
        input  io_writeback_14_bits_debugInfo_eliminatedMove;
        input  io_writeback_14_bits_debugInfo_renameTime;
        input  io_writeback_14_bits_debugInfo_dispatchTime;
        input  io_writeback_14_bits_debugInfo_enqRsTime;
        input  io_writeback_14_bits_debugInfo_selectTime;
        input  io_writeback_14_bits_debugInfo_issueTime;
        input  io_writeback_14_bits_debugInfo_writebackTime;
        input  io_writeback_14_bits_debugInfo_runahead_checkpoint_id;
        input  io_writeback_14_bits_debugInfo_tlbFirstReqTime;
        input  io_writeback_14_bits_debugInfo_tlbRespTime;
        input  io_writeback_14_bits_debug_seqNum;
        input  io_writeback_13_valid;
        input  io_writeback_13_bits_data_0;
        input  io_writeback_13_bits_data_1;
        input  io_writeback_13_bits_data_2;
        input  io_writeback_13_bits_pdest;
        input  io_writeback_13_bits_robIdx_flag;
        input  io_writeback_13_bits_robIdx_value;
        input  io_writeback_13_bits_vecWen;
        input  io_writeback_13_bits_v0Wen;
        input  io_writeback_13_bits_fflags;
        input  io_writeback_13_bits_wflags;
        input  io_writeback_13_bits_vxsat;
        input  io_writeback_13_bits_exceptionVec_2;
        input  io_writeback_13_bits_debugInfo_eliminatedMove;
        input  io_writeback_13_bits_debugInfo_renameTime;
        input  io_writeback_13_bits_debugInfo_dispatchTime;
        input  io_writeback_13_bits_debugInfo_enqRsTime;
        input  io_writeback_13_bits_debugInfo_selectTime;
        input  io_writeback_13_bits_debugInfo_issueTime;
        input  io_writeback_13_bits_debugInfo_writebackTime;
        input  io_writeback_13_bits_debugInfo_runahead_checkpoint_id;
        input  io_writeback_13_bits_debugInfo_tlbFirstReqTime;
        input  io_writeback_13_bits_debugInfo_tlbRespTime;
        input  io_writeback_13_bits_debug_seqNum;
        input  io_writeback_7_valid;
        input  io_writeback_7_bits_data_0;
        input  io_writeback_7_bits_data_1;
        input  io_writeback_7_bits_pdest;
        input  io_writeback_7_bits_robIdx_flag;
        input  io_writeback_7_bits_robIdx_value;
        input  io_writeback_7_bits_intWen;
        input  io_writeback_7_bits_redirect_valid;
        input  io_writeback_7_bits_redirect_bits_isRVC;
        input  io_writeback_7_bits_redirect_bits_robIdx_flag;
        input  io_writeback_7_bits_redirect_bits_robIdx_value;
        input  io_writeback_7_bits_redirect_bits_ftqIdx_flag;
        input  io_writeback_7_bits_redirect_bits_ftqIdx_value;
        input  io_writeback_7_bits_redirect_bits_ftqOffset;
        input  io_writeback_7_bits_redirect_bits_level;
        input  io_writeback_7_bits_redirect_bits_interrupt;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_pc;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_ssp;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_sctr;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_ghr;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_target;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_taken;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_shift;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF;
        input  io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF;
        input  io_writeback_7_bits_redirect_bits_fullTarget;
        input  io_writeback_7_bits_redirect_bits_stFtqIdx_flag;
        input  io_writeback_7_bits_redirect_bits_stFtqIdx_value;
        input  io_writeback_7_bits_redirect_bits_stFtqOffset;
        input  io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id;
        input  io_writeback_7_bits_redirect_bits_debugIsCtrl;
        input  io_writeback_7_bits_redirect_bits_debugIsMemVio;
        input  io_writeback_7_bits_exceptionVec_2;
        input  io_writeback_7_bits_exceptionVec_3;
        input  io_writeback_7_bits_exceptionVec_8;
        input  io_writeback_7_bits_exceptionVec_9;
        input  io_writeback_7_bits_exceptionVec_10;
        input  io_writeback_7_bits_exceptionVec_11;
        input  io_writeback_7_bits_exceptionVec_22;
        input  io_writeback_7_bits_flushPipe;
        input  io_writeback_7_bits_predecodeInfo_valid;
        input  io_writeback_7_bits_predecodeInfo_isRVC;
        input  io_writeback_7_bits_predecodeInfo_brType;
        input  io_writeback_7_bits_predecodeInfo_isCall;
        input  io_writeback_7_bits_predecodeInfo_isRet;
        input  io_writeback_7_bits_debug_isPerfCnt;
        input  io_writeback_7_bits_debugInfo_eliminatedMove;
        input  io_writeback_7_bits_debugInfo_renameTime;
        input  io_writeback_7_bits_debugInfo_dispatchTime;
        input  io_writeback_7_bits_debugInfo_enqRsTime;
        input  io_writeback_7_bits_debugInfo_selectTime;
        input  io_writeback_7_bits_debugInfo_issueTime;
        input  io_writeback_7_bits_debugInfo_writebackTime;
        input  io_writeback_7_bits_debugInfo_runahead_checkpoint_id;
        input  io_writeback_7_bits_debugInfo_tlbFirstReqTime;
        input  io_writeback_7_bits_debugInfo_tlbRespTime;
        input  io_writeback_7_bits_debug_seqNum;
        input  io_writeback_5_valid;
        input  io_writeback_5_bits_redirect_valid;
        input  io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred;
        input  io_writeback_3_valid;
        input  io_writeback_3_bits_redirect_valid;
        input  io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred;
        input  io_writeback_1_valid;
        input  io_writeback_1_bits_redirect_valid;
        input  io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred;
        input  io_exuWriteback_26_valid;
        input  io_exuWriteback_26_bits_robIdx_value;
        input  io_exuWriteback_25_valid;
        input  io_exuWriteback_25_bits_robIdx_value;
        input  io_exuWriteback_24_valid;
        input  io_exuWriteback_24_bits_data_0;
        input  io_exuWriteback_24_bits_pdest;
        input  io_exuWriteback_24_bits_robIdx_value;
        input  io_exuWriteback_24_bits_vecWen;
        input  io_exuWriteback_24_bits_v0Wen;
        input  io_exuWriteback_24_bits_vls_vdIdx;
        input  io_exuWriteback_24_bits_debug_isMMIO;
        input  io_exuWriteback_24_bits_debug_isNCIO;
        input  io_exuWriteback_24_bits_debug_isPerfCnt;
        input  io_exuWriteback_24_bits_debug_paddr;
        input  io_exuWriteback_23_valid;
        input  io_exuWriteback_23_bits_data_0;
        input  io_exuWriteback_23_bits_pdest;
        input  io_exuWriteback_23_bits_robIdx_value;
        input  io_exuWriteback_23_bits_vecWen;
        input  io_exuWriteback_23_bits_v0Wen;
        input  io_exuWriteback_23_bits_vls_vdIdx;
        input  io_exuWriteback_23_bits_debug_isMMIO;
        input  io_exuWriteback_23_bits_debug_isNCIO;
        input  io_exuWriteback_23_bits_debug_isPerfCnt;
        input  io_exuWriteback_23_bits_debug_paddr;
        input  io_exuWriteback_22_valid;
        input  io_exuWriteback_22_bits_data_0;
        input  io_exuWriteback_22_bits_robIdx_value;
        input  io_exuWriteback_22_bits_lqIdx_value;
        input  io_exuWriteback_22_bits_debug_isMMIO;
        input  io_exuWriteback_22_bits_debug_isNCIO;
        input  io_exuWriteback_22_bits_debug_isPerfCnt;
        input  io_exuWriteback_22_bits_debug_paddr;
        input  io_exuWriteback_21_valid;
        input  io_exuWriteback_21_bits_data_0;
        input  io_exuWriteback_21_bits_robIdx_value;
        input  io_exuWriteback_21_bits_lqIdx_value;
        input  io_exuWriteback_21_bits_debug_isMMIO;
        input  io_exuWriteback_21_bits_debug_isNCIO;
        input  io_exuWriteback_21_bits_debug_isPerfCnt;
        input  io_exuWriteback_21_bits_debug_paddr;
        input  io_exuWriteback_20_valid;
        input  io_exuWriteback_20_bits_data_0;
        input  io_exuWriteback_20_bits_robIdx_value;
        input  io_exuWriteback_20_bits_lqIdx_value;
        input  io_exuWriteback_20_bits_debug_isMMIO;
        input  io_exuWriteback_20_bits_debug_isNCIO;
        input  io_exuWriteback_20_bits_debug_isPerfCnt;
        input  io_exuWriteback_20_bits_debug_paddr;
        input  io_exuWriteback_19_valid;
        input  io_exuWriteback_19_bits_data_0;
        input  io_exuWriteback_19_bits_robIdx_value;
        input  io_exuWriteback_19_bits_sqIdx_value;
        input  io_exuWriteback_19_bits_debug_isMMIO;
        input  io_exuWriteback_19_bits_debug_isNCIO;
        input  io_exuWriteback_19_bits_debug_isPerfCnt;
        input  io_exuWriteback_19_bits_debug_paddr;
        input  io_exuWriteback_18_valid;
        input  io_exuWriteback_18_bits_data_0;
        input  io_exuWriteback_18_bits_robIdx_value;
        input  io_exuWriteback_18_bits_sqIdx_value;
        input  io_exuWriteback_18_bits_debug_isMMIO;
        input  io_exuWriteback_18_bits_debug_isNCIO;
        input  io_exuWriteback_18_bits_debug_isPerfCnt;
        input  io_exuWriteback_18_bits_debug_paddr;
        input  io_exuWriteback_17_valid;
        input  io_exuWriteback_17_bits_data_0;
        input  io_exuWriteback_17_bits_robIdx_value;
        input  io_exuWriteback_17_bits_fflags;
        input  io_exuWriteback_17_bits_wflags;
        input  io_exuWriteback_16_valid;
        input  io_exuWriteback_16_bits_data_0;
        input  io_exuWriteback_16_bits_robIdx_value;
        input  io_exuWriteback_16_bits_fflags;
        input  io_exuWriteback_16_bits_wflags;
        input  io_exuWriteback_15_valid;
        input  io_exuWriteback_15_bits_data_0;
        input  io_exuWriteback_15_bits_robIdx_value;
        input  io_exuWriteback_15_bits_fflags;
        input  io_exuWriteback_15_bits_wflags;
        input  io_exuWriteback_15_bits_vxsat;
        input  io_exuWriteback_14_valid;
        input  io_exuWriteback_14_bits_data_0;
        input  io_exuWriteback_14_bits_robIdx_value;
        input  io_exuWriteback_14_bits_fflags;
        input  io_exuWriteback_14_bits_wflags;
        input  io_exuWriteback_13_valid;
        input  io_exuWriteback_13_bits_data_0;
        input  io_exuWriteback_13_bits_robIdx_value;
        input  io_exuWriteback_13_bits_fflags;
        input  io_exuWriteback_13_bits_wflags;
        input  io_exuWriteback_13_bits_vxsat;
        input  io_exuWriteback_12_valid;
        input  io_exuWriteback_12_bits_data_0;
        input  io_exuWriteback_12_bits_robIdx_value;
        input  io_exuWriteback_12_bits_fflags;
        input  io_exuWriteback_12_bits_wflags;
        input  io_exuWriteback_11_valid;
        input  io_exuWriteback_11_bits_data_0;
        input  io_exuWriteback_11_bits_robIdx_value;
        input  io_exuWriteback_11_bits_fflags;
        input  io_exuWriteback_11_bits_wflags;
        input  io_exuWriteback_10_valid;
        input  io_exuWriteback_10_bits_data_0;
        input  io_exuWriteback_10_bits_robIdx_value;
        input  io_exuWriteback_10_bits_fflags;
        input  io_exuWriteback_10_bits_wflags;
        input  io_exuWriteback_9_valid;
        input  io_exuWriteback_9_bits_data_0;
        input  io_exuWriteback_9_bits_robIdx_value;
        input  io_exuWriteback_9_bits_fflags;
        input  io_exuWriteback_9_bits_wflags;
        input  io_exuWriteback_8_valid;
        input  io_exuWriteback_8_bits_data_0;
        input  io_exuWriteback_8_bits_robIdx_value;
        input  io_exuWriteback_8_bits_fflags;
        input  io_exuWriteback_8_bits_wflags;
        input  io_exuWriteback_7_valid;
        input  io_exuWriteback_7_bits_data_0;
        input  io_exuWriteback_7_bits_robIdx_value;
        input  io_exuWriteback_7_bits_debug_isPerfCnt;
        input  io_exuWriteback_6_valid;
        input  io_exuWriteback_6_bits_data_0;
        input  io_exuWriteback_6_bits_robIdx_value;
        input  io_exuWriteback_5_valid;
        input  io_exuWriteback_5_bits_data_0;
        input  io_exuWriteback_5_bits_robIdx_value;
        input  io_exuWriteback_5_bits_redirect_valid;
        input  io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken;
        input  io_exuWriteback_5_bits_fflags;
        input  io_exuWriteback_5_bits_wflags;
        input  io_exuWriteback_4_valid;
        input  io_exuWriteback_4_bits_data_0;
        input  io_exuWriteback_4_bits_robIdx_value;
        input  io_exuWriteback_3_valid;
        input  io_exuWriteback_3_bits_data_0;
        input  io_exuWriteback_3_bits_robIdx_value;
        input  io_exuWriteback_3_bits_redirect_valid;
        input  io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken;
        input  io_exuWriteback_2_valid;
        input  io_exuWriteback_2_bits_data_0;
        input  io_exuWriteback_2_bits_robIdx_value;
        input  io_exuWriteback_1_valid;
        input  io_exuWriteback_1_bits_data_0;
        input  io_exuWriteback_1_bits_robIdx_value;
        input  io_exuWriteback_1_bits_redirect_valid;
        input  io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken;
        input  io_exuWriteback_0_valid;
        input  io_exuWriteback_0_bits_data_0;
        input  io_exuWriteback_0_bits_robIdx_value;
        input  io_writebackNums_0_bits;
        input  io_writebackNums_1_bits;
        input  io_writebackNums_2_bits;
        input  io_writebackNums_3_bits;
        input  io_writebackNums_4_bits;
        input  io_writebackNums_5_bits;
        input  io_writebackNums_6_bits;
        input  io_writebackNums_7_bits;
        input  io_writebackNums_8_bits;
        input  io_writebackNums_9_bits;
        input  io_writebackNums_10_bits;
        input  io_writebackNums_11_bits;
        input  io_writebackNums_12_bits;
        input  io_writebackNums_13_bits;
        input  io_writebackNums_14_bits;
        input  io_writebackNums_15_bits;
        input  io_writebackNums_16_bits;
        input  io_writebackNums_17_bits;
        input  io_writebackNums_18_bits;
        input  io_writebackNums_19_bits;
        input  io_writebackNums_20_bits;
        input  io_writebackNums_21_bits;
        input  io_writebackNums_22_bits;
        input  io_writebackNums_23_bits;
        input  io_writebackNums_24_bits;
        input  io_writebackNeedFlush_0;
        input  io_writebackNeedFlush_1;
        input  io_writebackNeedFlush_2;
        input  io_writebackNeedFlush_6;
        input  io_writebackNeedFlush_7;
        input  io_writebackNeedFlush_8;
        input  io_writebackNeedFlush_9;
        input  io_writebackNeedFlush_10;
        input  io_writebackNeedFlush_11;
        input  io_writebackNeedFlush_12;

    endclocking:mon_cb

    modport drv_mp (clocking drv_cb);
    modport mon_mp (clocking mon_cb);

endinterface:WriteBack_in_agent_interface

`endif


//=========================================================
//File name    : WriteBack_in_agent_driver.sv
//Author       : nanyunhao
//Module name  : WriteBack_in_agent_driver
//Discribution : WriteBack_in_agent_driver : driver
//Date         : 2026-01-22
//=========================================================
`ifndef WRITEBACK_IN_AGENT_DRIVER__SV
`define WRITEBACK_IN_AGENT_DRIVER__SV

class WriteBack_in_agent_driver  extends tcnt_driver_base#(virtual WriteBack_in_agent_interface,WriteBack_in_agent_cfg,WriteBack_in_agent_xaction);

    `uvm_component_utils(WriteBack_in_agent_driver)

    extern function new(string name, uvm_component parent);
    extern virtual function void build_phase(uvm_phase phase);
    extern virtual task reset_phase(uvm_phase phase);
    extern task main_phase(uvm_phase phase);
    extern task send_pkt(WriteBack_in_agent_xaction tr);
    extern task drive_idle(tcnt_dec_base::drv_mode_e drv_mode);
endclass:WriteBack_in_agent_driver

function WriteBack_in_agent_driver::new(string name, uvm_component parent);
    super.new(name,parent);
endfunction:new

function void WriteBack_in_agent_driver::build_phase(uvm_phase phase);
    super.build_phase(phase);
endfunction:build_phase

task WriteBack_in_agent_driver::reset_phase(uvm_phase phase);

    super.reset_phase(phase);
    phase.raise_objection(this);

    repeat(2) begin
        @this.vif.drv_mp.drv_cb;
        this.drive_idle(this.cfg.drv_mode);
    end
    wait(vif.rst_n == 1'b1);
    repeat(20) begin
        @this.vif.drv_mp.drv_cb;
        this.drive_idle(this.cfg.drv_mode);
    end

    phase.drop_objection(this);
endtask:reset_phase

task WriteBack_in_agent_driver::main_phase(uvm_phase phase);
    super.main_phase(phase);
    //while(1) begin
    if(this.cfg.sqr_sw==tcnt_dec_base::ON && this.cfg.drv_sw==tcnt_dec_base::ON) begin
        while(1) begin
            seq_item_port.try_next_item(req);
            if(req!=null) begin
                repeat(req.pre_pkt_gap) begin
                    @this.vif.drv_mp.drv_cb;
                    this.drive_idle(this.cfg.drv_mode);
                end
                @this.vif.drv_mp.drv_cb;
                this.send_pkt(req);
                repeat(req.post_pkt_gap) begin
                    @this.vif.drv_mp.drv_cb;
                    this.drive_idle(this.cfg.drv_mode);
                end
                seq_item_port.item_done();
            end
            else begin
                @this.vif.drv_mp.drv_cb;
                this.drive_idle(this.cfg.drv_mode);
            end
        end
    end
    else if (this.cfg.drv_sw==tcnt_dec_base::ON) begin
        while(1) begin
            @this.vif.drv_mp.drv_cb;
            `uvm_fatal(get_type_name(), $sformatf("sqr_sw==OFF & drv_sw==ON, please give a driver send task!"))
            //send task
        end
    end
endtask:main_phase

task WriteBack_in_agent_driver::send_pkt(WriteBack_in_agent_xaction tr);
    vif.drv_mp.drv_cb.io_writeback_24_valid <= tr.io_writeback_24_valid; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_data_0 <= tr.io_writeback_24_bits_data_0; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_pdest <= tr.io_writeback_24_bits_pdest; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_robIdx_flag <= tr.io_writeback_24_bits_robIdx_flag; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_robIdx_value <= tr.io_writeback_24_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vecWen <= tr.io_writeback_24_bits_vecWen; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_v0Wen <= tr.io_writeback_24_bits_v0Wen; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vlWen <= tr.io_writeback_24_bits_vlWen; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_0 <= tr.io_writeback_24_bits_exceptionVec_0; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_1 <= tr.io_writeback_24_bits_exceptionVec_1; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_2 <= tr.io_writeback_24_bits_exceptionVec_2; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_3 <= tr.io_writeback_24_bits_exceptionVec_3; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_4 <= tr.io_writeback_24_bits_exceptionVec_4; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_5 <= tr.io_writeback_24_bits_exceptionVec_5; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_6 <= tr.io_writeback_24_bits_exceptionVec_6; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_7 <= tr.io_writeback_24_bits_exceptionVec_7; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_8 <= tr.io_writeback_24_bits_exceptionVec_8; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_9 <= tr.io_writeback_24_bits_exceptionVec_9; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_10 <= tr.io_writeback_24_bits_exceptionVec_10; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_11 <= tr.io_writeback_24_bits_exceptionVec_11; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_12 <= tr.io_writeback_24_bits_exceptionVec_12; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_13 <= tr.io_writeback_24_bits_exceptionVec_13; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_14 <= tr.io_writeback_24_bits_exceptionVec_14; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_15 <= tr.io_writeback_24_bits_exceptionVec_15; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_16 <= tr.io_writeback_24_bits_exceptionVec_16; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_17 <= tr.io_writeback_24_bits_exceptionVec_17; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_18 <= tr.io_writeback_24_bits_exceptionVec_18; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_19 <= tr.io_writeback_24_bits_exceptionVec_19; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_20 <= tr.io_writeback_24_bits_exceptionVec_20; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_21 <= tr.io_writeback_24_bits_exceptionVec_21; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_22 <= tr.io_writeback_24_bits_exceptionVec_22; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_23 <= tr.io_writeback_24_bits_exceptionVec_23; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_flushPipe <= tr.io_writeback_24_bits_flushPipe; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_replay <= tr.io_writeback_24_bits_replay; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_trigger <= tr.io_writeback_24_bits_trigger; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vill <= tr.io_writeback_24_bits_vls_vpu_vill; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vma <= tr.io_writeback_24_bits_vls_vpu_vma; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vta <= tr.io_writeback_24_bits_vls_vpu_vta; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vsew <= tr.io_writeback_24_bits_vls_vpu_vsew; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vlmul <= tr.io_writeback_24_bits_vls_vpu_vlmul; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVill <= tr.io_writeback_24_bits_vls_vpu_specVill; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVma <= tr.io_writeback_24_bits_vls_vpu_specVma; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVta <= tr.io_writeback_24_bits_vls_vpu_specVta; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVsew <= tr.io_writeback_24_bits_vls_vpu_specVsew; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVlmul <= tr.io_writeback_24_bits_vls_vpu_specVlmul; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vm <= tr.io_writeback_24_bits_vls_vpu_vm; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vstart <= tr.io_writeback_24_bits_vls_vpu_vstart; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_frm <= tr.io_writeback_24_bits_vls_vpu_frm; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst <= tr.io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFP32Instr <= tr.io_writeback_24_bits_vls_vpu_fpu_isFP32Instr; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFP64Instr <= tr.io_writeback_24_bits_vls_vpu_fpu_isFP64Instr; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isReduction <= tr.io_writeback_24_bits_vls_vpu_fpu_isReduction; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2 <= tr.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4 <= tr.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8 <= tr.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vxrm <= tr.io_writeback_24_bits_vls_vpu_vxrm; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vuopIdx <= tr.io_writeback_24_bits_vls_vpu_vuopIdx; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_lastUop <= tr.io_writeback_24_bits_vls_vpu_lastUop; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vmask <= tr.io_writeback_24_bits_vls_vpu_vmask; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vl <= tr.io_writeback_24_bits_vls_vpu_vl; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_nf <= tr.io_writeback_24_bits_vls_vpu_nf; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_veew <= tr.io_writeback_24_bits_vls_vpu_veew; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isReverse <= tr.io_writeback_24_bits_vls_vpu_isReverse; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isExt <= tr.io_writeback_24_bits_vls_vpu_isExt; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isNarrow <= tr.io_writeback_24_bits_vls_vpu_isNarrow; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isDstMask <= tr.io_writeback_24_bits_vls_vpu_isDstMask; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isOpMask <= tr.io_writeback_24_bits_vls_vpu_isOpMask; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isMove <= tr.io_writeback_24_bits_vls_vpu_isMove; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isDependOldVd <= tr.io_writeback_24_bits_vls_vpu_isDependOldVd; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isWritePartVd <= tr.io_writeback_24_bits_vls_vpu_isWritePartVd; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isVleff <= tr.io_writeback_24_bits_vls_vpu_isVleff; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_oldVdPsrc <= tr.io_writeback_24_bits_vls_oldVdPsrc; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vdIdx <= tr.io_writeback_24_bits_vls_vdIdx; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vdIdxInField <= tr.io_writeback_24_bits_vls_vdIdxInField; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isIndexed <= tr.io_writeback_24_bits_vls_isIndexed; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isMasked <= tr.io_writeback_24_bits_vls_isMasked; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isStrided <= tr.io_writeback_24_bits_vls_isStrided; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isWhole <= tr.io_writeback_24_bits_vls_isWhole; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isVecLoad <= tr.io_writeback_24_bits_vls_isVecLoad; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isVlm <= tr.io_writeback_24_bits_vls_isVlm; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_debug_isMMIO <= tr.io_writeback_24_bits_debug_isMMIO; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_debug_isNCIO <= tr.io_writeback_24_bits_debug_isNCIO; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_debug_isPerfCnt <= tr.io_writeback_24_bits_debug_isPerfCnt; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_debug_paddr <= tr.io_writeback_24_bits_debug_paddr; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_debug_vaddr <= tr.io_writeback_24_bits_debug_vaddr; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_eliminatedMove <= tr.io_writeback_24_bits_debugInfo_eliminatedMove; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_renameTime <= tr.io_writeback_24_bits_debugInfo_renameTime; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_dispatchTime <= tr.io_writeback_24_bits_debugInfo_dispatchTime; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_enqRsTime <= tr.io_writeback_24_bits_debugInfo_enqRsTime; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_selectTime <= tr.io_writeback_24_bits_debugInfo_selectTime; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_issueTime <= tr.io_writeback_24_bits_debugInfo_issueTime; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_writebackTime <= tr.io_writeback_24_bits_debugInfo_writebackTime; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_runahead_checkpoint_id <= tr.io_writeback_24_bits_debugInfo_runahead_checkpoint_id; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_tlbFirstReqTime <= tr.io_writeback_24_bits_debugInfo_tlbFirstReqTime; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_tlbRespTime <= tr.io_writeback_24_bits_debugInfo_tlbRespTime; 
    vif.drv_mp.drv_cb.io_writeback_24_bits_debug_seqNum <= tr.io_writeback_24_bits_debug_seqNum; 
    vif.drv_mp.drv_cb.io_writeback_23_valid <= tr.io_writeback_23_valid; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_data_0 <= tr.io_writeback_23_bits_data_0; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_pdest <= tr.io_writeback_23_bits_pdest; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_robIdx_flag <= tr.io_writeback_23_bits_robIdx_flag; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_robIdx_value <= tr.io_writeback_23_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vecWen <= tr.io_writeback_23_bits_vecWen; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_v0Wen <= tr.io_writeback_23_bits_v0Wen; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vlWen <= tr.io_writeback_23_bits_vlWen; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_0 <= tr.io_writeback_23_bits_exceptionVec_0; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_1 <= tr.io_writeback_23_bits_exceptionVec_1; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_2 <= tr.io_writeback_23_bits_exceptionVec_2; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_3 <= tr.io_writeback_23_bits_exceptionVec_3; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_4 <= tr.io_writeback_23_bits_exceptionVec_4; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_5 <= tr.io_writeback_23_bits_exceptionVec_5; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_6 <= tr.io_writeback_23_bits_exceptionVec_6; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_7 <= tr.io_writeback_23_bits_exceptionVec_7; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_8 <= tr.io_writeback_23_bits_exceptionVec_8; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_9 <= tr.io_writeback_23_bits_exceptionVec_9; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_10 <= tr.io_writeback_23_bits_exceptionVec_10; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_11 <= tr.io_writeback_23_bits_exceptionVec_11; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_12 <= tr.io_writeback_23_bits_exceptionVec_12; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_13 <= tr.io_writeback_23_bits_exceptionVec_13; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_14 <= tr.io_writeback_23_bits_exceptionVec_14; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_15 <= tr.io_writeback_23_bits_exceptionVec_15; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_16 <= tr.io_writeback_23_bits_exceptionVec_16; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_17 <= tr.io_writeback_23_bits_exceptionVec_17; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_18 <= tr.io_writeback_23_bits_exceptionVec_18; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_19 <= tr.io_writeback_23_bits_exceptionVec_19; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_20 <= tr.io_writeback_23_bits_exceptionVec_20; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_21 <= tr.io_writeback_23_bits_exceptionVec_21; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_22 <= tr.io_writeback_23_bits_exceptionVec_22; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_23 <= tr.io_writeback_23_bits_exceptionVec_23; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_flushPipe <= tr.io_writeback_23_bits_flushPipe; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_replay <= tr.io_writeback_23_bits_replay; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_trigger <= tr.io_writeback_23_bits_trigger; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vill <= tr.io_writeback_23_bits_vls_vpu_vill; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vma <= tr.io_writeback_23_bits_vls_vpu_vma; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vta <= tr.io_writeback_23_bits_vls_vpu_vta; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vsew <= tr.io_writeback_23_bits_vls_vpu_vsew; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vlmul <= tr.io_writeback_23_bits_vls_vpu_vlmul; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVill <= tr.io_writeback_23_bits_vls_vpu_specVill; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVma <= tr.io_writeback_23_bits_vls_vpu_specVma; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVta <= tr.io_writeback_23_bits_vls_vpu_specVta; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVsew <= tr.io_writeback_23_bits_vls_vpu_specVsew; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVlmul <= tr.io_writeback_23_bits_vls_vpu_specVlmul; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vm <= tr.io_writeback_23_bits_vls_vpu_vm; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vstart <= tr.io_writeback_23_bits_vls_vpu_vstart; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_frm <= tr.io_writeback_23_bits_vls_vpu_frm; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst <= tr.io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFP32Instr <= tr.io_writeback_23_bits_vls_vpu_fpu_isFP32Instr; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFP64Instr <= tr.io_writeback_23_bits_vls_vpu_fpu_isFP64Instr; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isReduction <= tr.io_writeback_23_bits_vls_vpu_fpu_isReduction; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2 <= tr.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4 <= tr.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8 <= tr.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vxrm <= tr.io_writeback_23_bits_vls_vpu_vxrm; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vuopIdx <= tr.io_writeback_23_bits_vls_vpu_vuopIdx; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_lastUop <= tr.io_writeback_23_bits_vls_vpu_lastUop; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vmask <= tr.io_writeback_23_bits_vls_vpu_vmask; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vl <= tr.io_writeback_23_bits_vls_vpu_vl; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_nf <= tr.io_writeback_23_bits_vls_vpu_nf; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_veew <= tr.io_writeback_23_bits_vls_vpu_veew; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isReverse <= tr.io_writeback_23_bits_vls_vpu_isReverse; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isExt <= tr.io_writeback_23_bits_vls_vpu_isExt; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isNarrow <= tr.io_writeback_23_bits_vls_vpu_isNarrow; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isDstMask <= tr.io_writeback_23_bits_vls_vpu_isDstMask; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isOpMask <= tr.io_writeback_23_bits_vls_vpu_isOpMask; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isMove <= tr.io_writeback_23_bits_vls_vpu_isMove; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isDependOldVd <= tr.io_writeback_23_bits_vls_vpu_isDependOldVd; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isWritePartVd <= tr.io_writeback_23_bits_vls_vpu_isWritePartVd; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isVleff <= tr.io_writeback_23_bits_vls_vpu_isVleff; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_oldVdPsrc <= tr.io_writeback_23_bits_vls_oldVdPsrc; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vdIdx <= tr.io_writeback_23_bits_vls_vdIdx; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vdIdxInField <= tr.io_writeback_23_bits_vls_vdIdxInField; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isIndexed <= tr.io_writeback_23_bits_vls_isIndexed; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isMasked <= tr.io_writeback_23_bits_vls_isMasked; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isStrided <= tr.io_writeback_23_bits_vls_isStrided; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isWhole <= tr.io_writeback_23_bits_vls_isWhole; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isVecLoad <= tr.io_writeback_23_bits_vls_isVecLoad; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isVlm <= tr.io_writeback_23_bits_vls_isVlm; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_debug_isMMIO <= tr.io_writeback_23_bits_debug_isMMIO; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_debug_isNCIO <= tr.io_writeback_23_bits_debug_isNCIO; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_debug_isPerfCnt <= tr.io_writeback_23_bits_debug_isPerfCnt; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_debug_paddr <= tr.io_writeback_23_bits_debug_paddr; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_debug_vaddr <= tr.io_writeback_23_bits_debug_vaddr; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_eliminatedMove <= tr.io_writeback_23_bits_debugInfo_eliminatedMove; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_renameTime <= tr.io_writeback_23_bits_debugInfo_renameTime; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_dispatchTime <= tr.io_writeback_23_bits_debugInfo_dispatchTime; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_enqRsTime <= tr.io_writeback_23_bits_debugInfo_enqRsTime; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_selectTime <= tr.io_writeback_23_bits_debugInfo_selectTime; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_issueTime <= tr.io_writeback_23_bits_debugInfo_issueTime; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_writebackTime <= tr.io_writeback_23_bits_debugInfo_writebackTime; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_runahead_checkpoint_id <= tr.io_writeback_23_bits_debugInfo_runahead_checkpoint_id; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_tlbFirstReqTime <= tr.io_writeback_23_bits_debugInfo_tlbFirstReqTime; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_tlbRespTime <= tr.io_writeback_23_bits_debugInfo_tlbRespTime; 
    vif.drv_mp.drv_cb.io_writeback_23_bits_debug_seqNum <= tr.io_writeback_23_bits_debug_seqNum; 
    vif.drv_mp.drv_cb.io_writeback_22_valid <= tr.io_writeback_22_valid; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_data_0 <= tr.io_writeback_22_bits_data_0; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_pdest <= tr.io_writeback_22_bits_pdest; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_robIdx_flag <= tr.io_writeback_22_bits_robIdx_flag; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_robIdx_value <= tr.io_writeback_22_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_intWen <= tr.io_writeback_22_bits_intWen; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_fpWen <= tr.io_writeback_22_bits_fpWen; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_0 <= tr.io_writeback_22_bits_exceptionVec_0; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_1 <= tr.io_writeback_22_bits_exceptionVec_1; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_2 <= tr.io_writeback_22_bits_exceptionVec_2; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_3 <= tr.io_writeback_22_bits_exceptionVec_3; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_4 <= tr.io_writeback_22_bits_exceptionVec_4; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_5 <= tr.io_writeback_22_bits_exceptionVec_5; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_6 <= tr.io_writeback_22_bits_exceptionVec_6; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_7 <= tr.io_writeback_22_bits_exceptionVec_7; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_8 <= tr.io_writeback_22_bits_exceptionVec_8; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_9 <= tr.io_writeback_22_bits_exceptionVec_9; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_10 <= tr.io_writeback_22_bits_exceptionVec_10; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_11 <= tr.io_writeback_22_bits_exceptionVec_11; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_12 <= tr.io_writeback_22_bits_exceptionVec_12; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_13 <= tr.io_writeback_22_bits_exceptionVec_13; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_14 <= tr.io_writeback_22_bits_exceptionVec_14; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_15 <= tr.io_writeback_22_bits_exceptionVec_15; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_16 <= tr.io_writeback_22_bits_exceptionVec_16; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_17 <= tr.io_writeback_22_bits_exceptionVec_17; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_18 <= tr.io_writeback_22_bits_exceptionVec_18; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_19 <= tr.io_writeback_22_bits_exceptionVec_19; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_20 <= tr.io_writeback_22_bits_exceptionVec_20; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_21 <= tr.io_writeback_22_bits_exceptionVec_21; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_22 <= tr.io_writeback_22_bits_exceptionVec_22; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_23 <= tr.io_writeback_22_bits_exceptionVec_23; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_flushPipe <= tr.io_writeback_22_bits_flushPipe; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_replay <= tr.io_writeback_22_bits_replay; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_lqIdx_flag <= tr.io_writeback_22_bits_lqIdx_flag; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_lqIdx_value <= tr.io_writeback_22_bits_lqIdx_value; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_trigger <= tr.io_writeback_22_bits_trigger; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_valid <= tr.io_writeback_22_bits_predecodeInfo_valid; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_isRVC <= tr.io_writeback_22_bits_predecodeInfo_isRVC; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_brType <= tr.io_writeback_22_bits_predecodeInfo_brType; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_isCall <= tr.io_writeback_22_bits_predecodeInfo_isCall; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_isRet <= tr.io_writeback_22_bits_predecodeInfo_isRet; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_debug_isMMIO <= tr.io_writeback_22_bits_debug_isMMIO; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_debug_isNCIO <= tr.io_writeback_22_bits_debug_isNCIO; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_debug_isPerfCnt <= tr.io_writeback_22_bits_debug_isPerfCnt; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_debug_paddr <= tr.io_writeback_22_bits_debug_paddr; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_debug_vaddr <= tr.io_writeback_22_bits_debug_vaddr; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_eliminatedMove <= tr.io_writeback_22_bits_debugInfo_eliminatedMove; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_renameTime <= tr.io_writeback_22_bits_debugInfo_renameTime; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_dispatchTime <= tr.io_writeback_22_bits_debugInfo_dispatchTime; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_enqRsTime <= tr.io_writeback_22_bits_debugInfo_enqRsTime; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_selectTime <= tr.io_writeback_22_bits_debugInfo_selectTime; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_issueTime <= tr.io_writeback_22_bits_debugInfo_issueTime; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_writebackTime <= tr.io_writeback_22_bits_debugInfo_writebackTime; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_runahead_checkpoint_id <= tr.io_writeback_22_bits_debugInfo_runahead_checkpoint_id; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_tlbFirstReqTime <= tr.io_writeback_22_bits_debugInfo_tlbFirstReqTime; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_tlbRespTime <= tr.io_writeback_22_bits_debugInfo_tlbRespTime; 
    vif.drv_mp.drv_cb.io_writeback_22_bits_debug_seqNum <= tr.io_writeback_22_bits_debug_seqNum; 
    vif.drv_mp.drv_cb.io_writeback_21_valid <= tr.io_writeback_21_valid; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_data_0 <= tr.io_writeback_21_bits_data_0; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_pdest <= tr.io_writeback_21_bits_pdest; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_robIdx_flag <= tr.io_writeback_21_bits_robIdx_flag; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_robIdx_value <= tr.io_writeback_21_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_intWen <= tr.io_writeback_21_bits_intWen; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_fpWen <= tr.io_writeback_21_bits_fpWen; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_0 <= tr.io_writeback_21_bits_exceptionVec_0; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_1 <= tr.io_writeback_21_bits_exceptionVec_1; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_2 <= tr.io_writeback_21_bits_exceptionVec_2; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_3 <= tr.io_writeback_21_bits_exceptionVec_3; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_4 <= tr.io_writeback_21_bits_exceptionVec_4; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_5 <= tr.io_writeback_21_bits_exceptionVec_5; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_6 <= tr.io_writeback_21_bits_exceptionVec_6; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_7 <= tr.io_writeback_21_bits_exceptionVec_7; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_8 <= tr.io_writeback_21_bits_exceptionVec_8; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_9 <= tr.io_writeback_21_bits_exceptionVec_9; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_10 <= tr.io_writeback_21_bits_exceptionVec_10; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_11 <= tr.io_writeback_21_bits_exceptionVec_11; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_12 <= tr.io_writeback_21_bits_exceptionVec_12; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_13 <= tr.io_writeback_21_bits_exceptionVec_13; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_14 <= tr.io_writeback_21_bits_exceptionVec_14; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_15 <= tr.io_writeback_21_bits_exceptionVec_15; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_16 <= tr.io_writeback_21_bits_exceptionVec_16; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_17 <= tr.io_writeback_21_bits_exceptionVec_17; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_18 <= tr.io_writeback_21_bits_exceptionVec_18; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_19 <= tr.io_writeback_21_bits_exceptionVec_19; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_20 <= tr.io_writeback_21_bits_exceptionVec_20; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_21 <= tr.io_writeback_21_bits_exceptionVec_21; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_22 <= tr.io_writeback_21_bits_exceptionVec_22; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_23 <= tr.io_writeback_21_bits_exceptionVec_23; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_flushPipe <= tr.io_writeback_21_bits_flushPipe; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_replay <= tr.io_writeback_21_bits_replay; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_lqIdx_flag <= tr.io_writeback_21_bits_lqIdx_flag; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_lqIdx_value <= tr.io_writeback_21_bits_lqIdx_value; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_trigger <= tr.io_writeback_21_bits_trigger; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_valid <= tr.io_writeback_21_bits_predecodeInfo_valid; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_isRVC <= tr.io_writeback_21_bits_predecodeInfo_isRVC; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_brType <= tr.io_writeback_21_bits_predecodeInfo_brType; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_isCall <= tr.io_writeback_21_bits_predecodeInfo_isCall; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_isRet <= tr.io_writeback_21_bits_predecodeInfo_isRet; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_debug_isMMIO <= tr.io_writeback_21_bits_debug_isMMIO; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_debug_isNCIO <= tr.io_writeback_21_bits_debug_isNCIO; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_debug_isPerfCnt <= tr.io_writeback_21_bits_debug_isPerfCnt; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_debug_paddr <= tr.io_writeback_21_bits_debug_paddr; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_debug_vaddr <= tr.io_writeback_21_bits_debug_vaddr; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_eliminatedMove <= tr.io_writeback_21_bits_debugInfo_eliminatedMove; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_renameTime <= tr.io_writeback_21_bits_debugInfo_renameTime; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_dispatchTime <= tr.io_writeback_21_bits_debugInfo_dispatchTime; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_enqRsTime <= tr.io_writeback_21_bits_debugInfo_enqRsTime; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_selectTime <= tr.io_writeback_21_bits_debugInfo_selectTime; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_issueTime <= tr.io_writeback_21_bits_debugInfo_issueTime; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_writebackTime <= tr.io_writeback_21_bits_debugInfo_writebackTime; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_runahead_checkpoint_id <= tr.io_writeback_21_bits_debugInfo_runahead_checkpoint_id; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_tlbFirstReqTime <= tr.io_writeback_21_bits_debugInfo_tlbFirstReqTime; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_tlbRespTime <= tr.io_writeback_21_bits_debugInfo_tlbRespTime; 
    vif.drv_mp.drv_cb.io_writeback_21_bits_debug_seqNum <= tr.io_writeback_21_bits_debug_seqNum; 
    vif.drv_mp.drv_cb.io_writeback_20_valid <= tr.io_writeback_20_valid; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_data_0 <= tr.io_writeback_20_bits_data_0; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_pdest <= tr.io_writeback_20_bits_pdest; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_robIdx_flag <= tr.io_writeback_20_bits_robIdx_flag; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_robIdx_value <= tr.io_writeback_20_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_intWen <= tr.io_writeback_20_bits_intWen; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_fpWen <= tr.io_writeback_20_bits_fpWen; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_0 <= tr.io_writeback_20_bits_exceptionVec_0; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_1 <= tr.io_writeback_20_bits_exceptionVec_1; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_2 <= tr.io_writeback_20_bits_exceptionVec_2; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_3 <= tr.io_writeback_20_bits_exceptionVec_3; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_4 <= tr.io_writeback_20_bits_exceptionVec_4; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_5 <= tr.io_writeback_20_bits_exceptionVec_5; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_6 <= tr.io_writeback_20_bits_exceptionVec_6; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_7 <= tr.io_writeback_20_bits_exceptionVec_7; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_8 <= tr.io_writeback_20_bits_exceptionVec_8; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_9 <= tr.io_writeback_20_bits_exceptionVec_9; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_10 <= tr.io_writeback_20_bits_exceptionVec_10; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_11 <= tr.io_writeback_20_bits_exceptionVec_11; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_12 <= tr.io_writeback_20_bits_exceptionVec_12; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_13 <= tr.io_writeback_20_bits_exceptionVec_13; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_14 <= tr.io_writeback_20_bits_exceptionVec_14; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_15 <= tr.io_writeback_20_bits_exceptionVec_15; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_16 <= tr.io_writeback_20_bits_exceptionVec_16; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_17 <= tr.io_writeback_20_bits_exceptionVec_17; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_18 <= tr.io_writeback_20_bits_exceptionVec_18; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_19 <= tr.io_writeback_20_bits_exceptionVec_19; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_20 <= tr.io_writeback_20_bits_exceptionVec_20; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_21 <= tr.io_writeback_20_bits_exceptionVec_21; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_22 <= tr.io_writeback_20_bits_exceptionVec_22; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_23 <= tr.io_writeback_20_bits_exceptionVec_23; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_flushPipe <= tr.io_writeback_20_bits_flushPipe; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_replay <= tr.io_writeback_20_bits_replay; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_lqIdx_flag <= tr.io_writeback_20_bits_lqIdx_flag; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_lqIdx_value <= tr.io_writeback_20_bits_lqIdx_value; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_trigger <= tr.io_writeback_20_bits_trigger; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_valid <= tr.io_writeback_20_bits_predecodeInfo_valid; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_isRVC <= tr.io_writeback_20_bits_predecodeInfo_isRVC; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_brType <= tr.io_writeback_20_bits_predecodeInfo_brType; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_isCall <= tr.io_writeback_20_bits_predecodeInfo_isCall; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_isRet <= tr.io_writeback_20_bits_predecodeInfo_isRet; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_debug_isMMIO <= tr.io_writeback_20_bits_debug_isMMIO; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_debug_isNCIO <= tr.io_writeback_20_bits_debug_isNCIO; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_debug_isPerfCnt <= tr.io_writeback_20_bits_debug_isPerfCnt; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_debug_paddr <= tr.io_writeback_20_bits_debug_paddr; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_debug_vaddr <= tr.io_writeback_20_bits_debug_vaddr; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_eliminatedMove <= tr.io_writeback_20_bits_debugInfo_eliminatedMove; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_renameTime <= tr.io_writeback_20_bits_debugInfo_renameTime; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_dispatchTime <= tr.io_writeback_20_bits_debugInfo_dispatchTime; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_enqRsTime <= tr.io_writeback_20_bits_debugInfo_enqRsTime; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_selectTime <= tr.io_writeback_20_bits_debugInfo_selectTime; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_issueTime <= tr.io_writeback_20_bits_debugInfo_issueTime; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_writebackTime <= tr.io_writeback_20_bits_debugInfo_writebackTime; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_runahead_checkpoint_id <= tr.io_writeback_20_bits_debugInfo_runahead_checkpoint_id; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_tlbFirstReqTime <= tr.io_writeback_20_bits_debugInfo_tlbFirstReqTime; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_tlbRespTime <= tr.io_writeback_20_bits_debugInfo_tlbRespTime; 
    vif.drv_mp.drv_cb.io_writeback_20_bits_debug_seqNum <= tr.io_writeback_20_bits_debug_seqNum; 
    vif.drv_mp.drv_cb.io_writeback_19_valid <= tr.io_writeback_19_valid; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_data_0 <= tr.io_writeback_19_bits_data_0; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_pdest <= tr.io_writeback_19_bits_pdest; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_robIdx_flag <= tr.io_writeback_19_bits_robIdx_flag; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_robIdx_value <= tr.io_writeback_19_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_intWen <= tr.io_writeback_19_bits_intWen; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_0 <= tr.io_writeback_19_bits_exceptionVec_0; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_1 <= tr.io_writeback_19_bits_exceptionVec_1; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_2 <= tr.io_writeback_19_bits_exceptionVec_2; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_3 <= tr.io_writeback_19_bits_exceptionVec_3; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_4 <= tr.io_writeback_19_bits_exceptionVec_4; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_5 <= tr.io_writeback_19_bits_exceptionVec_5; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_6 <= tr.io_writeback_19_bits_exceptionVec_6; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_7 <= tr.io_writeback_19_bits_exceptionVec_7; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_8 <= tr.io_writeback_19_bits_exceptionVec_8; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_9 <= tr.io_writeback_19_bits_exceptionVec_9; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_10 <= tr.io_writeback_19_bits_exceptionVec_10; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_11 <= tr.io_writeback_19_bits_exceptionVec_11; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_12 <= tr.io_writeback_19_bits_exceptionVec_12; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_13 <= tr.io_writeback_19_bits_exceptionVec_13; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_14 <= tr.io_writeback_19_bits_exceptionVec_14; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_15 <= tr.io_writeback_19_bits_exceptionVec_15; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_16 <= tr.io_writeback_19_bits_exceptionVec_16; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_17 <= tr.io_writeback_19_bits_exceptionVec_17; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_18 <= tr.io_writeback_19_bits_exceptionVec_18; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_19 <= tr.io_writeback_19_bits_exceptionVec_19; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_20 <= tr.io_writeback_19_bits_exceptionVec_20; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_21 <= tr.io_writeback_19_bits_exceptionVec_21; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_22 <= tr.io_writeback_19_bits_exceptionVec_22; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_23 <= tr.io_writeback_19_bits_exceptionVec_23; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_flushPipe <= tr.io_writeback_19_bits_flushPipe; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_sqIdx_flag <= tr.io_writeback_19_bits_sqIdx_flag; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_sqIdx_value <= tr.io_writeback_19_bits_sqIdx_value; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_trigger <= tr.io_writeback_19_bits_trigger; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_debug_isMMIO <= tr.io_writeback_19_bits_debug_isMMIO; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_debug_isNCIO <= tr.io_writeback_19_bits_debug_isNCIO; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_debug_isPerfCnt <= tr.io_writeback_19_bits_debug_isPerfCnt; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_debug_paddr <= tr.io_writeback_19_bits_debug_paddr; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_debug_vaddr <= tr.io_writeback_19_bits_debug_vaddr; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_eliminatedMove <= tr.io_writeback_19_bits_debugInfo_eliminatedMove; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_renameTime <= tr.io_writeback_19_bits_debugInfo_renameTime; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_dispatchTime <= tr.io_writeback_19_bits_debugInfo_dispatchTime; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_enqRsTime <= tr.io_writeback_19_bits_debugInfo_enqRsTime; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_selectTime <= tr.io_writeback_19_bits_debugInfo_selectTime; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_issueTime <= tr.io_writeback_19_bits_debugInfo_issueTime; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_writebackTime <= tr.io_writeback_19_bits_debugInfo_writebackTime; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_runahead_checkpoint_id <= tr.io_writeback_19_bits_debugInfo_runahead_checkpoint_id; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_tlbFirstReqTime <= tr.io_writeback_19_bits_debugInfo_tlbFirstReqTime; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_tlbRespTime <= tr.io_writeback_19_bits_debugInfo_tlbRespTime; 
    vif.drv_mp.drv_cb.io_writeback_19_bits_debug_seqNum <= tr.io_writeback_19_bits_debug_seqNum; 
    vif.drv_mp.drv_cb.io_writeback_18_valid <= tr.io_writeback_18_valid; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_data_0 <= tr.io_writeback_18_bits_data_0; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_pdest <= tr.io_writeback_18_bits_pdest; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_robIdx_flag <= tr.io_writeback_18_bits_robIdx_flag; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_robIdx_value <= tr.io_writeback_18_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_intWen <= tr.io_writeback_18_bits_intWen; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_0 <= tr.io_writeback_18_bits_exceptionVec_0; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_1 <= tr.io_writeback_18_bits_exceptionVec_1; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_2 <= tr.io_writeback_18_bits_exceptionVec_2; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_3 <= tr.io_writeback_18_bits_exceptionVec_3; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_4 <= tr.io_writeback_18_bits_exceptionVec_4; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_5 <= tr.io_writeback_18_bits_exceptionVec_5; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_6 <= tr.io_writeback_18_bits_exceptionVec_6; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_7 <= tr.io_writeback_18_bits_exceptionVec_7; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_8 <= tr.io_writeback_18_bits_exceptionVec_8; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_9 <= tr.io_writeback_18_bits_exceptionVec_9; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_10 <= tr.io_writeback_18_bits_exceptionVec_10; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_11 <= tr.io_writeback_18_bits_exceptionVec_11; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_12 <= tr.io_writeback_18_bits_exceptionVec_12; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_13 <= tr.io_writeback_18_bits_exceptionVec_13; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_14 <= tr.io_writeback_18_bits_exceptionVec_14; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_15 <= tr.io_writeback_18_bits_exceptionVec_15; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_16 <= tr.io_writeback_18_bits_exceptionVec_16; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_17 <= tr.io_writeback_18_bits_exceptionVec_17; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_18 <= tr.io_writeback_18_bits_exceptionVec_18; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_19 <= tr.io_writeback_18_bits_exceptionVec_19; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_20 <= tr.io_writeback_18_bits_exceptionVec_20; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_21 <= tr.io_writeback_18_bits_exceptionVec_21; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_22 <= tr.io_writeback_18_bits_exceptionVec_22; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_23 <= tr.io_writeback_18_bits_exceptionVec_23; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_flushPipe <= tr.io_writeback_18_bits_flushPipe; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_sqIdx_flag <= tr.io_writeback_18_bits_sqIdx_flag; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_sqIdx_value <= tr.io_writeback_18_bits_sqIdx_value; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_trigger <= tr.io_writeback_18_bits_trigger; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_debug_isMMIO <= tr.io_writeback_18_bits_debug_isMMIO; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_debug_isNCIO <= tr.io_writeback_18_bits_debug_isNCIO; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_debug_isPerfCnt <= tr.io_writeback_18_bits_debug_isPerfCnt; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_debug_paddr <= tr.io_writeback_18_bits_debug_paddr; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_debug_vaddr <= tr.io_writeback_18_bits_debug_vaddr; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_eliminatedMove <= tr.io_writeback_18_bits_debugInfo_eliminatedMove; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_renameTime <= tr.io_writeback_18_bits_debugInfo_renameTime; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_dispatchTime <= tr.io_writeback_18_bits_debugInfo_dispatchTime; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_enqRsTime <= tr.io_writeback_18_bits_debugInfo_enqRsTime; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_selectTime <= tr.io_writeback_18_bits_debugInfo_selectTime; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_issueTime <= tr.io_writeback_18_bits_debugInfo_issueTime; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_writebackTime <= tr.io_writeback_18_bits_debugInfo_writebackTime; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_runahead_checkpoint_id <= tr.io_writeback_18_bits_debugInfo_runahead_checkpoint_id; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_tlbFirstReqTime <= tr.io_writeback_18_bits_debugInfo_tlbFirstReqTime; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_tlbRespTime <= tr.io_writeback_18_bits_debugInfo_tlbRespTime; 
    vif.drv_mp.drv_cb.io_writeback_18_bits_debug_seqNum <= tr.io_writeback_18_bits_debug_seqNum; 
    vif.drv_mp.drv_cb.io_writeback_17_valid <= tr.io_writeback_17_valid; 
    vif.drv_mp.drv_cb.io_writeback_17_bits_data_0 <= tr.io_writeback_17_bits_data_0; 
    vif.drv_mp.drv_cb.io_writeback_17_bits_data_1 <= tr.io_writeback_17_bits_data_1; 
    vif.drv_mp.drv_cb.io_writeback_17_bits_data_2 <= tr.io_writeback_17_bits_data_2; 
    vif.drv_mp.drv_cb.io_writeback_17_bits_pdest <= tr.io_writeback_17_bits_pdest; 
    vif.drv_mp.drv_cb.io_writeback_17_bits_robIdx_flag <= tr.io_writeback_17_bits_robIdx_flag; 
    vif.drv_mp.drv_cb.io_writeback_17_bits_robIdx_value <= tr.io_writeback_17_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_writeback_17_bits_vecWen <= tr.io_writeback_17_bits_vecWen; 
    vif.drv_mp.drv_cb.io_writeback_17_bits_v0Wen <= tr.io_writeback_17_bits_v0Wen; 
    vif.drv_mp.drv_cb.io_writeback_17_bits_fflags <= tr.io_writeback_17_bits_fflags; 
    vif.drv_mp.drv_cb.io_writeback_17_bits_wflags <= tr.io_writeback_17_bits_wflags; 
    vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_eliminatedMove <= tr.io_writeback_17_bits_debugInfo_eliminatedMove; 
    vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_renameTime <= tr.io_writeback_17_bits_debugInfo_renameTime; 
    vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_dispatchTime <= tr.io_writeback_17_bits_debugInfo_dispatchTime; 
    vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_enqRsTime <= tr.io_writeback_17_bits_debugInfo_enqRsTime; 
    vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_selectTime <= tr.io_writeback_17_bits_debugInfo_selectTime; 
    vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_issueTime <= tr.io_writeback_17_bits_debugInfo_issueTime; 
    vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_writebackTime <= tr.io_writeback_17_bits_debugInfo_writebackTime; 
    vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_runahead_checkpoint_id <= tr.io_writeback_17_bits_debugInfo_runahead_checkpoint_id; 
    vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_tlbFirstReqTime <= tr.io_writeback_17_bits_debugInfo_tlbFirstReqTime; 
    vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_tlbRespTime <= tr.io_writeback_17_bits_debugInfo_tlbRespTime; 
    vif.drv_mp.drv_cb.io_writeback_17_bits_debug_seqNum <= tr.io_writeback_17_bits_debug_seqNum; 
    vif.drv_mp.drv_cb.io_writeback_16_valid <= tr.io_writeback_16_valid; 
    vif.drv_mp.drv_cb.io_writeback_16_bits_data_0 <= tr.io_writeback_16_bits_data_0; 
    vif.drv_mp.drv_cb.io_writeback_16_bits_data_1 <= tr.io_writeback_16_bits_data_1; 
    vif.drv_mp.drv_cb.io_writeback_16_bits_data_2 <= tr.io_writeback_16_bits_data_2; 
    vif.drv_mp.drv_cb.io_writeback_16_bits_data_3 <= tr.io_writeback_16_bits_data_3; 
    vif.drv_mp.drv_cb.io_writeback_16_bits_pdest <= tr.io_writeback_16_bits_pdest; 
    vif.drv_mp.drv_cb.io_writeback_16_bits_robIdx_flag <= tr.io_writeback_16_bits_robIdx_flag; 
    vif.drv_mp.drv_cb.io_writeback_16_bits_robIdx_value <= tr.io_writeback_16_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_writeback_16_bits_fpWen <= tr.io_writeback_16_bits_fpWen; 
    vif.drv_mp.drv_cb.io_writeback_16_bits_vecWen <= tr.io_writeback_16_bits_vecWen; 
    vif.drv_mp.drv_cb.io_writeback_16_bits_v0Wen <= tr.io_writeback_16_bits_v0Wen; 
    vif.drv_mp.drv_cb.io_writeback_16_bits_fflags <= tr.io_writeback_16_bits_fflags; 
    vif.drv_mp.drv_cb.io_writeback_16_bits_wflags <= tr.io_writeback_16_bits_wflags; 
    vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_eliminatedMove <= tr.io_writeback_16_bits_debugInfo_eliminatedMove; 
    vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_renameTime <= tr.io_writeback_16_bits_debugInfo_renameTime; 
    vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_dispatchTime <= tr.io_writeback_16_bits_debugInfo_dispatchTime; 
    vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_enqRsTime <= tr.io_writeback_16_bits_debugInfo_enqRsTime; 
    vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_selectTime <= tr.io_writeback_16_bits_debugInfo_selectTime; 
    vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_issueTime <= tr.io_writeback_16_bits_debugInfo_issueTime; 
    vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_writebackTime <= tr.io_writeback_16_bits_debugInfo_writebackTime; 
    vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_runahead_checkpoint_id <= tr.io_writeback_16_bits_debugInfo_runahead_checkpoint_id; 
    vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_tlbFirstReqTime <= tr.io_writeback_16_bits_debugInfo_tlbFirstReqTime; 
    vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_tlbRespTime <= tr.io_writeback_16_bits_debugInfo_tlbRespTime; 
    vif.drv_mp.drv_cb.io_writeback_16_bits_debug_seqNum <= tr.io_writeback_16_bits_debug_seqNum; 
    vif.drv_mp.drv_cb.io_writeback_15_valid <= tr.io_writeback_15_valid; 
    vif.drv_mp.drv_cb.io_writeback_15_bits_data_0 <= tr.io_writeback_15_bits_data_0; 
    vif.drv_mp.drv_cb.io_writeback_15_bits_data_1 <= tr.io_writeback_15_bits_data_1; 
    vif.drv_mp.drv_cb.io_writeback_15_bits_data_2 <= tr.io_writeback_15_bits_data_2; 
    vif.drv_mp.drv_cb.io_writeback_15_bits_pdest <= tr.io_writeback_15_bits_pdest; 
    vif.drv_mp.drv_cb.io_writeback_15_bits_robIdx_flag <= tr.io_writeback_15_bits_robIdx_flag; 
    vif.drv_mp.drv_cb.io_writeback_15_bits_robIdx_value <= tr.io_writeback_15_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_writeback_15_bits_vecWen <= tr.io_writeback_15_bits_vecWen; 
    vif.drv_mp.drv_cb.io_writeback_15_bits_v0Wen <= tr.io_writeback_15_bits_v0Wen; 
    vif.drv_mp.drv_cb.io_writeback_15_bits_fflags <= tr.io_writeback_15_bits_fflags; 
    vif.drv_mp.drv_cb.io_writeback_15_bits_wflags <= tr.io_writeback_15_bits_wflags; 
    vif.drv_mp.drv_cb.io_writeback_15_bits_vxsat <= tr.io_writeback_15_bits_vxsat; 
    vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_eliminatedMove <= tr.io_writeback_15_bits_debugInfo_eliminatedMove; 
    vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_renameTime <= tr.io_writeback_15_bits_debugInfo_renameTime; 
    vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_dispatchTime <= tr.io_writeback_15_bits_debugInfo_dispatchTime; 
    vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_enqRsTime <= tr.io_writeback_15_bits_debugInfo_enqRsTime; 
    vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_selectTime <= tr.io_writeback_15_bits_debugInfo_selectTime; 
    vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_issueTime <= tr.io_writeback_15_bits_debugInfo_issueTime; 
    vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_writebackTime <= tr.io_writeback_15_bits_debugInfo_writebackTime; 
    vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_runahead_checkpoint_id <= tr.io_writeback_15_bits_debugInfo_runahead_checkpoint_id; 
    vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_tlbFirstReqTime <= tr.io_writeback_15_bits_debugInfo_tlbFirstReqTime; 
    vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_tlbRespTime <= tr.io_writeback_15_bits_debugInfo_tlbRespTime; 
    vif.drv_mp.drv_cb.io_writeback_15_bits_debug_seqNum <= tr.io_writeback_15_bits_debug_seqNum; 
    vif.drv_mp.drv_cb.io_writeback_14_valid <= tr.io_writeback_14_valid; 
    vif.drv_mp.drv_cb.io_writeback_14_bits_data_0 <= tr.io_writeback_14_bits_data_0; 
    vif.drv_mp.drv_cb.io_writeback_14_bits_data_1 <= tr.io_writeback_14_bits_data_1; 
    vif.drv_mp.drv_cb.io_writeback_14_bits_data_2 <= tr.io_writeback_14_bits_data_2; 
    vif.drv_mp.drv_cb.io_writeback_14_bits_data_3 <= tr.io_writeback_14_bits_data_3; 
    vif.drv_mp.drv_cb.io_writeback_14_bits_data_4 <= tr.io_writeback_14_bits_data_4; 
    vif.drv_mp.drv_cb.io_writeback_14_bits_data_5 <= tr.io_writeback_14_bits_data_5; 
    vif.drv_mp.drv_cb.io_writeback_14_bits_pdest <= tr.io_writeback_14_bits_pdest; 
    vif.drv_mp.drv_cb.io_writeback_14_bits_robIdx_flag <= tr.io_writeback_14_bits_robIdx_flag; 
    vif.drv_mp.drv_cb.io_writeback_14_bits_robIdx_value <= tr.io_writeback_14_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_writeback_14_bits_intWen <= tr.io_writeback_14_bits_intWen; 
    vif.drv_mp.drv_cb.io_writeback_14_bits_fpWen <= tr.io_writeback_14_bits_fpWen; 
    vif.drv_mp.drv_cb.io_writeback_14_bits_vecWen <= tr.io_writeback_14_bits_vecWen; 
    vif.drv_mp.drv_cb.io_writeback_14_bits_v0Wen <= tr.io_writeback_14_bits_v0Wen; 
    vif.drv_mp.drv_cb.io_writeback_14_bits_vlWen <= tr.io_writeback_14_bits_vlWen; 
    vif.drv_mp.drv_cb.io_writeback_14_bits_fflags <= tr.io_writeback_14_bits_fflags; 
    vif.drv_mp.drv_cb.io_writeback_14_bits_wflags <= tr.io_writeback_14_bits_wflags; 
    vif.drv_mp.drv_cb.io_writeback_14_bits_exceptionVec_2 <= tr.io_writeback_14_bits_exceptionVec_2; 
    vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_eliminatedMove <= tr.io_writeback_14_bits_debugInfo_eliminatedMove; 
    vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_renameTime <= tr.io_writeback_14_bits_debugInfo_renameTime; 
    vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_dispatchTime <= tr.io_writeback_14_bits_debugInfo_dispatchTime; 
    vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_enqRsTime <= tr.io_writeback_14_bits_debugInfo_enqRsTime; 
    vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_selectTime <= tr.io_writeback_14_bits_debugInfo_selectTime; 
    vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_issueTime <= tr.io_writeback_14_bits_debugInfo_issueTime; 
    vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_writebackTime <= tr.io_writeback_14_bits_debugInfo_writebackTime; 
    vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_runahead_checkpoint_id <= tr.io_writeback_14_bits_debugInfo_runahead_checkpoint_id; 
    vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_tlbFirstReqTime <= tr.io_writeback_14_bits_debugInfo_tlbFirstReqTime; 
    vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_tlbRespTime <= tr.io_writeback_14_bits_debugInfo_tlbRespTime; 
    vif.drv_mp.drv_cb.io_writeback_14_bits_debug_seqNum <= tr.io_writeback_14_bits_debug_seqNum; 
    vif.drv_mp.drv_cb.io_writeback_13_valid <= tr.io_writeback_13_valid; 
    vif.drv_mp.drv_cb.io_writeback_13_bits_data_0 <= tr.io_writeback_13_bits_data_0; 
    vif.drv_mp.drv_cb.io_writeback_13_bits_data_1 <= tr.io_writeback_13_bits_data_1; 
    vif.drv_mp.drv_cb.io_writeback_13_bits_data_2 <= tr.io_writeback_13_bits_data_2; 
    vif.drv_mp.drv_cb.io_writeback_13_bits_pdest <= tr.io_writeback_13_bits_pdest; 
    vif.drv_mp.drv_cb.io_writeback_13_bits_robIdx_flag <= tr.io_writeback_13_bits_robIdx_flag; 
    vif.drv_mp.drv_cb.io_writeback_13_bits_robIdx_value <= tr.io_writeback_13_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_writeback_13_bits_vecWen <= tr.io_writeback_13_bits_vecWen; 
    vif.drv_mp.drv_cb.io_writeback_13_bits_v0Wen <= tr.io_writeback_13_bits_v0Wen; 
    vif.drv_mp.drv_cb.io_writeback_13_bits_fflags <= tr.io_writeback_13_bits_fflags; 
    vif.drv_mp.drv_cb.io_writeback_13_bits_wflags <= tr.io_writeback_13_bits_wflags; 
    vif.drv_mp.drv_cb.io_writeback_13_bits_vxsat <= tr.io_writeback_13_bits_vxsat; 
    vif.drv_mp.drv_cb.io_writeback_13_bits_exceptionVec_2 <= tr.io_writeback_13_bits_exceptionVec_2; 
    vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_eliminatedMove <= tr.io_writeback_13_bits_debugInfo_eliminatedMove; 
    vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_renameTime <= tr.io_writeback_13_bits_debugInfo_renameTime; 
    vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_dispatchTime <= tr.io_writeback_13_bits_debugInfo_dispatchTime; 
    vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_enqRsTime <= tr.io_writeback_13_bits_debugInfo_enqRsTime; 
    vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_selectTime <= tr.io_writeback_13_bits_debugInfo_selectTime; 
    vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_issueTime <= tr.io_writeback_13_bits_debugInfo_issueTime; 
    vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_writebackTime <= tr.io_writeback_13_bits_debugInfo_writebackTime; 
    vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_runahead_checkpoint_id <= tr.io_writeback_13_bits_debugInfo_runahead_checkpoint_id; 
    vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_tlbFirstReqTime <= tr.io_writeback_13_bits_debugInfo_tlbFirstReqTime; 
    vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_tlbRespTime <= tr.io_writeback_13_bits_debugInfo_tlbRespTime; 
    vif.drv_mp.drv_cb.io_writeback_13_bits_debug_seqNum <= tr.io_writeback_13_bits_debug_seqNum; 
    vif.drv_mp.drv_cb.io_writeback_7_valid <= tr.io_writeback_7_valid; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_data_0 <= tr.io_writeback_7_bits_data_0; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_data_1 <= tr.io_writeback_7_bits_data_1; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_pdest <= tr.io_writeback_7_bits_pdest; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_robIdx_flag <= tr.io_writeback_7_bits_robIdx_flag; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_robIdx_value <= tr.io_writeback_7_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_intWen <= tr.io_writeback_7_bits_intWen; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_valid <= tr.io_writeback_7_bits_redirect_valid; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_isRVC <= tr.io_writeback_7_bits_redirect_bits_isRVC; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_robIdx_flag <= tr.io_writeback_7_bits_redirect_bits_robIdx_flag; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_robIdx_value <= tr.io_writeback_7_bits_redirect_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_ftqIdx_flag <= tr.io_writeback_7_bits_redirect_bits_ftqIdx_flag; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_ftqIdx_value <= tr.io_writeback_7_bits_redirect_bits_ftqIdx_value; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_ftqOffset <= tr.io_writeback_7_bits_redirect_bits_ftqOffset; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_level <= tr.io_writeback_7_bits_redirect_bits_level; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_interrupt <= tr.io_writeback_7_bits_redirect_bits_interrupt; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pc <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_pc; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_ssp <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_ssp; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_sctr <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_sctr; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0 <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1 <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2 <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3 <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0 <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1 <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2 <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3 <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0 <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1 <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2 <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3 <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0 <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1 <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2 <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3 <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0 <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1 <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2 <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3 <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0 <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1 <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2 <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3 <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_ghr <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_ghr; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0 <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1 <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_target <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_target; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_taken <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_taken; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_shift <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_shift; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF <= tr.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_fullTarget <= tr.io_writeback_7_bits_redirect_bits_fullTarget; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_stFtqIdx_flag <= tr.io_writeback_7_bits_redirect_bits_stFtqIdx_flag; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_stFtqIdx_value <= tr.io_writeback_7_bits_redirect_bits_stFtqIdx_value; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_stFtqOffset <= tr.io_writeback_7_bits_redirect_bits_stFtqOffset; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id <= tr.io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_debugIsCtrl <= tr.io_writeback_7_bits_redirect_bits_debugIsCtrl; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_debugIsMemVio <= tr.io_writeback_7_bits_redirect_bits_debugIsMemVio; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_2 <= tr.io_writeback_7_bits_exceptionVec_2; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_3 <= tr.io_writeback_7_bits_exceptionVec_3; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_8 <= tr.io_writeback_7_bits_exceptionVec_8; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_9 <= tr.io_writeback_7_bits_exceptionVec_9; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_10 <= tr.io_writeback_7_bits_exceptionVec_10; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_11 <= tr.io_writeback_7_bits_exceptionVec_11; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_22 <= tr.io_writeback_7_bits_exceptionVec_22; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_flushPipe <= tr.io_writeback_7_bits_flushPipe; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_valid <= tr.io_writeback_7_bits_predecodeInfo_valid; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_isRVC <= tr.io_writeback_7_bits_predecodeInfo_isRVC; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_brType <= tr.io_writeback_7_bits_predecodeInfo_brType; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_isCall <= tr.io_writeback_7_bits_predecodeInfo_isCall; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_isRet <= tr.io_writeback_7_bits_predecodeInfo_isRet; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_debug_isPerfCnt <= tr.io_writeback_7_bits_debug_isPerfCnt; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_eliminatedMove <= tr.io_writeback_7_bits_debugInfo_eliminatedMove; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_renameTime <= tr.io_writeback_7_bits_debugInfo_renameTime; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_dispatchTime <= tr.io_writeback_7_bits_debugInfo_dispatchTime; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_enqRsTime <= tr.io_writeback_7_bits_debugInfo_enqRsTime; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_selectTime <= tr.io_writeback_7_bits_debugInfo_selectTime; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_issueTime <= tr.io_writeback_7_bits_debugInfo_issueTime; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_writebackTime <= tr.io_writeback_7_bits_debugInfo_writebackTime; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_runahead_checkpoint_id <= tr.io_writeback_7_bits_debugInfo_runahead_checkpoint_id; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_tlbFirstReqTime <= tr.io_writeback_7_bits_debugInfo_tlbFirstReqTime; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_tlbRespTime <= tr.io_writeback_7_bits_debugInfo_tlbRespTime; 
    vif.drv_mp.drv_cb.io_writeback_7_bits_debug_seqNum <= tr.io_writeback_7_bits_debug_seqNum; 
    vif.drv_mp.drv_cb.io_writeback_5_valid <= tr.io_writeback_5_valid; 
    vif.drv_mp.drv_cb.io_writeback_5_bits_redirect_valid <= tr.io_writeback_5_bits_redirect_valid; 
    vif.drv_mp.drv_cb.io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred <= tr.io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred; 
    vif.drv_mp.drv_cb.io_writeback_3_valid <= tr.io_writeback_3_valid; 
    vif.drv_mp.drv_cb.io_writeback_3_bits_redirect_valid <= tr.io_writeback_3_bits_redirect_valid; 
    vif.drv_mp.drv_cb.io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred <= tr.io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred; 
    vif.drv_mp.drv_cb.io_writeback_1_valid <= tr.io_writeback_1_valid; 
    vif.drv_mp.drv_cb.io_writeback_1_bits_redirect_valid <= tr.io_writeback_1_bits_redirect_valid; 
    vif.drv_mp.drv_cb.io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred <= tr.io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred; 
    vif.drv_mp.drv_cb.io_exuWriteback_26_valid <= tr.io_exuWriteback_26_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_26_bits_robIdx_value <= tr.io_exuWriteback_26_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_25_valid <= tr.io_exuWriteback_25_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_25_bits_robIdx_value <= tr.io_exuWriteback_25_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_24_valid <= tr.io_exuWriteback_24_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_24_bits_data_0 <= tr.io_exuWriteback_24_bits_data_0; 
    vif.drv_mp.drv_cb.io_exuWriteback_24_bits_pdest <= tr.io_exuWriteback_24_bits_pdest; 
    vif.drv_mp.drv_cb.io_exuWriteback_24_bits_robIdx_value <= tr.io_exuWriteback_24_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_24_bits_vecWen <= tr.io_exuWriteback_24_bits_vecWen; 
    vif.drv_mp.drv_cb.io_exuWriteback_24_bits_v0Wen <= tr.io_exuWriteback_24_bits_v0Wen; 
    vif.drv_mp.drv_cb.io_exuWriteback_24_bits_vls_vdIdx <= tr.io_exuWriteback_24_bits_vls_vdIdx; 
    vif.drv_mp.drv_cb.io_exuWriteback_24_bits_debug_isMMIO <= tr.io_exuWriteback_24_bits_debug_isMMIO; 
    vif.drv_mp.drv_cb.io_exuWriteback_24_bits_debug_isNCIO <= tr.io_exuWriteback_24_bits_debug_isNCIO; 
    vif.drv_mp.drv_cb.io_exuWriteback_24_bits_debug_isPerfCnt <= tr.io_exuWriteback_24_bits_debug_isPerfCnt; 
    vif.drv_mp.drv_cb.io_exuWriteback_24_bits_debug_paddr <= tr.io_exuWriteback_24_bits_debug_paddr; 
    vif.drv_mp.drv_cb.io_exuWriteback_23_valid <= tr.io_exuWriteback_23_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_23_bits_data_0 <= tr.io_exuWriteback_23_bits_data_0; 
    vif.drv_mp.drv_cb.io_exuWriteback_23_bits_pdest <= tr.io_exuWriteback_23_bits_pdest; 
    vif.drv_mp.drv_cb.io_exuWriteback_23_bits_robIdx_value <= tr.io_exuWriteback_23_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_23_bits_vecWen <= tr.io_exuWriteback_23_bits_vecWen; 
    vif.drv_mp.drv_cb.io_exuWriteback_23_bits_v0Wen <= tr.io_exuWriteback_23_bits_v0Wen; 
    vif.drv_mp.drv_cb.io_exuWriteback_23_bits_vls_vdIdx <= tr.io_exuWriteback_23_bits_vls_vdIdx; 
    vif.drv_mp.drv_cb.io_exuWriteback_23_bits_debug_isMMIO <= tr.io_exuWriteback_23_bits_debug_isMMIO; 
    vif.drv_mp.drv_cb.io_exuWriteback_23_bits_debug_isNCIO <= tr.io_exuWriteback_23_bits_debug_isNCIO; 
    vif.drv_mp.drv_cb.io_exuWriteback_23_bits_debug_isPerfCnt <= tr.io_exuWriteback_23_bits_debug_isPerfCnt; 
    vif.drv_mp.drv_cb.io_exuWriteback_23_bits_debug_paddr <= tr.io_exuWriteback_23_bits_debug_paddr; 
    vif.drv_mp.drv_cb.io_exuWriteback_22_valid <= tr.io_exuWriteback_22_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_22_bits_data_0 <= tr.io_exuWriteback_22_bits_data_0; 
    vif.drv_mp.drv_cb.io_exuWriteback_22_bits_robIdx_value <= tr.io_exuWriteback_22_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_22_bits_lqIdx_value <= tr.io_exuWriteback_22_bits_lqIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_22_bits_debug_isMMIO <= tr.io_exuWriteback_22_bits_debug_isMMIO; 
    vif.drv_mp.drv_cb.io_exuWriteback_22_bits_debug_isNCIO <= tr.io_exuWriteback_22_bits_debug_isNCIO; 
    vif.drv_mp.drv_cb.io_exuWriteback_22_bits_debug_isPerfCnt <= tr.io_exuWriteback_22_bits_debug_isPerfCnt; 
    vif.drv_mp.drv_cb.io_exuWriteback_22_bits_debug_paddr <= tr.io_exuWriteback_22_bits_debug_paddr; 
    vif.drv_mp.drv_cb.io_exuWriteback_21_valid <= tr.io_exuWriteback_21_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_21_bits_data_0 <= tr.io_exuWriteback_21_bits_data_0; 
    vif.drv_mp.drv_cb.io_exuWriteback_21_bits_robIdx_value <= tr.io_exuWriteback_21_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_21_bits_lqIdx_value <= tr.io_exuWriteback_21_bits_lqIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_21_bits_debug_isMMIO <= tr.io_exuWriteback_21_bits_debug_isMMIO; 
    vif.drv_mp.drv_cb.io_exuWriteback_21_bits_debug_isNCIO <= tr.io_exuWriteback_21_bits_debug_isNCIO; 
    vif.drv_mp.drv_cb.io_exuWriteback_21_bits_debug_isPerfCnt <= tr.io_exuWriteback_21_bits_debug_isPerfCnt; 
    vif.drv_mp.drv_cb.io_exuWriteback_21_bits_debug_paddr <= tr.io_exuWriteback_21_bits_debug_paddr; 
    vif.drv_mp.drv_cb.io_exuWriteback_20_valid <= tr.io_exuWriteback_20_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_20_bits_data_0 <= tr.io_exuWriteback_20_bits_data_0; 
    vif.drv_mp.drv_cb.io_exuWriteback_20_bits_robIdx_value <= tr.io_exuWriteback_20_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_20_bits_lqIdx_value <= tr.io_exuWriteback_20_bits_lqIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_20_bits_debug_isMMIO <= tr.io_exuWriteback_20_bits_debug_isMMIO; 
    vif.drv_mp.drv_cb.io_exuWriteback_20_bits_debug_isNCIO <= tr.io_exuWriteback_20_bits_debug_isNCIO; 
    vif.drv_mp.drv_cb.io_exuWriteback_20_bits_debug_isPerfCnt <= tr.io_exuWriteback_20_bits_debug_isPerfCnt; 
    vif.drv_mp.drv_cb.io_exuWriteback_20_bits_debug_paddr <= tr.io_exuWriteback_20_bits_debug_paddr; 
    vif.drv_mp.drv_cb.io_exuWriteback_19_valid <= tr.io_exuWriteback_19_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_19_bits_data_0 <= tr.io_exuWriteback_19_bits_data_0; 
    vif.drv_mp.drv_cb.io_exuWriteback_19_bits_robIdx_value <= tr.io_exuWriteback_19_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_19_bits_sqIdx_value <= tr.io_exuWriteback_19_bits_sqIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_19_bits_debug_isMMIO <= tr.io_exuWriteback_19_bits_debug_isMMIO; 
    vif.drv_mp.drv_cb.io_exuWriteback_19_bits_debug_isNCIO <= tr.io_exuWriteback_19_bits_debug_isNCIO; 
    vif.drv_mp.drv_cb.io_exuWriteback_19_bits_debug_isPerfCnt <= tr.io_exuWriteback_19_bits_debug_isPerfCnt; 
    vif.drv_mp.drv_cb.io_exuWriteback_19_bits_debug_paddr <= tr.io_exuWriteback_19_bits_debug_paddr; 
    vif.drv_mp.drv_cb.io_exuWriteback_18_valid <= tr.io_exuWriteback_18_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_18_bits_data_0 <= tr.io_exuWriteback_18_bits_data_0; 
    vif.drv_mp.drv_cb.io_exuWriteback_18_bits_robIdx_value <= tr.io_exuWriteback_18_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_18_bits_sqIdx_value <= tr.io_exuWriteback_18_bits_sqIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_18_bits_debug_isMMIO <= tr.io_exuWriteback_18_bits_debug_isMMIO; 
    vif.drv_mp.drv_cb.io_exuWriteback_18_bits_debug_isNCIO <= tr.io_exuWriteback_18_bits_debug_isNCIO; 
    vif.drv_mp.drv_cb.io_exuWriteback_18_bits_debug_isPerfCnt <= tr.io_exuWriteback_18_bits_debug_isPerfCnt; 
    vif.drv_mp.drv_cb.io_exuWriteback_18_bits_debug_paddr <= tr.io_exuWriteback_18_bits_debug_paddr; 
    vif.drv_mp.drv_cb.io_exuWriteback_17_valid <= tr.io_exuWriteback_17_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_17_bits_data_0 <= tr.io_exuWriteback_17_bits_data_0; 
    vif.drv_mp.drv_cb.io_exuWriteback_17_bits_robIdx_value <= tr.io_exuWriteback_17_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_17_bits_fflags <= tr.io_exuWriteback_17_bits_fflags; 
    vif.drv_mp.drv_cb.io_exuWriteback_17_bits_wflags <= tr.io_exuWriteback_17_bits_wflags; 
    vif.drv_mp.drv_cb.io_exuWriteback_16_valid <= tr.io_exuWriteback_16_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_16_bits_data_0 <= tr.io_exuWriteback_16_bits_data_0; 
    vif.drv_mp.drv_cb.io_exuWriteback_16_bits_robIdx_value <= tr.io_exuWriteback_16_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_16_bits_fflags <= tr.io_exuWriteback_16_bits_fflags; 
    vif.drv_mp.drv_cb.io_exuWriteback_16_bits_wflags <= tr.io_exuWriteback_16_bits_wflags; 
    vif.drv_mp.drv_cb.io_exuWriteback_15_valid <= tr.io_exuWriteback_15_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_15_bits_data_0 <= tr.io_exuWriteback_15_bits_data_0; 
    vif.drv_mp.drv_cb.io_exuWriteback_15_bits_robIdx_value <= tr.io_exuWriteback_15_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_15_bits_fflags <= tr.io_exuWriteback_15_bits_fflags; 
    vif.drv_mp.drv_cb.io_exuWriteback_15_bits_wflags <= tr.io_exuWriteback_15_bits_wflags; 
    vif.drv_mp.drv_cb.io_exuWriteback_15_bits_vxsat <= tr.io_exuWriteback_15_bits_vxsat; 
    vif.drv_mp.drv_cb.io_exuWriteback_14_valid <= tr.io_exuWriteback_14_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_14_bits_data_0 <= tr.io_exuWriteback_14_bits_data_0; 
    vif.drv_mp.drv_cb.io_exuWriteback_14_bits_robIdx_value <= tr.io_exuWriteback_14_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_14_bits_fflags <= tr.io_exuWriteback_14_bits_fflags; 
    vif.drv_mp.drv_cb.io_exuWriteback_14_bits_wflags <= tr.io_exuWriteback_14_bits_wflags; 
    vif.drv_mp.drv_cb.io_exuWriteback_13_valid <= tr.io_exuWriteback_13_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_13_bits_data_0 <= tr.io_exuWriteback_13_bits_data_0; 
    vif.drv_mp.drv_cb.io_exuWriteback_13_bits_robIdx_value <= tr.io_exuWriteback_13_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_13_bits_fflags <= tr.io_exuWriteback_13_bits_fflags; 
    vif.drv_mp.drv_cb.io_exuWriteback_13_bits_wflags <= tr.io_exuWriteback_13_bits_wflags; 
    vif.drv_mp.drv_cb.io_exuWriteback_13_bits_vxsat <= tr.io_exuWriteback_13_bits_vxsat; 
    vif.drv_mp.drv_cb.io_exuWriteback_12_valid <= tr.io_exuWriteback_12_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_12_bits_data_0 <= tr.io_exuWriteback_12_bits_data_0; 
    vif.drv_mp.drv_cb.io_exuWriteback_12_bits_robIdx_value <= tr.io_exuWriteback_12_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_12_bits_fflags <= tr.io_exuWriteback_12_bits_fflags; 
    vif.drv_mp.drv_cb.io_exuWriteback_12_bits_wflags <= tr.io_exuWriteback_12_bits_wflags; 
    vif.drv_mp.drv_cb.io_exuWriteback_11_valid <= tr.io_exuWriteback_11_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_11_bits_data_0 <= tr.io_exuWriteback_11_bits_data_0; 
    vif.drv_mp.drv_cb.io_exuWriteback_11_bits_robIdx_value <= tr.io_exuWriteback_11_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_11_bits_fflags <= tr.io_exuWriteback_11_bits_fflags; 
    vif.drv_mp.drv_cb.io_exuWriteback_11_bits_wflags <= tr.io_exuWriteback_11_bits_wflags; 
    vif.drv_mp.drv_cb.io_exuWriteback_10_valid <= tr.io_exuWriteback_10_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_10_bits_data_0 <= tr.io_exuWriteback_10_bits_data_0; 
    vif.drv_mp.drv_cb.io_exuWriteback_10_bits_robIdx_value <= tr.io_exuWriteback_10_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_10_bits_fflags <= tr.io_exuWriteback_10_bits_fflags; 
    vif.drv_mp.drv_cb.io_exuWriteback_10_bits_wflags <= tr.io_exuWriteback_10_bits_wflags; 
    vif.drv_mp.drv_cb.io_exuWriteback_9_valid <= tr.io_exuWriteback_9_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_9_bits_data_0 <= tr.io_exuWriteback_9_bits_data_0; 
    vif.drv_mp.drv_cb.io_exuWriteback_9_bits_robIdx_value <= tr.io_exuWriteback_9_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_9_bits_fflags <= tr.io_exuWriteback_9_bits_fflags; 
    vif.drv_mp.drv_cb.io_exuWriteback_9_bits_wflags <= tr.io_exuWriteback_9_bits_wflags; 
    vif.drv_mp.drv_cb.io_exuWriteback_8_valid <= tr.io_exuWriteback_8_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_8_bits_data_0 <= tr.io_exuWriteback_8_bits_data_0; 
    vif.drv_mp.drv_cb.io_exuWriteback_8_bits_robIdx_value <= tr.io_exuWriteback_8_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_8_bits_fflags <= tr.io_exuWriteback_8_bits_fflags; 
    vif.drv_mp.drv_cb.io_exuWriteback_8_bits_wflags <= tr.io_exuWriteback_8_bits_wflags; 
    vif.drv_mp.drv_cb.io_exuWriteback_7_valid <= tr.io_exuWriteback_7_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_7_bits_data_0 <= tr.io_exuWriteback_7_bits_data_0; 
    vif.drv_mp.drv_cb.io_exuWriteback_7_bits_robIdx_value <= tr.io_exuWriteback_7_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_7_bits_debug_isPerfCnt <= tr.io_exuWriteback_7_bits_debug_isPerfCnt; 
    vif.drv_mp.drv_cb.io_exuWriteback_6_valid <= tr.io_exuWriteback_6_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_6_bits_data_0 <= tr.io_exuWriteback_6_bits_data_0; 
    vif.drv_mp.drv_cb.io_exuWriteback_6_bits_robIdx_value <= tr.io_exuWriteback_6_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_5_valid <= tr.io_exuWriteback_5_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_5_bits_data_0 <= tr.io_exuWriteback_5_bits_data_0; 
    vif.drv_mp.drv_cb.io_exuWriteback_5_bits_robIdx_value <= tr.io_exuWriteback_5_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_5_bits_redirect_valid <= tr.io_exuWriteback_5_bits_redirect_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken <= tr.io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken; 
    vif.drv_mp.drv_cb.io_exuWriteback_5_bits_fflags <= tr.io_exuWriteback_5_bits_fflags; 
    vif.drv_mp.drv_cb.io_exuWriteback_5_bits_wflags <= tr.io_exuWriteback_5_bits_wflags; 
    vif.drv_mp.drv_cb.io_exuWriteback_4_valid <= tr.io_exuWriteback_4_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_4_bits_data_0 <= tr.io_exuWriteback_4_bits_data_0; 
    vif.drv_mp.drv_cb.io_exuWriteback_4_bits_robIdx_value <= tr.io_exuWriteback_4_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_3_valid <= tr.io_exuWriteback_3_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_3_bits_data_0 <= tr.io_exuWriteback_3_bits_data_0; 
    vif.drv_mp.drv_cb.io_exuWriteback_3_bits_robIdx_value <= tr.io_exuWriteback_3_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_3_bits_redirect_valid <= tr.io_exuWriteback_3_bits_redirect_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken <= tr.io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken; 
    vif.drv_mp.drv_cb.io_exuWriteback_2_valid <= tr.io_exuWriteback_2_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_2_bits_data_0 <= tr.io_exuWriteback_2_bits_data_0; 
    vif.drv_mp.drv_cb.io_exuWriteback_2_bits_robIdx_value <= tr.io_exuWriteback_2_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_1_valid <= tr.io_exuWriteback_1_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_1_bits_data_0 <= tr.io_exuWriteback_1_bits_data_0; 
    vif.drv_mp.drv_cb.io_exuWriteback_1_bits_robIdx_value <= tr.io_exuWriteback_1_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_exuWriteback_1_bits_redirect_valid <= tr.io_exuWriteback_1_bits_redirect_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken <= tr.io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken; 
    vif.drv_mp.drv_cb.io_exuWriteback_0_valid <= tr.io_exuWriteback_0_valid; 
    vif.drv_mp.drv_cb.io_exuWriteback_0_bits_data_0 <= tr.io_exuWriteback_0_bits_data_0; 
    vif.drv_mp.drv_cb.io_exuWriteback_0_bits_robIdx_value <= tr.io_exuWriteback_0_bits_robIdx_value; 
    vif.drv_mp.drv_cb.io_writebackNums_0_bits <= tr.io_writebackNums_0_bits; 
    vif.drv_mp.drv_cb.io_writebackNums_1_bits <= tr.io_writebackNums_1_bits; 
    vif.drv_mp.drv_cb.io_writebackNums_2_bits <= tr.io_writebackNums_2_bits; 
    vif.drv_mp.drv_cb.io_writebackNums_3_bits <= tr.io_writebackNums_3_bits; 
    vif.drv_mp.drv_cb.io_writebackNums_4_bits <= tr.io_writebackNums_4_bits; 
    vif.drv_mp.drv_cb.io_writebackNums_5_bits <= tr.io_writebackNums_5_bits; 
    vif.drv_mp.drv_cb.io_writebackNums_6_bits <= tr.io_writebackNums_6_bits; 
    vif.drv_mp.drv_cb.io_writebackNums_7_bits <= tr.io_writebackNums_7_bits; 
    vif.drv_mp.drv_cb.io_writebackNums_8_bits <= tr.io_writebackNums_8_bits; 
    vif.drv_mp.drv_cb.io_writebackNums_9_bits <= tr.io_writebackNums_9_bits; 
    vif.drv_mp.drv_cb.io_writebackNums_10_bits <= tr.io_writebackNums_10_bits; 
    vif.drv_mp.drv_cb.io_writebackNums_11_bits <= tr.io_writebackNums_11_bits; 
    vif.drv_mp.drv_cb.io_writebackNums_12_bits <= tr.io_writebackNums_12_bits; 
    vif.drv_mp.drv_cb.io_writebackNums_13_bits <= tr.io_writebackNums_13_bits; 
    vif.drv_mp.drv_cb.io_writebackNums_14_bits <= tr.io_writebackNums_14_bits; 
    vif.drv_mp.drv_cb.io_writebackNums_15_bits <= tr.io_writebackNums_15_bits; 
    vif.drv_mp.drv_cb.io_writebackNums_16_bits <= tr.io_writebackNums_16_bits; 
    vif.drv_mp.drv_cb.io_writebackNums_17_bits <= tr.io_writebackNums_17_bits; 
    vif.drv_mp.drv_cb.io_writebackNums_18_bits <= tr.io_writebackNums_18_bits; 
    vif.drv_mp.drv_cb.io_writebackNums_19_bits <= tr.io_writebackNums_19_bits; 
    vif.drv_mp.drv_cb.io_writebackNums_20_bits <= tr.io_writebackNums_20_bits; 
    vif.drv_mp.drv_cb.io_writebackNums_21_bits <= tr.io_writebackNums_21_bits; 
    vif.drv_mp.drv_cb.io_writebackNums_22_bits <= tr.io_writebackNums_22_bits; 
    vif.drv_mp.drv_cb.io_writebackNums_23_bits <= tr.io_writebackNums_23_bits; 
    vif.drv_mp.drv_cb.io_writebackNums_24_bits <= tr.io_writebackNums_24_bits; 
    vif.drv_mp.drv_cb.io_writebackNeedFlush_0 <= tr.io_writebackNeedFlush_0; 
    vif.drv_mp.drv_cb.io_writebackNeedFlush_1 <= tr.io_writebackNeedFlush_1; 
    vif.drv_mp.drv_cb.io_writebackNeedFlush_2 <= tr.io_writebackNeedFlush_2; 
    vif.drv_mp.drv_cb.io_writebackNeedFlush_6 <= tr.io_writebackNeedFlush_6; 
    vif.drv_mp.drv_cb.io_writebackNeedFlush_7 <= tr.io_writebackNeedFlush_7; 
    vif.drv_mp.drv_cb.io_writebackNeedFlush_8 <= tr.io_writebackNeedFlush_8; 
    vif.drv_mp.drv_cb.io_writebackNeedFlush_9 <= tr.io_writebackNeedFlush_9; 
    vif.drv_mp.drv_cb.io_writebackNeedFlush_10 <= tr.io_writebackNeedFlush_10; 
    vif.drv_mp.drv_cb.io_writebackNeedFlush_11 <= tr.io_writebackNeedFlush_11; 
    vif.drv_mp.drv_cb.io_writebackNeedFlush_12 <= tr.io_writebackNeedFlush_12; 

endtask:send_pkt

task WriteBack_in_agent_driver::drive_idle(tcnt_dec_base::drv_mode_e drv_mode);

    if(drv_mode==tcnt_dec_base::DRV_0) begin
        vif.drv_mp.drv_cb.io_writeback_24_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vlWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_4 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_5 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_6 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_7 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_8 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_9 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_10 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_11 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_12 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_13 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_14 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_15 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_16 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_17 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_18 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_19 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_20 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_21 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_22 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_23 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_flushPipe <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_replay <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_trigger <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vill <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vma <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vta <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vsew <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vlmul <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVill <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVma <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVta <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVsew <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVlmul <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vm <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vstart <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_frm <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFP32Instr <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFP64Instr <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isReduction <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vxrm <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vuopIdx <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_lastUop <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vmask <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vl <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_nf <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_veew <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isReverse <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isExt <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isNarrow <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isDstMask <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isOpMask <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isDependOldVd <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isWritePartVd <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isVleff <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_oldVdPsrc <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vdIdx <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vdIdxInField <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isIndexed <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isMasked <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isStrided <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isWhole <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isVecLoad <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isVlm <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_isMMIO <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_isNCIO <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_paddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_vaddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_renameTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_dispatchTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_enqRsTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_selectTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_issueTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_writebackTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_runahead_checkpoint_id <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_tlbFirstReqTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_tlbRespTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_seqNum <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vlWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_4 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_5 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_6 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_7 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_8 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_9 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_10 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_11 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_12 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_13 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_14 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_15 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_16 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_17 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_18 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_19 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_20 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_21 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_22 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_23 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_flushPipe <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_replay <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_trigger <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vill <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vma <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vta <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vsew <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vlmul <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVill <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVma <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVta <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVsew <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVlmul <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vm <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vstart <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_frm <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFP32Instr <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFP64Instr <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isReduction <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vxrm <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vuopIdx <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_lastUop <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vmask <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vl <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_nf <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_veew <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isReverse <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isExt <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isNarrow <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isDstMask <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isOpMask <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isDependOldVd <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isWritePartVd <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isVleff <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_oldVdPsrc <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vdIdx <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vdIdxInField <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isIndexed <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isMasked <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isStrided <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isWhole <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isVecLoad <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isVlm <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_isMMIO <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_isNCIO <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_paddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_vaddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_renameTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_dispatchTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_enqRsTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_selectTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_issueTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_writebackTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_runahead_checkpoint_id <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_tlbFirstReqTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_tlbRespTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_seqNum <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_intWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_fpWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_4 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_5 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_6 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_7 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_8 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_9 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_10 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_11 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_12 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_13 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_14 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_15 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_16 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_17 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_18 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_19 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_20 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_21 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_22 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_23 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_flushPipe <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_replay <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_lqIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_lqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_trigger <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_isRVC <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_brType <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_isCall <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_isRet <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_isMMIO <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_isNCIO <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_paddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_vaddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_renameTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_dispatchTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_enqRsTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_selectTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_issueTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_writebackTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_runahead_checkpoint_id <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_tlbFirstReqTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_tlbRespTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_seqNum <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_intWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_fpWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_4 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_5 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_6 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_7 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_8 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_9 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_10 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_11 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_12 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_13 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_14 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_15 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_16 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_17 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_18 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_19 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_20 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_21 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_22 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_23 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_flushPipe <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_replay <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_lqIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_lqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_trigger <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_isRVC <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_brType <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_isCall <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_isRet <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_isMMIO <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_isNCIO <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_paddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_vaddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_renameTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_dispatchTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_enqRsTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_selectTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_issueTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_writebackTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_runahead_checkpoint_id <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_tlbFirstReqTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_tlbRespTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_seqNum <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_intWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_fpWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_4 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_5 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_6 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_7 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_8 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_9 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_10 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_11 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_12 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_13 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_14 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_15 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_16 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_17 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_18 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_19 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_20 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_21 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_22 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_23 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_flushPipe <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_replay <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_lqIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_lqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_trigger <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_isRVC <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_brType <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_isCall <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_isRet <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_isMMIO <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_isNCIO <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_paddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_vaddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_renameTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_dispatchTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_enqRsTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_selectTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_issueTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_writebackTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_runahead_checkpoint_id <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_tlbFirstReqTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_tlbRespTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_seqNum <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_intWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_4 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_5 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_6 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_7 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_8 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_9 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_10 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_11 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_12 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_13 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_14 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_15 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_16 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_17 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_18 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_19 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_20 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_21 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_22 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_23 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_flushPipe <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_sqIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_sqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_trigger <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_isMMIO <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_isNCIO <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_paddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_vaddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_renameTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_dispatchTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_enqRsTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_selectTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_issueTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_writebackTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_runahead_checkpoint_id <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_tlbFirstReqTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_tlbRespTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_seqNum <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_intWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_4 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_5 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_6 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_7 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_8 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_9 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_10 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_11 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_12 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_13 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_14 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_15 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_16 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_17 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_18 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_19 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_20 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_21 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_22 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_23 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_flushPipe <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_sqIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_sqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_trigger <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_isMMIO <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_isNCIO <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_paddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_vaddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_renameTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_dispatchTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_enqRsTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_selectTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_issueTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_writebackTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_runahead_checkpoint_id <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_tlbFirstReqTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_tlbRespTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_seqNum <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_data_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_data_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_renameTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_dispatchTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_enqRsTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_selectTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_issueTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_writebackTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_runahead_checkpoint_id <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_tlbFirstReqTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_tlbRespTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debug_seqNum <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_data_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_data_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_data_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_fpWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_renameTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_dispatchTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_enqRsTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_selectTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_issueTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_writebackTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_runahead_checkpoint_id <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_tlbFirstReqTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_tlbRespTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debug_seqNum <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_data_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_data_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_vxsat <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_renameTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_dispatchTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_enqRsTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_selectTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_issueTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_writebackTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_runahead_checkpoint_id <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_tlbFirstReqTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_tlbRespTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debug_seqNum <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_4 <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_5 <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_intWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_fpWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_vlWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_renameTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_dispatchTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_enqRsTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_selectTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_issueTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_writebackTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_runahead_checkpoint_id <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_tlbFirstReqTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_tlbRespTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debug_seqNum <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_data_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_data_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_vxsat <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_renameTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_dispatchTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_enqRsTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_selectTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_issueTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_writebackTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_runahead_checkpoint_id <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_tlbFirstReqTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_tlbRespTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debug_seqNum <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_data_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_intWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_isRVC <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_ftqIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_ftqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_ftqOffset <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_level <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_interrupt <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pc <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_ssp <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_sctr <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_ghr <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_target <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_taken <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_shift <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_fullTarget <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_stFtqIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_stFtqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_stFtqOffset <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_debugIsCtrl <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_debugIsMemVio <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_8 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_9 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_10 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_11 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_22 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_flushPipe <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_isRVC <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_brType <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_isCall <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_isRet <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_renameTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_dispatchTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_enqRsTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_selectTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_issueTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_writebackTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_runahead_checkpoint_id <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_tlbFirstReqTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_tlbRespTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debug_seqNum <= '0;
        vif.drv_mp.drv_cb.io_writeback_5_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_5_bits_redirect_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred <= '0;
        vif.drv_mp.drv_cb.io_writeback_3_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_3_bits_redirect_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred <= '0;
        vif.drv_mp.drv_cb.io_writeback_1_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_1_bits_redirect_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_26_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_26_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_25_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_25_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_24_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_vls_vdIdx <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_debug_isMMIO <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_debug_isNCIO <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_debug_paddr <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_23_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_vls_vdIdx <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_debug_isMMIO <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_debug_isNCIO <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_debug_paddr <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_22_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_lqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_debug_isMMIO <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_debug_isNCIO <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_debug_paddr <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_21_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_lqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_debug_isMMIO <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_debug_isNCIO <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_debug_paddr <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_20_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_lqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_debug_isMMIO <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_debug_isNCIO <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_debug_paddr <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_19_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_sqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_debug_isMMIO <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_debug_isNCIO <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_debug_paddr <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_18_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_sqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_debug_isMMIO <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_debug_isNCIO <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_debug_paddr <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_17_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_17_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_17_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_17_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_17_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_16_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_16_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_16_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_16_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_16_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_15_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_15_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_15_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_15_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_15_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_15_bits_vxsat <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_14_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_14_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_14_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_14_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_14_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_13_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_13_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_13_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_13_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_13_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_13_bits_vxsat <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_12_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_12_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_12_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_12_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_12_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_11_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_11_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_11_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_11_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_11_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_10_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_10_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_10_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_10_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_10_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_9_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_9_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_9_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_9_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_9_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_8_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_8_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_8_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_8_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_8_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_7_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_7_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_7_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_7_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_6_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_6_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_6_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_5_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_redirect_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_4_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_4_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_4_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_3_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_3_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_3_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_3_bits_redirect_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_2_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_2_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_2_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_1_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_1_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_1_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_1_bits_redirect_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_0_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_0_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_0_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_0_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_1_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_2_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_3_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_4_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_5_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_6_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_7_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_8_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_9_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_10_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_11_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_12_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_13_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_14_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_15_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_16_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_17_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_18_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_19_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_20_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_21_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_22_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_23_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_24_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_0 <= '0;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_1 <= '0;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_2 <= '0;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_6 <= '0;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_7 <= '0;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_8 <= '0;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_9 <= '0;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_10 <= '0;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_11 <= '0;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_12 <= '0;

    end
    else if(drv_mode==tcnt_dec_base::DRV_1) begin
        vif.drv_mp.drv_cb.io_writeback_24_valid <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_pdest <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_robIdx_flag <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vecWen <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_v0Wen <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vlWen <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_0 <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_1 <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_2 <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_3 <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_4 <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_5 <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_6 <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_7 <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_8 <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_9 <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_10 <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_11 <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_12 <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_13 <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_14 <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_15 <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_16 <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_17 <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_18 <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_19 <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_20 <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_21 <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_22 <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_23 <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_flushPipe <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_replay <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_trigger <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vill <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vma <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vta <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vsew <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vlmul <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVill <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVma <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVta <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVsew <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVlmul <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vm <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vstart <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_frm <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFP32Instr <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFP64Instr <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isReduction <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2 <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4 <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8 <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vxrm <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vuopIdx <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_lastUop <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vmask <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vl <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_nf <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_veew <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isReverse <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isExt <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isNarrow <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isDstMask <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isOpMask <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isMove <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isDependOldVd <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isWritePartVd <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isVleff <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_oldVdPsrc <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vdIdx <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vdIdxInField <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isIndexed <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isMasked <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isStrided <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isWhole <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isVecLoad <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isVlm <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_isMMIO <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_isNCIO <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_isPerfCnt <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_paddr <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_vaddr <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_eliminatedMove <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_renameTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_dispatchTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_enqRsTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_selectTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_issueTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_writebackTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_runahead_checkpoint_id <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_tlbFirstReqTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_tlbRespTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_seqNum <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_valid <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_pdest <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_robIdx_flag <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vecWen <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_v0Wen <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vlWen <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_0 <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_1 <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_2 <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_3 <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_4 <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_5 <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_6 <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_7 <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_8 <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_9 <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_10 <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_11 <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_12 <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_13 <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_14 <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_15 <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_16 <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_17 <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_18 <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_19 <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_20 <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_21 <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_22 <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_23 <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_flushPipe <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_replay <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_trigger <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vill <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vma <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vta <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vsew <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vlmul <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVill <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVma <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVta <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVsew <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVlmul <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vm <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vstart <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_frm <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFP32Instr <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFP64Instr <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isReduction <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2 <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4 <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8 <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vxrm <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vuopIdx <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_lastUop <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vmask <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vl <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_nf <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_veew <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isReverse <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isExt <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isNarrow <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isDstMask <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isOpMask <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isMove <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isDependOldVd <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isWritePartVd <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isVleff <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_oldVdPsrc <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vdIdx <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vdIdxInField <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isIndexed <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isMasked <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isStrided <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isWhole <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isVecLoad <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isVlm <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_isMMIO <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_isNCIO <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_isPerfCnt <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_paddr <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_vaddr <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_eliminatedMove <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_renameTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_dispatchTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_enqRsTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_selectTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_issueTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_writebackTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_runahead_checkpoint_id <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_tlbFirstReqTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_tlbRespTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_seqNum <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_valid <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_pdest <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_robIdx_flag <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_intWen <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_fpWen <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_0 <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_1 <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_2 <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_3 <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_4 <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_5 <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_6 <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_7 <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_8 <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_9 <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_10 <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_11 <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_12 <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_13 <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_14 <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_15 <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_16 <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_17 <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_18 <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_19 <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_20 <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_21 <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_22 <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_23 <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_flushPipe <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_replay <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_lqIdx_flag <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_lqIdx_value <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_trigger <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_valid <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_isRVC <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_brType <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_isCall <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_isRet <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_isMMIO <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_isNCIO <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_isPerfCnt <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_paddr <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_vaddr <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_eliminatedMove <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_renameTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_dispatchTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_enqRsTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_selectTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_issueTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_writebackTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_runahead_checkpoint_id <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_tlbFirstReqTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_tlbRespTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_seqNum <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_valid <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_pdest <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_robIdx_flag <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_intWen <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_fpWen <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_0 <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_1 <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_2 <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_3 <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_4 <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_5 <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_6 <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_7 <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_8 <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_9 <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_10 <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_11 <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_12 <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_13 <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_14 <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_15 <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_16 <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_17 <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_18 <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_19 <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_20 <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_21 <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_22 <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_23 <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_flushPipe <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_replay <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_lqIdx_flag <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_lqIdx_value <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_trigger <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_valid <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_isRVC <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_brType <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_isCall <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_isRet <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_isMMIO <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_isNCIO <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_isPerfCnt <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_paddr <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_vaddr <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_eliminatedMove <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_renameTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_dispatchTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_enqRsTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_selectTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_issueTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_writebackTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_runahead_checkpoint_id <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_tlbFirstReqTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_tlbRespTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_seqNum <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_valid <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_pdest <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_robIdx_flag <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_intWen <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_fpWen <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_0 <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_1 <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_2 <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_3 <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_4 <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_5 <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_6 <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_7 <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_8 <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_9 <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_10 <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_11 <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_12 <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_13 <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_14 <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_15 <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_16 <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_17 <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_18 <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_19 <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_20 <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_21 <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_22 <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_23 <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_flushPipe <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_replay <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_lqIdx_flag <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_lqIdx_value <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_trigger <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_valid <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_isRVC <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_brType <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_isCall <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_isRet <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_isMMIO <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_isNCIO <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_isPerfCnt <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_paddr <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_vaddr <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_eliminatedMove <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_renameTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_dispatchTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_enqRsTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_selectTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_issueTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_writebackTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_runahead_checkpoint_id <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_tlbFirstReqTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_tlbRespTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_seqNum <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_valid <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_pdest <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_robIdx_flag <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_intWen <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_0 <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_1 <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_2 <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_3 <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_4 <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_5 <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_6 <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_7 <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_8 <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_9 <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_10 <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_11 <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_12 <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_13 <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_14 <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_15 <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_16 <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_17 <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_18 <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_19 <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_20 <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_21 <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_22 <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_23 <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_flushPipe <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_sqIdx_flag <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_sqIdx_value <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_trigger <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_isMMIO <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_isNCIO <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_isPerfCnt <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_paddr <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_vaddr <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_eliminatedMove <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_renameTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_dispatchTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_enqRsTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_selectTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_issueTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_writebackTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_runahead_checkpoint_id <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_tlbFirstReqTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_tlbRespTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_seqNum <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_valid <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_pdest <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_robIdx_flag <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_intWen <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_0 <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_1 <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_2 <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_3 <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_4 <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_5 <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_6 <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_7 <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_8 <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_9 <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_10 <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_11 <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_12 <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_13 <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_14 <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_15 <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_16 <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_17 <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_18 <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_19 <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_20 <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_21 <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_22 <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_23 <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_flushPipe <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_sqIdx_flag <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_sqIdx_value <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_trigger <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_isMMIO <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_isNCIO <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_isPerfCnt <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_paddr <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_vaddr <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_eliminatedMove <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_renameTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_dispatchTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_enqRsTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_selectTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_issueTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_writebackTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_runahead_checkpoint_id <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_tlbFirstReqTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_tlbRespTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_seqNum <= '1;
        vif.drv_mp.drv_cb.io_writeback_17_valid <= '1;
        vif.drv_mp.drv_cb.io_writeback_17_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_writeback_17_bits_data_1 <= '1;
        vif.drv_mp.drv_cb.io_writeback_17_bits_data_2 <= '1;
        vif.drv_mp.drv_cb.io_writeback_17_bits_pdest <= '1;
        vif.drv_mp.drv_cb.io_writeback_17_bits_robIdx_flag <= '1;
        vif.drv_mp.drv_cb.io_writeback_17_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_writeback_17_bits_vecWen <= '1;
        vif.drv_mp.drv_cb.io_writeback_17_bits_v0Wen <= '1;
        vif.drv_mp.drv_cb.io_writeback_17_bits_fflags <= '1;
        vif.drv_mp.drv_cb.io_writeback_17_bits_wflags <= '1;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_eliminatedMove <= '1;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_renameTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_dispatchTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_enqRsTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_selectTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_issueTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_writebackTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_runahead_checkpoint_id <= '1;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_tlbFirstReqTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_tlbRespTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debug_seqNum <= '1;
        vif.drv_mp.drv_cb.io_writeback_16_valid <= '1;
        vif.drv_mp.drv_cb.io_writeback_16_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_writeback_16_bits_data_1 <= '1;
        vif.drv_mp.drv_cb.io_writeback_16_bits_data_2 <= '1;
        vif.drv_mp.drv_cb.io_writeback_16_bits_data_3 <= '1;
        vif.drv_mp.drv_cb.io_writeback_16_bits_pdest <= '1;
        vif.drv_mp.drv_cb.io_writeback_16_bits_robIdx_flag <= '1;
        vif.drv_mp.drv_cb.io_writeback_16_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_writeback_16_bits_fpWen <= '1;
        vif.drv_mp.drv_cb.io_writeback_16_bits_vecWen <= '1;
        vif.drv_mp.drv_cb.io_writeback_16_bits_v0Wen <= '1;
        vif.drv_mp.drv_cb.io_writeback_16_bits_fflags <= '1;
        vif.drv_mp.drv_cb.io_writeback_16_bits_wflags <= '1;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_eliminatedMove <= '1;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_renameTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_dispatchTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_enqRsTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_selectTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_issueTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_writebackTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_runahead_checkpoint_id <= '1;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_tlbFirstReqTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_tlbRespTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debug_seqNum <= '1;
        vif.drv_mp.drv_cb.io_writeback_15_valid <= '1;
        vif.drv_mp.drv_cb.io_writeback_15_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_writeback_15_bits_data_1 <= '1;
        vif.drv_mp.drv_cb.io_writeback_15_bits_data_2 <= '1;
        vif.drv_mp.drv_cb.io_writeback_15_bits_pdest <= '1;
        vif.drv_mp.drv_cb.io_writeback_15_bits_robIdx_flag <= '1;
        vif.drv_mp.drv_cb.io_writeback_15_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_writeback_15_bits_vecWen <= '1;
        vif.drv_mp.drv_cb.io_writeback_15_bits_v0Wen <= '1;
        vif.drv_mp.drv_cb.io_writeback_15_bits_fflags <= '1;
        vif.drv_mp.drv_cb.io_writeback_15_bits_wflags <= '1;
        vif.drv_mp.drv_cb.io_writeback_15_bits_vxsat <= '1;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_eliminatedMove <= '1;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_renameTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_dispatchTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_enqRsTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_selectTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_issueTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_writebackTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_runahead_checkpoint_id <= '1;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_tlbFirstReqTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_tlbRespTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debug_seqNum <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_valid <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_1 <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_2 <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_3 <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_4 <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_5 <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_bits_pdest <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_bits_robIdx_flag <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_bits_intWen <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_bits_fpWen <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_bits_vecWen <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_bits_v0Wen <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_bits_vlWen <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_bits_fflags <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_bits_wflags <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_bits_exceptionVec_2 <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_eliminatedMove <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_renameTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_dispatchTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_enqRsTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_selectTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_issueTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_writebackTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_runahead_checkpoint_id <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_tlbFirstReqTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_tlbRespTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debug_seqNum <= '1;
        vif.drv_mp.drv_cb.io_writeback_13_valid <= '1;
        vif.drv_mp.drv_cb.io_writeback_13_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_writeback_13_bits_data_1 <= '1;
        vif.drv_mp.drv_cb.io_writeback_13_bits_data_2 <= '1;
        vif.drv_mp.drv_cb.io_writeback_13_bits_pdest <= '1;
        vif.drv_mp.drv_cb.io_writeback_13_bits_robIdx_flag <= '1;
        vif.drv_mp.drv_cb.io_writeback_13_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_writeback_13_bits_vecWen <= '1;
        vif.drv_mp.drv_cb.io_writeback_13_bits_v0Wen <= '1;
        vif.drv_mp.drv_cb.io_writeback_13_bits_fflags <= '1;
        vif.drv_mp.drv_cb.io_writeback_13_bits_wflags <= '1;
        vif.drv_mp.drv_cb.io_writeback_13_bits_vxsat <= '1;
        vif.drv_mp.drv_cb.io_writeback_13_bits_exceptionVec_2 <= '1;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_eliminatedMove <= '1;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_renameTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_dispatchTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_enqRsTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_selectTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_issueTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_writebackTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_runahead_checkpoint_id <= '1;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_tlbFirstReqTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_tlbRespTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debug_seqNum <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_valid <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_data_1 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_pdest <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_robIdx_flag <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_intWen <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_valid <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_isRVC <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_robIdx_flag <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_ftqIdx_flag <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_ftqIdx_value <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_ftqOffset <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_level <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_interrupt <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pc <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_ssp <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_sctr <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_ghr <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_target <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_taken <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_shift <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_fullTarget <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_stFtqIdx_flag <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_stFtqIdx_value <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_stFtqOffset <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_debugIsCtrl <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_debugIsMemVio <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_2 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_3 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_8 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_9 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_10 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_11 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_22 <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_flushPipe <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_valid <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_isRVC <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_brType <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_isCall <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_isRet <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debug_isPerfCnt <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_eliminatedMove <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_renameTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_dispatchTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_enqRsTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_selectTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_issueTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_writebackTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_runahead_checkpoint_id <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_tlbFirstReqTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_tlbRespTime <= '1;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debug_seqNum <= '1;
        vif.drv_mp.drv_cb.io_writeback_5_valid <= '1;
        vif.drv_mp.drv_cb.io_writeback_5_bits_redirect_valid <= '1;
        vif.drv_mp.drv_cb.io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred <= '1;
        vif.drv_mp.drv_cb.io_writeback_3_valid <= '1;
        vif.drv_mp.drv_cb.io_writeback_3_bits_redirect_valid <= '1;
        vif.drv_mp.drv_cb.io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred <= '1;
        vif.drv_mp.drv_cb.io_writeback_1_valid <= '1;
        vif.drv_mp.drv_cb.io_writeback_1_bits_redirect_valid <= '1;
        vif.drv_mp.drv_cb.io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_26_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_26_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_25_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_25_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_24_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_pdest <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_vecWen <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_v0Wen <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_vls_vdIdx <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_debug_isMMIO <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_debug_isNCIO <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_debug_isPerfCnt <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_debug_paddr <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_23_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_pdest <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_vecWen <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_v0Wen <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_vls_vdIdx <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_debug_isMMIO <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_debug_isNCIO <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_debug_isPerfCnt <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_debug_paddr <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_22_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_lqIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_debug_isMMIO <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_debug_isNCIO <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_debug_isPerfCnt <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_debug_paddr <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_21_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_lqIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_debug_isMMIO <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_debug_isNCIO <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_debug_isPerfCnt <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_debug_paddr <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_20_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_lqIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_debug_isMMIO <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_debug_isNCIO <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_debug_isPerfCnt <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_debug_paddr <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_19_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_sqIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_debug_isMMIO <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_debug_isNCIO <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_debug_isPerfCnt <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_debug_paddr <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_18_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_sqIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_debug_isMMIO <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_debug_isNCIO <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_debug_isPerfCnt <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_debug_paddr <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_17_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_17_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_17_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_17_bits_fflags <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_17_bits_wflags <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_16_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_16_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_16_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_16_bits_fflags <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_16_bits_wflags <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_15_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_15_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_15_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_15_bits_fflags <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_15_bits_wflags <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_15_bits_vxsat <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_14_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_14_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_14_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_14_bits_fflags <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_14_bits_wflags <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_13_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_13_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_13_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_13_bits_fflags <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_13_bits_wflags <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_13_bits_vxsat <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_12_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_12_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_12_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_12_bits_fflags <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_12_bits_wflags <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_11_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_11_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_11_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_11_bits_fflags <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_11_bits_wflags <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_10_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_10_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_10_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_10_bits_fflags <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_10_bits_wflags <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_9_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_9_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_9_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_9_bits_fflags <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_9_bits_wflags <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_8_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_8_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_8_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_8_bits_fflags <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_8_bits_wflags <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_7_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_7_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_7_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_7_bits_debug_isPerfCnt <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_6_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_6_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_6_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_5_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_redirect_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_fflags <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_wflags <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_4_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_4_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_4_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_3_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_3_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_3_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_3_bits_redirect_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_2_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_2_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_2_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_1_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_1_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_1_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_1_bits_redirect_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_0_valid <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_0_bits_data_0 <= '1;
        vif.drv_mp.drv_cb.io_exuWriteback_0_bits_robIdx_value <= '1;
        vif.drv_mp.drv_cb.io_writebackNums_0_bits <= '1;
        vif.drv_mp.drv_cb.io_writebackNums_1_bits <= '1;
        vif.drv_mp.drv_cb.io_writebackNums_2_bits <= '1;
        vif.drv_mp.drv_cb.io_writebackNums_3_bits <= '1;
        vif.drv_mp.drv_cb.io_writebackNums_4_bits <= '1;
        vif.drv_mp.drv_cb.io_writebackNums_5_bits <= '1;
        vif.drv_mp.drv_cb.io_writebackNums_6_bits <= '1;
        vif.drv_mp.drv_cb.io_writebackNums_7_bits <= '1;
        vif.drv_mp.drv_cb.io_writebackNums_8_bits <= '1;
        vif.drv_mp.drv_cb.io_writebackNums_9_bits <= '1;
        vif.drv_mp.drv_cb.io_writebackNums_10_bits <= '1;
        vif.drv_mp.drv_cb.io_writebackNums_11_bits <= '1;
        vif.drv_mp.drv_cb.io_writebackNums_12_bits <= '1;
        vif.drv_mp.drv_cb.io_writebackNums_13_bits <= '1;
        vif.drv_mp.drv_cb.io_writebackNums_14_bits <= '1;
        vif.drv_mp.drv_cb.io_writebackNums_15_bits <= '1;
        vif.drv_mp.drv_cb.io_writebackNums_16_bits <= '1;
        vif.drv_mp.drv_cb.io_writebackNums_17_bits <= '1;
        vif.drv_mp.drv_cb.io_writebackNums_18_bits <= '1;
        vif.drv_mp.drv_cb.io_writebackNums_19_bits <= '1;
        vif.drv_mp.drv_cb.io_writebackNums_20_bits <= '1;
        vif.drv_mp.drv_cb.io_writebackNums_21_bits <= '1;
        vif.drv_mp.drv_cb.io_writebackNums_22_bits <= '1;
        vif.drv_mp.drv_cb.io_writebackNums_23_bits <= '1;
        vif.drv_mp.drv_cb.io_writebackNums_24_bits <= '1;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_0 <= '1;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_1 <= '1;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_2 <= '1;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_6 <= '1;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_7 <= '1;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_8 <= '1;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_9 <= '1;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_10 <= '1;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_11 <= '1;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_12 <= '1;

    end
    else if(drv_mode==tcnt_dec_base::DRV_X) begin
        vif.drv_mp.drv_cb.io_writeback_24_valid <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_pdest <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_robIdx_flag <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vecWen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_v0Wen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vlWen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_0 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_1 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_2 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_3 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_4 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_5 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_6 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_7 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_8 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_9 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_10 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_11 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_12 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_13 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_14 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_15 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_16 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_17 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_18 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_19 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_20 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_21 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_22 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_23 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_flushPipe <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_replay <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_trigger <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vill <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vma <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vta <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vsew <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vlmul <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVill <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVma <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVta <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVsew <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVlmul <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vm <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vstart <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_frm <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFP32Instr <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFP64Instr <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isReduction <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vxrm <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vuopIdx <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_lastUop <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vmask <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vl <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_nf <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_veew <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isReverse <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isExt <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isNarrow <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isDstMask <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isOpMask <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isMove <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isDependOldVd <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isWritePartVd <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isVleff <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_oldVdPsrc <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vdIdx <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vdIdxInField <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isIndexed <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isMasked <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isStrided <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isWhole <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isVecLoad <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isVlm <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_isMMIO <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_isNCIO <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_isPerfCnt <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_paddr <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_vaddr <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_eliminatedMove <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_renameTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_dispatchTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_enqRsTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_selectTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_issueTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_writebackTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_runahead_checkpoint_id <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_tlbFirstReqTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_tlbRespTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_seqNum <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_valid <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_pdest <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_robIdx_flag <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vecWen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_v0Wen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vlWen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_0 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_1 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_2 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_3 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_4 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_5 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_6 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_7 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_8 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_9 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_10 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_11 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_12 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_13 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_14 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_15 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_16 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_17 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_18 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_19 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_20 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_21 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_22 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_23 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_flushPipe <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_replay <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_trigger <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vill <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vma <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vta <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vsew <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vlmul <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVill <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVma <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVta <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVsew <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVlmul <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vm <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vstart <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_frm <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFP32Instr <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFP64Instr <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isReduction <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vxrm <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vuopIdx <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_lastUop <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vmask <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vl <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_nf <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_veew <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isReverse <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isExt <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isNarrow <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isDstMask <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isOpMask <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isMove <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isDependOldVd <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isWritePartVd <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isVleff <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_oldVdPsrc <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vdIdx <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vdIdxInField <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isIndexed <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isMasked <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isStrided <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isWhole <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isVecLoad <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isVlm <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_isMMIO <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_isNCIO <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_isPerfCnt <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_paddr <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_vaddr <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_eliminatedMove <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_renameTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_dispatchTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_enqRsTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_selectTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_issueTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_writebackTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_runahead_checkpoint_id <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_tlbFirstReqTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_tlbRespTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_seqNum <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_valid <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_pdest <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_robIdx_flag <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_intWen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_fpWen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_0 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_1 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_2 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_3 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_4 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_5 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_6 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_7 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_8 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_9 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_10 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_11 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_12 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_13 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_14 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_15 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_16 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_17 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_18 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_19 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_20 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_21 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_22 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_23 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_flushPipe <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_replay <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_lqIdx_flag <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_lqIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_trigger <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_valid <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_isRVC <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_brType <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_isCall <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_isRet <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_isMMIO <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_isNCIO <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_isPerfCnt <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_paddr <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_vaddr <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_eliminatedMove <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_renameTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_dispatchTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_enqRsTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_selectTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_issueTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_writebackTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_runahead_checkpoint_id <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_tlbFirstReqTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_tlbRespTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_seqNum <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_valid <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_pdest <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_robIdx_flag <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_intWen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_fpWen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_0 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_1 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_2 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_3 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_4 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_5 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_6 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_7 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_8 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_9 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_10 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_11 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_12 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_13 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_14 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_15 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_16 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_17 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_18 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_19 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_20 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_21 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_22 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_23 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_flushPipe <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_replay <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_lqIdx_flag <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_lqIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_trigger <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_valid <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_isRVC <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_brType <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_isCall <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_isRet <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_isMMIO <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_isNCIO <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_isPerfCnt <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_paddr <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_vaddr <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_eliminatedMove <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_renameTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_dispatchTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_enqRsTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_selectTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_issueTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_writebackTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_runahead_checkpoint_id <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_tlbFirstReqTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_tlbRespTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_seqNum <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_valid <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_pdest <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_robIdx_flag <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_intWen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_fpWen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_0 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_1 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_2 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_3 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_4 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_5 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_6 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_7 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_8 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_9 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_10 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_11 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_12 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_13 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_14 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_15 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_16 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_17 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_18 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_19 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_20 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_21 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_22 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_23 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_flushPipe <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_replay <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_lqIdx_flag <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_lqIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_trigger <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_valid <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_isRVC <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_brType <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_isCall <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_isRet <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_isMMIO <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_isNCIO <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_isPerfCnt <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_paddr <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_vaddr <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_eliminatedMove <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_renameTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_dispatchTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_enqRsTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_selectTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_issueTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_writebackTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_runahead_checkpoint_id <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_tlbFirstReqTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_tlbRespTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_seqNum <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_valid <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_pdest <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_robIdx_flag <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_intWen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_0 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_1 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_2 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_3 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_4 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_5 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_6 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_7 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_8 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_9 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_10 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_11 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_12 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_13 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_14 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_15 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_16 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_17 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_18 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_19 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_20 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_21 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_22 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_23 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_flushPipe <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_sqIdx_flag <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_sqIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_trigger <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_isMMIO <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_isNCIO <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_isPerfCnt <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_paddr <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_vaddr <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_eliminatedMove <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_renameTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_dispatchTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_enqRsTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_selectTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_issueTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_writebackTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_runahead_checkpoint_id <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_tlbFirstReqTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_tlbRespTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_seqNum <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_valid <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_pdest <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_robIdx_flag <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_intWen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_0 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_1 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_2 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_3 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_4 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_5 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_6 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_7 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_8 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_9 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_10 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_11 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_12 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_13 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_14 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_15 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_16 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_17 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_18 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_19 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_20 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_21 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_22 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_23 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_flushPipe <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_sqIdx_flag <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_sqIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_trigger <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_isMMIO <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_isNCIO <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_isPerfCnt <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_paddr <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_vaddr <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_eliminatedMove <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_renameTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_dispatchTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_enqRsTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_selectTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_issueTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_writebackTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_runahead_checkpoint_id <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_tlbFirstReqTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_tlbRespTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_seqNum <= 'x;
        vif.drv_mp.drv_cb.io_writeback_17_valid <= 'x;
        vif.drv_mp.drv_cb.io_writeback_17_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_17_bits_data_1 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_17_bits_data_2 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_17_bits_pdest <= 'x;
        vif.drv_mp.drv_cb.io_writeback_17_bits_robIdx_flag <= 'x;
        vif.drv_mp.drv_cb.io_writeback_17_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_writeback_17_bits_vecWen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_17_bits_v0Wen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_17_bits_fflags <= 'x;
        vif.drv_mp.drv_cb.io_writeback_17_bits_wflags <= 'x;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_eliminatedMove <= 'x;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_renameTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_dispatchTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_enqRsTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_selectTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_issueTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_writebackTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_runahead_checkpoint_id <= 'x;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_tlbFirstReqTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_tlbRespTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debug_seqNum <= 'x;
        vif.drv_mp.drv_cb.io_writeback_16_valid <= 'x;
        vif.drv_mp.drv_cb.io_writeback_16_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_16_bits_data_1 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_16_bits_data_2 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_16_bits_data_3 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_16_bits_pdest <= 'x;
        vif.drv_mp.drv_cb.io_writeback_16_bits_robIdx_flag <= 'x;
        vif.drv_mp.drv_cb.io_writeback_16_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_writeback_16_bits_fpWen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_16_bits_vecWen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_16_bits_v0Wen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_16_bits_fflags <= 'x;
        vif.drv_mp.drv_cb.io_writeback_16_bits_wflags <= 'x;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_eliminatedMove <= 'x;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_renameTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_dispatchTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_enqRsTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_selectTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_issueTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_writebackTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_runahead_checkpoint_id <= 'x;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_tlbFirstReqTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_tlbRespTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debug_seqNum <= 'x;
        vif.drv_mp.drv_cb.io_writeback_15_valid <= 'x;
        vif.drv_mp.drv_cb.io_writeback_15_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_15_bits_data_1 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_15_bits_data_2 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_15_bits_pdest <= 'x;
        vif.drv_mp.drv_cb.io_writeback_15_bits_robIdx_flag <= 'x;
        vif.drv_mp.drv_cb.io_writeback_15_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_writeback_15_bits_vecWen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_15_bits_v0Wen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_15_bits_fflags <= 'x;
        vif.drv_mp.drv_cb.io_writeback_15_bits_wflags <= 'x;
        vif.drv_mp.drv_cb.io_writeback_15_bits_vxsat <= 'x;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_eliminatedMove <= 'x;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_renameTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_dispatchTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_enqRsTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_selectTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_issueTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_writebackTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_runahead_checkpoint_id <= 'x;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_tlbFirstReqTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_tlbRespTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debug_seqNum <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_valid <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_1 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_2 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_3 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_4 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_5 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_bits_pdest <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_bits_robIdx_flag <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_bits_intWen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_bits_fpWen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_bits_vecWen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_bits_v0Wen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_bits_vlWen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_bits_fflags <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_bits_wflags <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_bits_exceptionVec_2 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_eliminatedMove <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_renameTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_dispatchTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_enqRsTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_selectTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_issueTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_writebackTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_runahead_checkpoint_id <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_tlbFirstReqTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_tlbRespTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debug_seqNum <= 'x;
        vif.drv_mp.drv_cb.io_writeback_13_valid <= 'x;
        vif.drv_mp.drv_cb.io_writeback_13_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_13_bits_data_1 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_13_bits_data_2 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_13_bits_pdest <= 'x;
        vif.drv_mp.drv_cb.io_writeback_13_bits_robIdx_flag <= 'x;
        vif.drv_mp.drv_cb.io_writeback_13_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_writeback_13_bits_vecWen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_13_bits_v0Wen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_13_bits_fflags <= 'x;
        vif.drv_mp.drv_cb.io_writeback_13_bits_wflags <= 'x;
        vif.drv_mp.drv_cb.io_writeback_13_bits_vxsat <= 'x;
        vif.drv_mp.drv_cb.io_writeback_13_bits_exceptionVec_2 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_eliminatedMove <= 'x;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_renameTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_dispatchTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_enqRsTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_selectTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_issueTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_writebackTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_runahead_checkpoint_id <= 'x;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_tlbFirstReqTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_tlbRespTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debug_seqNum <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_valid <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_data_1 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_pdest <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_robIdx_flag <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_intWen <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_valid <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_isRVC <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_robIdx_flag <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_ftqIdx_flag <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_ftqIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_ftqOffset <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_level <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_interrupt <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pc <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_ssp <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_sctr <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_ghr <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_target <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_taken <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_shift <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_fullTarget <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_stFtqIdx_flag <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_stFtqIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_stFtqOffset <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_debugIsCtrl <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_debugIsMemVio <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_2 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_3 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_8 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_9 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_10 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_11 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_22 <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_flushPipe <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_valid <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_isRVC <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_brType <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_isCall <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_isRet <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debug_isPerfCnt <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_eliminatedMove <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_renameTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_dispatchTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_enqRsTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_selectTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_issueTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_writebackTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_runahead_checkpoint_id <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_tlbFirstReqTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_tlbRespTime <= 'x;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debug_seqNum <= 'x;
        vif.drv_mp.drv_cb.io_writeback_5_valid <= 'x;
        vif.drv_mp.drv_cb.io_writeback_5_bits_redirect_valid <= 'x;
        vif.drv_mp.drv_cb.io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred <= 'x;
        vif.drv_mp.drv_cb.io_writeback_3_valid <= 'x;
        vif.drv_mp.drv_cb.io_writeback_3_bits_redirect_valid <= 'x;
        vif.drv_mp.drv_cb.io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred <= 'x;
        vif.drv_mp.drv_cb.io_writeback_1_valid <= 'x;
        vif.drv_mp.drv_cb.io_writeback_1_bits_redirect_valid <= 'x;
        vif.drv_mp.drv_cb.io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_26_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_26_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_25_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_25_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_24_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_pdest <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_vecWen <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_v0Wen <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_vls_vdIdx <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_debug_isMMIO <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_debug_isNCIO <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_debug_isPerfCnt <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_debug_paddr <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_23_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_pdest <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_vecWen <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_v0Wen <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_vls_vdIdx <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_debug_isMMIO <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_debug_isNCIO <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_debug_isPerfCnt <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_debug_paddr <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_22_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_lqIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_debug_isMMIO <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_debug_isNCIO <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_debug_isPerfCnt <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_debug_paddr <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_21_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_lqIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_debug_isMMIO <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_debug_isNCIO <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_debug_isPerfCnt <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_debug_paddr <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_20_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_lqIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_debug_isMMIO <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_debug_isNCIO <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_debug_isPerfCnt <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_debug_paddr <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_19_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_sqIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_debug_isMMIO <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_debug_isNCIO <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_debug_isPerfCnt <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_debug_paddr <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_18_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_sqIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_debug_isMMIO <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_debug_isNCIO <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_debug_isPerfCnt <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_debug_paddr <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_17_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_17_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_17_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_17_bits_fflags <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_17_bits_wflags <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_16_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_16_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_16_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_16_bits_fflags <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_16_bits_wflags <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_15_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_15_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_15_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_15_bits_fflags <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_15_bits_wflags <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_15_bits_vxsat <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_14_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_14_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_14_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_14_bits_fflags <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_14_bits_wflags <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_13_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_13_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_13_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_13_bits_fflags <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_13_bits_wflags <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_13_bits_vxsat <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_12_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_12_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_12_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_12_bits_fflags <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_12_bits_wflags <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_11_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_11_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_11_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_11_bits_fflags <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_11_bits_wflags <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_10_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_10_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_10_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_10_bits_fflags <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_10_bits_wflags <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_9_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_9_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_9_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_9_bits_fflags <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_9_bits_wflags <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_8_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_8_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_8_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_8_bits_fflags <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_8_bits_wflags <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_7_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_7_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_7_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_7_bits_debug_isPerfCnt <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_6_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_6_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_6_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_5_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_redirect_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_fflags <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_wflags <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_4_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_4_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_4_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_3_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_3_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_3_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_3_bits_redirect_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_2_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_2_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_2_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_1_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_1_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_1_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_1_bits_redirect_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_0_valid <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_0_bits_data_0 <= 'x;
        vif.drv_mp.drv_cb.io_exuWriteback_0_bits_robIdx_value <= 'x;
        vif.drv_mp.drv_cb.io_writebackNums_0_bits <= 'x;
        vif.drv_mp.drv_cb.io_writebackNums_1_bits <= 'x;
        vif.drv_mp.drv_cb.io_writebackNums_2_bits <= 'x;
        vif.drv_mp.drv_cb.io_writebackNums_3_bits <= 'x;
        vif.drv_mp.drv_cb.io_writebackNums_4_bits <= 'x;
        vif.drv_mp.drv_cb.io_writebackNums_5_bits <= 'x;
        vif.drv_mp.drv_cb.io_writebackNums_6_bits <= 'x;
        vif.drv_mp.drv_cb.io_writebackNums_7_bits <= 'x;
        vif.drv_mp.drv_cb.io_writebackNums_8_bits <= 'x;
        vif.drv_mp.drv_cb.io_writebackNums_9_bits <= 'x;
        vif.drv_mp.drv_cb.io_writebackNums_10_bits <= 'x;
        vif.drv_mp.drv_cb.io_writebackNums_11_bits <= 'x;
        vif.drv_mp.drv_cb.io_writebackNums_12_bits <= 'x;
        vif.drv_mp.drv_cb.io_writebackNums_13_bits <= 'x;
        vif.drv_mp.drv_cb.io_writebackNums_14_bits <= 'x;
        vif.drv_mp.drv_cb.io_writebackNums_15_bits <= 'x;
        vif.drv_mp.drv_cb.io_writebackNums_16_bits <= 'x;
        vif.drv_mp.drv_cb.io_writebackNums_17_bits <= 'x;
        vif.drv_mp.drv_cb.io_writebackNums_18_bits <= 'x;
        vif.drv_mp.drv_cb.io_writebackNums_19_bits <= 'x;
        vif.drv_mp.drv_cb.io_writebackNums_20_bits <= 'x;
        vif.drv_mp.drv_cb.io_writebackNums_21_bits <= 'x;
        vif.drv_mp.drv_cb.io_writebackNums_22_bits <= 'x;
        vif.drv_mp.drv_cb.io_writebackNums_23_bits <= 'x;
        vif.drv_mp.drv_cb.io_writebackNums_24_bits <= 'x;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_0 <= 'x;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_1 <= 'x;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_2 <= 'x;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_6 <= 'x;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_7 <= 'x;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_8 <= 'x;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_9 <= 'x;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_10 <= 'x;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_11 <= 'x;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_12 <= 'x;

    end
    else if(drv_mode==tcnt_dec_base::DRV_RAND) begin
        vif.drv_mp.drv_cb.io_writeback_24_valid <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_pdest <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_robIdx_flag <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vecWen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_v0Wen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vlWen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_0 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_1 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_2 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_3 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_4 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_5 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_6 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_7 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_8 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_9 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_10 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_11 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_12 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_13 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_14 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_15 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_16 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_17 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_18 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_19 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_20 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_21 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_22 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_23 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_flushPipe <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_replay <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_trigger <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vill <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vma <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vta <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vsew <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vlmul <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVill <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVma <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVta <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVsew <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVlmul <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vm <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vstart <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_frm <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFP32Instr <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFP64Instr <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isReduction <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vxrm <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vuopIdx <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_lastUop <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vmask <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vl <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_nf <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_veew <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isReverse <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isExt <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isNarrow <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isDstMask <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isOpMask <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isMove <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isDependOldVd <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isWritePartVd <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isVleff <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_oldVdPsrc <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vdIdx <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vdIdxInField <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isIndexed <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isMasked <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isStrided <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isWhole <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isVecLoad <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isVlm <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_isMMIO <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_isNCIO <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_isPerfCnt <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_paddr <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_vaddr <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_eliminatedMove <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_renameTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_dispatchTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_enqRsTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_selectTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_issueTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_writebackTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_runahead_checkpoint_id <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_tlbFirstReqTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_tlbRespTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_seqNum <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_valid <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_pdest <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_robIdx_flag <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vecWen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_v0Wen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vlWen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_0 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_1 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_2 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_3 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_4 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_5 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_6 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_7 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_8 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_9 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_10 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_11 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_12 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_13 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_14 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_15 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_16 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_17 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_18 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_19 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_20 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_21 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_22 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_23 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_flushPipe <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_replay <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_trigger <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vill <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vma <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vta <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vsew <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vlmul <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVill <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVma <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVta <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVsew <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVlmul <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vm <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vstart <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_frm <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFP32Instr <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFP64Instr <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isReduction <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vxrm <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vuopIdx <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_lastUop <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vmask <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vl <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_nf <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_veew <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isReverse <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isExt <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isNarrow <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isDstMask <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isOpMask <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isMove <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isDependOldVd <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isWritePartVd <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isVleff <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_oldVdPsrc <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vdIdx <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vdIdxInField <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isIndexed <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isMasked <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isStrided <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isWhole <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isVecLoad <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isVlm <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_isMMIO <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_isNCIO <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_isPerfCnt <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_paddr <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_vaddr <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_eliminatedMove <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_renameTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_dispatchTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_enqRsTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_selectTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_issueTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_writebackTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_runahead_checkpoint_id <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_tlbFirstReqTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_tlbRespTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_seqNum <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_valid <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_pdest <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_robIdx_flag <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_intWen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_fpWen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_0 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_1 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_2 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_3 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_4 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_5 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_6 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_7 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_8 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_9 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_10 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_11 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_12 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_13 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_14 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_15 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_16 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_17 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_18 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_19 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_20 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_21 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_22 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_23 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_flushPipe <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_replay <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_lqIdx_flag <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_lqIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_trigger <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_valid <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_isRVC <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_brType <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_isCall <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_isRet <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_isMMIO <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_isNCIO <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_isPerfCnt <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_paddr <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_vaddr <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_eliminatedMove <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_renameTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_dispatchTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_enqRsTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_selectTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_issueTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_writebackTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_runahead_checkpoint_id <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_tlbFirstReqTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_tlbRespTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_seqNum <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_valid <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_pdest <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_robIdx_flag <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_intWen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_fpWen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_0 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_1 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_2 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_3 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_4 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_5 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_6 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_7 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_8 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_9 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_10 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_11 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_12 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_13 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_14 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_15 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_16 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_17 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_18 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_19 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_20 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_21 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_22 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_23 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_flushPipe <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_replay <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_lqIdx_flag <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_lqIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_trigger <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_valid <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_isRVC <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_brType <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_isCall <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_isRet <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_isMMIO <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_isNCIO <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_isPerfCnt <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_paddr <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_vaddr <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_eliminatedMove <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_renameTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_dispatchTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_enqRsTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_selectTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_issueTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_writebackTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_runahead_checkpoint_id <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_tlbFirstReqTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_tlbRespTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_seqNum <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_valid <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_pdest <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_robIdx_flag <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_intWen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_fpWen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_0 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_1 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_2 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_3 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_4 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_5 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_6 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_7 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_8 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_9 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_10 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_11 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_12 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_13 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_14 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_15 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_16 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_17 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_18 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_19 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_20 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_21 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_22 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_23 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_flushPipe <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_replay <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_lqIdx_flag <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_lqIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_trigger <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_valid <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_isRVC <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_brType <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_isCall <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_isRet <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_isMMIO <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_isNCIO <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_isPerfCnt <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_paddr <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_vaddr <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_eliminatedMove <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_renameTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_dispatchTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_enqRsTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_selectTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_issueTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_writebackTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_runahead_checkpoint_id <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_tlbFirstReqTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_tlbRespTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_seqNum <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_valid <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_pdest <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_robIdx_flag <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_intWen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_0 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_1 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_2 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_3 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_4 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_5 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_6 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_7 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_8 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_9 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_10 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_11 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_12 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_13 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_14 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_15 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_16 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_17 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_18 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_19 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_20 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_21 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_22 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_23 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_flushPipe <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_sqIdx_flag <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_sqIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_trigger <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_isMMIO <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_isNCIO <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_isPerfCnt <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_paddr <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_vaddr <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_eliminatedMove <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_renameTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_dispatchTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_enqRsTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_selectTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_issueTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_writebackTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_runahead_checkpoint_id <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_tlbFirstReqTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_tlbRespTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_seqNum <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_valid <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_pdest <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_robIdx_flag <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_intWen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_0 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_1 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_2 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_3 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_4 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_5 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_6 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_7 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_8 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_9 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_10 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_11 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_12 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_13 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_14 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_15 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_16 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_17 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_18 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_19 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_20 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_21 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_22 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_23 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_flushPipe <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_sqIdx_flag <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_sqIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_trigger <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_isMMIO <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_isNCIO <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_isPerfCnt <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_paddr <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_vaddr <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_eliminatedMove <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_renameTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_dispatchTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_enqRsTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_selectTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_issueTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_writebackTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_runahead_checkpoint_id <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_tlbFirstReqTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_tlbRespTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_seqNum <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_17_valid <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_17_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_17_bits_data_1 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_17_bits_data_2 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_17_bits_pdest <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_17_bits_robIdx_flag <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_17_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_17_bits_vecWen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_17_bits_v0Wen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_17_bits_fflags <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_17_bits_wflags <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_eliminatedMove <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_renameTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_dispatchTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_enqRsTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_selectTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_issueTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_writebackTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_runahead_checkpoint_id <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_tlbFirstReqTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_tlbRespTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debug_seqNum <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_16_valid <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_16_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_16_bits_data_1 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_16_bits_data_2 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_16_bits_data_3 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_16_bits_pdest <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_16_bits_robIdx_flag <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_16_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_16_bits_fpWen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_16_bits_vecWen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_16_bits_v0Wen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_16_bits_fflags <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_16_bits_wflags <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_eliminatedMove <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_renameTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_dispatchTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_enqRsTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_selectTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_issueTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_writebackTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_runahead_checkpoint_id <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_tlbFirstReqTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_tlbRespTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debug_seqNum <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_15_valid <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_15_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_15_bits_data_1 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_15_bits_data_2 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_15_bits_pdest <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_15_bits_robIdx_flag <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_15_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_15_bits_vecWen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_15_bits_v0Wen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_15_bits_fflags <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_15_bits_wflags <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_15_bits_vxsat <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_eliminatedMove <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_renameTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_dispatchTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_enqRsTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_selectTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_issueTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_writebackTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_runahead_checkpoint_id <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_tlbFirstReqTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_tlbRespTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debug_seqNum <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_valid <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_1 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_2 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_3 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_4 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_5 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_bits_pdest <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_bits_robIdx_flag <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_bits_intWen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_bits_fpWen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_bits_vecWen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_bits_v0Wen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_bits_vlWen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_bits_fflags <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_bits_wflags <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_bits_exceptionVec_2 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_eliminatedMove <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_renameTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_dispatchTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_enqRsTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_selectTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_issueTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_writebackTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_runahead_checkpoint_id <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_tlbFirstReqTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_tlbRespTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debug_seqNum <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_13_valid <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_13_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_13_bits_data_1 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_13_bits_data_2 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_13_bits_pdest <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_13_bits_robIdx_flag <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_13_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_13_bits_vecWen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_13_bits_v0Wen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_13_bits_fflags <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_13_bits_wflags <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_13_bits_vxsat <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_13_bits_exceptionVec_2 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_eliminatedMove <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_renameTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_dispatchTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_enqRsTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_selectTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_issueTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_writebackTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_runahead_checkpoint_id <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_tlbFirstReqTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_tlbRespTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debug_seqNum <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_valid <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_data_1 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_pdest <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_robIdx_flag <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_intWen <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_valid <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_isRVC <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_robIdx_flag <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_ftqIdx_flag <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_ftqIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_ftqOffset <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_level <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_interrupt <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pc <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_ssp <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_sctr <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_ghr <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_target <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_taken <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_shift <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_fullTarget <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_stFtqIdx_flag <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_stFtqIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_stFtqOffset <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_debugIsCtrl <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_debugIsMemVio <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_2 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_3 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_8 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_9 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_10 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_11 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_22 <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_flushPipe <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_valid <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_isRVC <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_brType <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_isCall <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_isRet <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debug_isPerfCnt <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_eliminatedMove <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_renameTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_dispatchTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_enqRsTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_selectTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_issueTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_writebackTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_runahead_checkpoint_id <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_tlbFirstReqTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_tlbRespTime <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debug_seqNum <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_5_valid <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_5_bits_redirect_valid <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_3_valid <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_3_bits_redirect_valid <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_1_valid <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_1_bits_redirect_valid <= $urandom;
        vif.drv_mp.drv_cb.io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_26_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_26_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_25_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_25_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_24_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_pdest <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_vecWen <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_v0Wen <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_vls_vdIdx <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_debug_isMMIO <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_debug_isNCIO <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_debug_isPerfCnt <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_debug_paddr <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_23_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_pdest <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_vecWen <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_v0Wen <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_vls_vdIdx <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_debug_isMMIO <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_debug_isNCIO <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_debug_isPerfCnt <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_debug_paddr <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_22_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_lqIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_debug_isMMIO <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_debug_isNCIO <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_debug_isPerfCnt <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_debug_paddr <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_21_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_lqIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_debug_isMMIO <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_debug_isNCIO <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_debug_isPerfCnt <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_debug_paddr <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_20_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_lqIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_debug_isMMIO <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_debug_isNCIO <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_debug_isPerfCnt <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_debug_paddr <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_19_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_sqIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_debug_isMMIO <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_debug_isNCIO <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_debug_isPerfCnt <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_debug_paddr <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_18_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_sqIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_debug_isMMIO <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_debug_isNCIO <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_debug_isPerfCnt <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_debug_paddr <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_17_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_17_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_17_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_17_bits_fflags <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_17_bits_wflags <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_16_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_16_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_16_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_16_bits_fflags <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_16_bits_wflags <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_15_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_15_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_15_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_15_bits_fflags <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_15_bits_wflags <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_15_bits_vxsat <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_14_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_14_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_14_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_14_bits_fflags <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_14_bits_wflags <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_13_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_13_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_13_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_13_bits_fflags <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_13_bits_wflags <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_13_bits_vxsat <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_12_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_12_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_12_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_12_bits_fflags <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_12_bits_wflags <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_11_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_11_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_11_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_11_bits_fflags <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_11_bits_wflags <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_10_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_10_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_10_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_10_bits_fflags <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_10_bits_wflags <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_9_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_9_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_9_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_9_bits_fflags <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_9_bits_wflags <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_8_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_8_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_8_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_8_bits_fflags <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_8_bits_wflags <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_7_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_7_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_7_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_7_bits_debug_isPerfCnt <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_6_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_6_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_6_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_5_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_redirect_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_fflags <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_wflags <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_4_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_4_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_4_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_3_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_3_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_3_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_3_bits_redirect_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_2_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_2_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_2_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_1_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_1_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_1_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_1_bits_redirect_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_0_valid <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_0_bits_data_0 <= $urandom;
        vif.drv_mp.drv_cb.io_exuWriteback_0_bits_robIdx_value <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNums_0_bits <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNums_1_bits <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNums_2_bits <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNums_3_bits <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNums_4_bits <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNums_5_bits <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNums_6_bits <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNums_7_bits <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNums_8_bits <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNums_9_bits <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNums_10_bits <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNums_11_bits <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNums_12_bits <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNums_13_bits <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNums_14_bits <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNums_15_bits <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNums_16_bits <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNums_17_bits <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNums_18_bits <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNums_19_bits <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNums_20_bits <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNums_21_bits <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNums_22_bits <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNums_23_bits <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNums_24_bits <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_0 <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_1 <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_2 <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_6 <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_7 <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_8 <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_9 <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_10 <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_11 <= $urandom;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_12 <= $urandom;

    end
    else if(drv_mode==tcnt_dec_base::DRV_LST) begin
        vif.drv_mp.drv_cb.io_writeback_24_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vlWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_4 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_5 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_6 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_7 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_8 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_9 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_10 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_11 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_12 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_13 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_14 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_15 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_16 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_17 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_18 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_19 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_20 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_21 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_22 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_exceptionVec_23 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_flushPipe <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_replay <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_trigger <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vill <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vma <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vta <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vsew <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vlmul <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVill <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVma <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVta <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVsew <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_specVlmul <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vm <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vstart <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_frm <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFP32Instr <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFP64Instr <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isReduction <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8 <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vxrm <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vuopIdx <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_lastUop <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vmask <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_vl <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_nf <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_veew <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isReverse <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isExt <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isNarrow <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isDstMask <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isOpMask <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isDependOldVd <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isWritePartVd <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vpu_isVleff <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_oldVdPsrc <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vdIdx <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_vdIdxInField <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isIndexed <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isMasked <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isStrided <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isWhole <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isVecLoad <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_vls_isVlm <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_isMMIO <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_isNCIO <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_paddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_vaddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_renameTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_dispatchTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_enqRsTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_selectTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_issueTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_writebackTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_runahead_checkpoint_id <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_tlbFirstReqTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debugInfo_tlbRespTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_24_bits_debug_seqNum <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vlWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_4 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_5 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_6 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_7 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_8 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_9 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_10 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_11 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_12 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_13 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_14 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_15 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_16 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_17 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_18 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_19 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_20 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_21 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_22 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_exceptionVec_23 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_flushPipe <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_replay <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_trigger <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vill <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vma <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vta <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vsew <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vlmul <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVill <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVma <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVta <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVsew <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_specVlmul <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vm <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vstart <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_frm <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFP32Instr <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFP64Instr <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isReduction <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8 <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vxrm <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vuopIdx <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_lastUop <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vmask <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_vl <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_nf <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_veew <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isReverse <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isExt <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isNarrow <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isDstMask <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isOpMask <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isDependOldVd <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isWritePartVd <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vpu_isVleff <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_oldVdPsrc <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vdIdx <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_vdIdxInField <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isIndexed <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isMasked <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isStrided <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isWhole <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isVecLoad <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_vls_isVlm <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_isMMIO <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_isNCIO <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_paddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_vaddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_renameTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_dispatchTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_enqRsTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_selectTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_issueTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_writebackTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_runahead_checkpoint_id <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_tlbFirstReqTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debugInfo_tlbRespTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_23_bits_debug_seqNum <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_intWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_fpWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_4 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_5 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_6 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_7 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_8 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_9 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_10 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_11 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_12 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_13 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_14 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_15 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_16 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_17 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_18 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_19 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_20 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_21 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_22 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_exceptionVec_23 <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_flushPipe <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_replay <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_lqIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_lqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_trigger <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_isRVC <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_brType <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_isCall <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_predecodeInfo_isRet <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_isMMIO <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_isNCIO <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_paddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_vaddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_renameTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_dispatchTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_enqRsTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_selectTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_issueTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_writebackTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_runahead_checkpoint_id <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_tlbFirstReqTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debugInfo_tlbRespTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_22_bits_debug_seqNum <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_intWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_fpWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_4 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_5 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_6 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_7 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_8 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_9 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_10 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_11 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_12 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_13 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_14 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_15 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_16 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_17 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_18 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_19 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_20 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_21 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_22 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_exceptionVec_23 <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_flushPipe <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_replay <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_lqIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_lqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_trigger <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_isRVC <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_brType <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_isCall <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_predecodeInfo_isRet <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_isMMIO <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_isNCIO <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_paddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_vaddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_renameTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_dispatchTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_enqRsTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_selectTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_issueTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_writebackTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_runahead_checkpoint_id <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_tlbFirstReqTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debugInfo_tlbRespTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_21_bits_debug_seqNum <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_intWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_fpWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_4 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_5 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_6 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_7 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_8 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_9 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_10 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_11 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_12 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_13 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_14 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_15 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_16 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_17 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_18 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_19 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_20 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_21 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_22 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_exceptionVec_23 <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_flushPipe <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_replay <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_lqIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_lqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_trigger <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_isRVC <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_brType <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_isCall <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_predecodeInfo_isRet <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_isMMIO <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_isNCIO <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_paddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_vaddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_renameTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_dispatchTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_enqRsTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_selectTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_issueTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_writebackTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_runahead_checkpoint_id <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_tlbFirstReqTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debugInfo_tlbRespTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_20_bits_debug_seqNum <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_intWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_4 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_5 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_6 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_7 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_8 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_9 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_10 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_11 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_12 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_13 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_14 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_15 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_16 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_17 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_18 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_19 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_20 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_21 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_22 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_exceptionVec_23 <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_flushPipe <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_sqIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_sqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_trigger <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_isMMIO <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_isNCIO <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_paddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_vaddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_renameTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_dispatchTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_enqRsTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_selectTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_issueTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_writebackTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_runahead_checkpoint_id <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_tlbFirstReqTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debugInfo_tlbRespTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_19_bits_debug_seqNum <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_intWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_4 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_5 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_6 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_7 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_8 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_9 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_10 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_11 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_12 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_13 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_14 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_15 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_16 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_17 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_18 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_19 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_20 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_21 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_22 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_exceptionVec_23 <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_flushPipe <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_sqIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_sqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_trigger <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_isMMIO <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_isNCIO <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_paddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_vaddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_renameTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_dispatchTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_enqRsTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_selectTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_issueTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_writebackTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_runahead_checkpoint_id <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_tlbFirstReqTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debugInfo_tlbRespTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_18_bits_debug_seqNum <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_data_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_data_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_renameTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_dispatchTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_enqRsTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_selectTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_issueTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_writebackTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_runahead_checkpoint_id <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_tlbFirstReqTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debugInfo_tlbRespTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_17_bits_debug_seqNum <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_data_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_data_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_data_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_fpWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_renameTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_dispatchTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_enqRsTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_selectTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_issueTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_writebackTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_runahead_checkpoint_id <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_tlbFirstReqTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debugInfo_tlbRespTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_16_bits_debug_seqNum <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_data_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_data_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_vxsat <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_renameTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_dispatchTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_enqRsTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_selectTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_issueTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_writebackTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_runahead_checkpoint_id <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_tlbFirstReqTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debugInfo_tlbRespTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_15_bits_debug_seqNum <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_4 <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_data_5 <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_intWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_fpWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_vlWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_renameTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_dispatchTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_enqRsTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_selectTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_issueTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_writebackTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_runahead_checkpoint_id <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_tlbFirstReqTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debugInfo_tlbRespTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_14_bits_debug_seqNum <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_data_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_data_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_vxsat <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_renameTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_dispatchTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_enqRsTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_selectTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_issueTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_writebackTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_runahead_checkpoint_id <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_tlbFirstReqTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debugInfo_tlbRespTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_13_bits_debug_seqNum <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_data_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_intWen <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_isRVC <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_robIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_ftqIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_ftqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_ftqOffset <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_level <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_interrupt <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pc <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_ssp <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_sctr <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_ghr <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_target <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_taken <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_shift <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_fullTarget <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_stFtqIdx_flag <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_stFtqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_stFtqOffset <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_debugIsCtrl <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_redirect_bits_debugIsMemVio <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_2 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_3 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_8 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_9 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_10 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_11 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_exceptionVec_22 <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_flushPipe <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_isRVC <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_brType <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_isCall <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_predecodeInfo_isRet <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_eliminatedMove <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_renameTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_dispatchTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_enqRsTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_selectTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_issueTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_writebackTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_runahead_checkpoint_id <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_tlbFirstReqTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debugInfo_tlbRespTime <= '0;
        vif.drv_mp.drv_cb.io_writeback_7_bits_debug_seqNum <= '0;
        vif.drv_mp.drv_cb.io_writeback_5_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_5_bits_redirect_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred <= '0;
        vif.drv_mp.drv_cb.io_writeback_3_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_3_bits_redirect_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred <= '0;
        vif.drv_mp.drv_cb.io_writeback_1_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_1_bits_redirect_valid <= '0;
        vif.drv_mp.drv_cb.io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_26_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_26_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_25_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_25_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_24_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_vls_vdIdx <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_debug_isMMIO <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_debug_isNCIO <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_24_bits_debug_paddr <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_23_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_pdest <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_vecWen <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_v0Wen <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_vls_vdIdx <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_debug_isMMIO <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_debug_isNCIO <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_23_bits_debug_paddr <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_22_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_lqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_debug_isMMIO <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_debug_isNCIO <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_22_bits_debug_paddr <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_21_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_lqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_debug_isMMIO <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_debug_isNCIO <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_21_bits_debug_paddr <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_20_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_lqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_debug_isMMIO <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_debug_isNCIO <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_20_bits_debug_paddr <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_19_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_sqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_debug_isMMIO <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_debug_isNCIO <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_19_bits_debug_paddr <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_18_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_sqIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_debug_isMMIO <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_debug_isNCIO <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_18_bits_debug_paddr <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_17_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_17_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_17_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_17_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_17_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_16_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_16_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_16_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_16_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_16_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_15_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_15_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_15_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_15_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_15_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_15_bits_vxsat <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_14_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_14_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_14_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_14_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_14_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_13_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_13_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_13_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_13_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_13_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_13_bits_vxsat <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_12_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_12_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_12_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_12_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_12_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_11_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_11_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_11_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_11_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_11_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_10_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_10_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_10_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_10_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_10_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_9_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_9_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_9_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_9_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_9_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_8_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_8_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_8_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_8_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_8_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_7_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_7_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_7_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_7_bits_debug_isPerfCnt <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_6_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_6_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_6_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_5_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_redirect_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_fflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_5_bits_wflags <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_4_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_4_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_4_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_3_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_3_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_3_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_3_bits_redirect_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_2_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_2_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_2_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_1_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_1_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_1_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_1_bits_redirect_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_0_valid <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_0_bits_data_0 <= '0;
        vif.drv_mp.drv_cb.io_exuWriteback_0_bits_robIdx_value <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_0_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_1_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_2_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_3_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_4_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_5_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_6_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_7_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_8_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_9_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_10_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_11_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_12_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_13_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_14_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_15_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_16_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_17_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_18_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_19_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_20_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_21_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_22_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_23_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNums_24_bits <= '0;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_0 <= '0;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_1 <= '0;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_2 <= '0;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_6 <= '0;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_7 <= '0;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_8 <= '0;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_9 <= '0;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_10 <= '0;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_11 <= '0;
        vif.drv_mp.drv_cb.io_writebackNeedFlush_12 <= '0;

    end

endtask:drive_idle

`endif


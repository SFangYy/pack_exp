//=========================================================
//File name    : WriteBack_in_agent_xaction.sv
//Author       : nanyunhao
//Module name  : WriteBack_in_agent_xaction
//Discribution : WriteBack_in_agent_xaction : agent transaction
//Date         : 2026-01-22
//=========================================================
`ifndef WRITEBACK_IN_AGENT_XACTION__SV
`define WRITEBACK_IN_AGENT_XACTION__SV

class WriteBack_in_agent_xaction  extends tcnt_data_base;
    rand bit         io_writeback_24_valid;
    rand bit [127:0] io_writeback_24_bits_data_0;
    rand bit [6:0]   io_writeback_24_bits_pdest;
    rand bit         io_writeback_24_bits_robIdx_flag;
    rand bit [7:0]   io_writeback_24_bits_robIdx_value;
    rand bit         io_writeback_24_bits_vecWen;
    rand bit         io_writeback_24_bits_v0Wen;
    rand bit         io_writeback_24_bits_vlWen;
    rand bit         io_writeback_24_bits_exceptionVec_0;
    rand bit         io_writeback_24_bits_exceptionVec_1;
    rand bit         io_writeback_24_bits_exceptionVec_2;
    rand bit         io_writeback_24_bits_exceptionVec_3;
    rand bit         io_writeback_24_bits_exceptionVec_4;
    rand bit         io_writeback_24_bits_exceptionVec_5;
    rand bit         io_writeback_24_bits_exceptionVec_6;
    rand bit         io_writeback_24_bits_exceptionVec_7;
    rand bit         io_writeback_24_bits_exceptionVec_8;
    rand bit         io_writeback_24_bits_exceptionVec_9;
    rand bit         io_writeback_24_bits_exceptionVec_10;
    rand bit         io_writeback_24_bits_exceptionVec_11;
    rand bit         io_writeback_24_bits_exceptionVec_12;
    rand bit         io_writeback_24_bits_exceptionVec_13;
    rand bit         io_writeback_24_bits_exceptionVec_14;
    rand bit         io_writeback_24_bits_exceptionVec_15;
    rand bit         io_writeback_24_bits_exceptionVec_16;
    rand bit         io_writeback_24_bits_exceptionVec_17;
    rand bit         io_writeback_24_bits_exceptionVec_18;
    rand bit         io_writeback_24_bits_exceptionVec_19;
    rand bit         io_writeback_24_bits_exceptionVec_20;
    rand bit         io_writeback_24_bits_exceptionVec_21;
    rand bit         io_writeback_24_bits_exceptionVec_22;
    rand bit         io_writeback_24_bits_exceptionVec_23;
    rand bit         io_writeback_24_bits_flushPipe;
    rand bit         io_writeback_24_bits_replay;
    rand bit [3:0]   io_writeback_24_bits_trigger;
    rand bit         io_writeback_24_bits_vls_vpu_vill;
    rand bit         io_writeback_24_bits_vls_vpu_vma;
    rand bit         io_writeback_24_bits_vls_vpu_vta;
    rand bit [1:0]   io_writeback_24_bits_vls_vpu_vsew;
    rand bit [2:0]   io_writeback_24_bits_vls_vpu_vlmul;
    rand bit         io_writeback_24_bits_vls_vpu_specVill;
    rand bit         io_writeback_24_bits_vls_vpu_specVma;
    rand bit         io_writeback_24_bits_vls_vpu_specVta;
    rand bit [1:0]   io_writeback_24_bits_vls_vpu_specVsew;
    rand bit [2:0]   io_writeback_24_bits_vls_vpu_specVlmul;
    rand bit         io_writeback_24_bits_vls_vpu_vm;
    rand bit [7:0]   io_writeback_24_bits_vls_vpu_vstart;
    rand bit [2:0]   io_writeback_24_bits_vls_vpu_frm;
    rand bit         io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst;
    rand bit         io_writeback_24_bits_vls_vpu_fpu_isFP32Instr;
    rand bit         io_writeback_24_bits_vls_vpu_fpu_isFP64Instr;
    rand bit         io_writeback_24_bits_vls_vpu_fpu_isReduction;
    rand bit         io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2;
    rand bit         io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4;
    rand bit         io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8;
    rand bit [1:0]   io_writeback_24_bits_vls_vpu_vxrm;
    rand bit [6:0]   io_writeback_24_bits_vls_vpu_vuopIdx;
    rand bit         io_writeback_24_bits_vls_vpu_lastUop;
    rand bit [127:0] io_writeback_24_bits_vls_vpu_vmask;
    rand bit [7:0]   io_writeback_24_bits_vls_vpu_vl;
    rand bit [2:0]   io_writeback_24_bits_vls_vpu_nf;
    rand bit [1:0]   io_writeback_24_bits_vls_vpu_veew;
    rand bit         io_writeback_24_bits_vls_vpu_isReverse;
    rand bit         io_writeback_24_bits_vls_vpu_isExt;
    rand bit         io_writeback_24_bits_vls_vpu_isNarrow;
    rand bit         io_writeback_24_bits_vls_vpu_isDstMask;
    rand bit         io_writeback_24_bits_vls_vpu_isOpMask;
    rand bit         io_writeback_24_bits_vls_vpu_isMove;
    rand bit         io_writeback_24_bits_vls_vpu_isDependOldVd;
    rand bit         io_writeback_24_bits_vls_vpu_isWritePartVd;
    rand bit         io_writeback_24_bits_vls_vpu_isVleff;
    rand bit [7:0]   io_writeback_24_bits_vls_oldVdPsrc;
    rand bit [2:0]   io_writeback_24_bits_vls_vdIdx;
    rand bit [2:0]   io_writeback_24_bits_vls_vdIdxInField;
    rand bit         io_writeback_24_bits_vls_isIndexed;
    rand bit         io_writeback_24_bits_vls_isMasked;
    rand bit         io_writeback_24_bits_vls_isStrided;
    rand bit         io_writeback_24_bits_vls_isWhole;
    rand bit         io_writeback_24_bits_vls_isVecLoad;
    rand bit         io_writeback_24_bits_vls_isVlm;
    rand bit         io_writeback_24_bits_debug_isMMIO;
    rand bit         io_writeback_24_bits_debug_isNCIO;
    rand bit         io_writeback_24_bits_debug_isPerfCnt;
    rand bit [47:0]  io_writeback_24_bits_debug_paddr;
    rand bit [49:0]  io_writeback_24_bits_debug_vaddr;
    rand bit         io_writeback_24_bits_debugInfo_eliminatedMove;
    rand bit [63:0]  io_writeback_24_bits_debugInfo_renameTime;
    rand bit [63:0]  io_writeback_24_bits_debugInfo_dispatchTime;
    rand bit [63:0]  io_writeback_24_bits_debugInfo_enqRsTime;
    rand bit [63:0]  io_writeback_24_bits_debugInfo_selectTime;
    rand bit [63:0]  io_writeback_24_bits_debugInfo_issueTime;
    rand bit [63:0]  io_writeback_24_bits_debugInfo_writebackTime;
    rand bit [63:0]  io_writeback_24_bits_debugInfo_runahead_checkpoint_id;
    rand bit [63:0]  io_writeback_24_bits_debugInfo_tlbFirstReqTime;
    rand bit [63:0]  io_writeback_24_bits_debugInfo_tlbRespTime;
    rand bit [63:0]  io_writeback_24_bits_debug_seqNum;
    rand bit         io_writeback_23_valid;
    rand bit [127:0] io_writeback_23_bits_data_0;
    rand bit [6:0]   io_writeback_23_bits_pdest;
    rand bit         io_writeback_23_bits_robIdx_flag;
    rand bit [7:0]   io_writeback_23_bits_robIdx_value;
    rand bit         io_writeback_23_bits_vecWen;
    rand bit         io_writeback_23_bits_v0Wen;
    rand bit         io_writeback_23_bits_vlWen;
    rand bit         io_writeback_23_bits_exceptionVec_0;
    rand bit         io_writeback_23_bits_exceptionVec_1;
    rand bit         io_writeback_23_bits_exceptionVec_2;
    rand bit         io_writeback_23_bits_exceptionVec_3;
    rand bit         io_writeback_23_bits_exceptionVec_4;
    rand bit         io_writeback_23_bits_exceptionVec_5;
    rand bit         io_writeback_23_bits_exceptionVec_6;
    rand bit         io_writeback_23_bits_exceptionVec_7;
    rand bit         io_writeback_23_bits_exceptionVec_8;
    rand bit         io_writeback_23_bits_exceptionVec_9;
    rand bit         io_writeback_23_bits_exceptionVec_10;
    rand bit         io_writeback_23_bits_exceptionVec_11;
    rand bit         io_writeback_23_bits_exceptionVec_12;
    rand bit         io_writeback_23_bits_exceptionVec_13;
    rand bit         io_writeback_23_bits_exceptionVec_14;
    rand bit         io_writeback_23_bits_exceptionVec_15;
    rand bit         io_writeback_23_bits_exceptionVec_16;
    rand bit         io_writeback_23_bits_exceptionVec_17;
    rand bit         io_writeback_23_bits_exceptionVec_18;
    rand bit         io_writeback_23_bits_exceptionVec_19;
    rand bit         io_writeback_23_bits_exceptionVec_20;
    rand bit         io_writeback_23_bits_exceptionVec_21;
    rand bit         io_writeback_23_bits_exceptionVec_22;
    rand bit         io_writeback_23_bits_exceptionVec_23;
    rand bit         io_writeback_23_bits_flushPipe;
    rand bit         io_writeback_23_bits_replay;
    rand bit [3:0]   io_writeback_23_bits_trigger;
    rand bit         io_writeback_23_bits_vls_vpu_vill;
    rand bit         io_writeback_23_bits_vls_vpu_vma;
    rand bit         io_writeback_23_bits_vls_vpu_vta;
    rand bit [1:0]   io_writeback_23_bits_vls_vpu_vsew;
    rand bit [2:0]   io_writeback_23_bits_vls_vpu_vlmul;
    rand bit         io_writeback_23_bits_vls_vpu_specVill;
    rand bit         io_writeback_23_bits_vls_vpu_specVma;
    rand bit         io_writeback_23_bits_vls_vpu_specVta;
    rand bit [1:0]   io_writeback_23_bits_vls_vpu_specVsew;
    rand bit [2:0]   io_writeback_23_bits_vls_vpu_specVlmul;
    rand bit         io_writeback_23_bits_vls_vpu_vm;
    rand bit [7:0]   io_writeback_23_bits_vls_vpu_vstart;
    rand bit [2:0]   io_writeback_23_bits_vls_vpu_frm;
    rand bit         io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst;
    rand bit         io_writeback_23_bits_vls_vpu_fpu_isFP32Instr;
    rand bit         io_writeback_23_bits_vls_vpu_fpu_isFP64Instr;
    rand bit         io_writeback_23_bits_vls_vpu_fpu_isReduction;
    rand bit         io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2;
    rand bit         io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4;
    rand bit         io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8;
    rand bit [1:0]   io_writeback_23_bits_vls_vpu_vxrm;
    rand bit [6:0]   io_writeback_23_bits_vls_vpu_vuopIdx;
    rand bit         io_writeback_23_bits_vls_vpu_lastUop;
    rand bit [127:0] io_writeback_23_bits_vls_vpu_vmask;
    rand bit [7:0]   io_writeback_23_bits_vls_vpu_vl;
    rand bit [2:0]   io_writeback_23_bits_vls_vpu_nf;
    rand bit [1:0]   io_writeback_23_bits_vls_vpu_veew;
    rand bit         io_writeback_23_bits_vls_vpu_isReverse;
    rand bit         io_writeback_23_bits_vls_vpu_isExt;
    rand bit         io_writeback_23_bits_vls_vpu_isNarrow;
    rand bit         io_writeback_23_bits_vls_vpu_isDstMask;
    rand bit         io_writeback_23_bits_vls_vpu_isOpMask;
    rand bit         io_writeback_23_bits_vls_vpu_isMove;
    rand bit         io_writeback_23_bits_vls_vpu_isDependOldVd;
    rand bit         io_writeback_23_bits_vls_vpu_isWritePartVd;
    rand bit         io_writeback_23_bits_vls_vpu_isVleff;
    rand bit [7:0]   io_writeback_23_bits_vls_oldVdPsrc;
    rand bit [2:0]   io_writeback_23_bits_vls_vdIdx;
    rand bit [2:0]   io_writeback_23_bits_vls_vdIdxInField;
    rand bit         io_writeback_23_bits_vls_isIndexed;
    rand bit         io_writeback_23_bits_vls_isMasked;
    rand bit         io_writeback_23_bits_vls_isStrided;
    rand bit         io_writeback_23_bits_vls_isWhole;
    rand bit         io_writeback_23_bits_vls_isVecLoad;
    rand bit         io_writeback_23_bits_vls_isVlm;
    rand bit         io_writeback_23_bits_debug_isMMIO;
    rand bit         io_writeback_23_bits_debug_isNCIO;
    rand bit         io_writeback_23_bits_debug_isPerfCnt;
    rand bit [47:0]  io_writeback_23_bits_debug_paddr;
    rand bit [49:0]  io_writeback_23_bits_debug_vaddr;
    rand bit         io_writeback_23_bits_debugInfo_eliminatedMove;
    rand bit [63:0]  io_writeback_23_bits_debugInfo_renameTime;
    rand bit [63:0]  io_writeback_23_bits_debugInfo_dispatchTime;
    rand bit [63:0]  io_writeback_23_bits_debugInfo_enqRsTime;
    rand bit [63:0]  io_writeback_23_bits_debugInfo_selectTime;
    rand bit [63:0]  io_writeback_23_bits_debugInfo_issueTime;
    rand bit [63:0]  io_writeback_23_bits_debugInfo_writebackTime;
    rand bit [63:0]  io_writeback_23_bits_debugInfo_runahead_checkpoint_id;
    rand bit [63:0]  io_writeback_23_bits_debugInfo_tlbFirstReqTime;
    rand bit [63:0]  io_writeback_23_bits_debugInfo_tlbRespTime;
    rand bit [63:0]  io_writeback_23_bits_debug_seqNum;
    rand bit         io_writeback_22_valid;
    rand bit [63:0]  io_writeback_22_bits_data_0;
    rand bit [7:0]   io_writeback_22_bits_pdest;
    rand bit         io_writeback_22_bits_robIdx_flag;
    rand bit [7:0]   io_writeback_22_bits_robIdx_value;
    rand bit         io_writeback_22_bits_intWen;
    rand bit         io_writeback_22_bits_fpWen;
    rand bit         io_writeback_22_bits_exceptionVec_0;
    rand bit         io_writeback_22_bits_exceptionVec_1;
    rand bit         io_writeback_22_bits_exceptionVec_2;
    rand bit         io_writeback_22_bits_exceptionVec_3;
    rand bit         io_writeback_22_bits_exceptionVec_4;
    rand bit         io_writeback_22_bits_exceptionVec_5;
    rand bit         io_writeback_22_bits_exceptionVec_6;
    rand bit         io_writeback_22_bits_exceptionVec_7;
    rand bit         io_writeback_22_bits_exceptionVec_8;
    rand bit         io_writeback_22_bits_exceptionVec_9;
    rand bit         io_writeback_22_bits_exceptionVec_10;
    rand bit         io_writeback_22_bits_exceptionVec_11;
    rand bit         io_writeback_22_bits_exceptionVec_12;
    rand bit         io_writeback_22_bits_exceptionVec_13;
    rand bit         io_writeback_22_bits_exceptionVec_14;
    rand bit         io_writeback_22_bits_exceptionVec_15;
    rand bit         io_writeback_22_bits_exceptionVec_16;
    rand bit         io_writeback_22_bits_exceptionVec_17;
    rand bit         io_writeback_22_bits_exceptionVec_18;
    rand bit         io_writeback_22_bits_exceptionVec_19;
    rand bit         io_writeback_22_bits_exceptionVec_20;
    rand bit         io_writeback_22_bits_exceptionVec_21;
    rand bit         io_writeback_22_bits_exceptionVec_22;
    rand bit         io_writeback_22_bits_exceptionVec_23;
    rand bit         io_writeback_22_bits_flushPipe;
    rand bit         io_writeback_22_bits_replay;
    rand bit         io_writeback_22_bits_lqIdx_flag;
    rand bit [6:0]   io_writeback_22_bits_lqIdx_value;
    rand bit [3:0]   io_writeback_22_bits_trigger;
    rand bit         io_writeback_22_bits_predecodeInfo_valid;
    rand bit         io_writeback_22_bits_predecodeInfo_isRVC;
    rand bit [1:0]   io_writeback_22_bits_predecodeInfo_brType;
    rand bit         io_writeback_22_bits_predecodeInfo_isCall;
    rand bit         io_writeback_22_bits_predecodeInfo_isRet;
    rand bit         io_writeback_22_bits_debug_isMMIO;
    rand bit         io_writeback_22_bits_debug_isNCIO;
    rand bit         io_writeback_22_bits_debug_isPerfCnt;
    rand bit [47:0]  io_writeback_22_bits_debug_paddr;
    rand bit [49:0]  io_writeback_22_bits_debug_vaddr;
    rand bit         io_writeback_22_bits_debugInfo_eliminatedMove;
    rand bit [63:0]  io_writeback_22_bits_debugInfo_renameTime;
    rand bit [63:0]  io_writeback_22_bits_debugInfo_dispatchTime;
    rand bit [63:0]  io_writeback_22_bits_debugInfo_enqRsTime;
    rand bit [63:0]  io_writeback_22_bits_debugInfo_selectTime;
    rand bit [63:0]  io_writeback_22_bits_debugInfo_issueTime;
    rand bit [63:0]  io_writeback_22_bits_debugInfo_writebackTime;
    rand bit [63:0]  io_writeback_22_bits_debugInfo_runahead_checkpoint_id;
    rand bit [63:0]  io_writeback_22_bits_debugInfo_tlbFirstReqTime;
    rand bit [63:0]  io_writeback_22_bits_debugInfo_tlbRespTime;
    rand bit [63:0]  io_writeback_22_bits_debug_seqNum;
    rand bit         io_writeback_21_valid;
    rand bit [63:0]  io_writeback_21_bits_data_0;
    rand bit [7:0]   io_writeback_21_bits_pdest;
    rand bit         io_writeback_21_bits_robIdx_flag;
    rand bit [7:0]   io_writeback_21_bits_robIdx_value;
    rand bit         io_writeback_21_bits_intWen;
    rand bit         io_writeback_21_bits_fpWen;
    rand bit         io_writeback_21_bits_exceptionVec_0;
    rand bit         io_writeback_21_bits_exceptionVec_1;
    rand bit         io_writeback_21_bits_exceptionVec_2;
    rand bit         io_writeback_21_bits_exceptionVec_3;
    rand bit         io_writeback_21_bits_exceptionVec_4;
    rand bit         io_writeback_21_bits_exceptionVec_5;
    rand bit         io_writeback_21_bits_exceptionVec_6;
    rand bit         io_writeback_21_bits_exceptionVec_7;
    rand bit         io_writeback_21_bits_exceptionVec_8;
    rand bit         io_writeback_21_bits_exceptionVec_9;
    rand bit         io_writeback_21_bits_exceptionVec_10;
    rand bit         io_writeback_21_bits_exceptionVec_11;
    rand bit         io_writeback_21_bits_exceptionVec_12;
    rand bit         io_writeback_21_bits_exceptionVec_13;
    rand bit         io_writeback_21_bits_exceptionVec_14;
    rand bit         io_writeback_21_bits_exceptionVec_15;
    rand bit         io_writeback_21_bits_exceptionVec_16;
    rand bit         io_writeback_21_bits_exceptionVec_17;
    rand bit         io_writeback_21_bits_exceptionVec_18;
    rand bit         io_writeback_21_bits_exceptionVec_19;
    rand bit         io_writeback_21_bits_exceptionVec_20;
    rand bit         io_writeback_21_bits_exceptionVec_21;
    rand bit         io_writeback_21_bits_exceptionVec_22;
    rand bit         io_writeback_21_bits_exceptionVec_23;
    rand bit         io_writeback_21_bits_flushPipe;
    rand bit         io_writeback_21_bits_replay;
    rand bit         io_writeback_21_bits_lqIdx_flag;
    rand bit [6:0]   io_writeback_21_bits_lqIdx_value;
    rand bit [3:0]   io_writeback_21_bits_trigger;
    rand bit         io_writeback_21_bits_predecodeInfo_valid;
    rand bit         io_writeback_21_bits_predecodeInfo_isRVC;
    rand bit [1:0]   io_writeback_21_bits_predecodeInfo_brType;
    rand bit         io_writeback_21_bits_predecodeInfo_isCall;
    rand bit         io_writeback_21_bits_predecodeInfo_isRet;
    rand bit         io_writeback_21_bits_debug_isMMIO;
    rand bit         io_writeback_21_bits_debug_isNCIO;
    rand bit         io_writeback_21_bits_debug_isPerfCnt;
    rand bit [47:0]  io_writeback_21_bits_debug_paddr;
    rand bit [49:0]  io_writeback_21_bits_debug_vaddr;
    rand bit         io_writeback_21_bits_debugInfo_eliminatedMove;
    rand bit [63:0]  io_writeback_21_bits_debugInfo_renameTime;
    rand bit [63:0]  io_writeback_21_bits_debugInfo_dispatchTime;
    rand bit [63:0]  io_writeback_21_bits_debugInfo_enqRsTime;
    rand bit [63:0]  io_writeback_21_bits_debugInfo_selectTime;
    rand bit [63:0]  io_writeback_21_bits_debugInfo_issueTime;
    rand bit [63:0]  io_writeback_21_bits_debugInfo_writebackTime;
    rand bit [63:0]  io_writeback_21_bits_debugInfo_runahead_checkpoint_id;
    rand bit [63:0]  io_writeback_21_bits_debugInfo_tlbFirstReqTime;
    rand bit [63:0]  io_writeback_21_bits_debugInfo_tlbRespTime;
    rand bit [63:0]  io_writeback_21_bits_debug_seqNum;
    rand bit         io_writeback_20_valid;
    rand bit [63:0]  io_writeback_20_bits_data_0;
    rand bit [7:0]   io_writeback_20_bits_pdest;
    rand bit         io_writeback_20_bits_robIdx_flag;
    rand bit [7:0]   io_writeback_20_bits_robIdx_value;
    rand bit         io_writeback_20_bits_intWen;
    rand bit         io_writeback_20_bits_fpWen;
    rand bit         io_writeback_20_bits_exceptionVec_0;
    rand bit         io_writeback_20_bits_exceptionVec_1;
    rand bit         io_writeback_20_bits_exceptionVec_2;
    rand bit         io_writeback_20_bits_exceptionVec_3;
    rand bit         io_writeback_20_bits_exceptionVec_4;
    rand bit         io_writeback_20_bits_exceptionVec_5;
    rand bit         io_writeback_20_bits_exceptionVec_6;
    rand bit         io_writeback_20_bits_exceptionVec_7;
    rand bit         io_writeback_20_bits_exceptionVec_8;
    rand bit         io_writeback_20_bits_exceptionVec_9;
    rand bit         io_writeback_20_bits_exceptionVec_10;
    rand bit         io_writeback_20_bits_exceptionVec_11;
    rand bit         io_writeback_20_bits_exceptionVec_12;
    rand bit         io_writeback_20_bits_exceptionVec_13;
    rand bit         io_writeback_20_bits_exceptionVec_14;
    rand bit         io_writeback_20_bits_exceptionVec_15;
    rand bit         io_writeback_20_bits_exceptionVec_16;
    rand bit         io_writeback_20_bits_exceptionVec_17;
    rand bit         io_writeback_20_bits_exceptionVec_18;
    rand bit         io_writeback_20_bits_exceptionVec_19;
    rand bit         io_writeback_20_bits_exceptionVec_20;
    rand bit         io_writeback_20_bits_exceptionVec_21;
    rand bit         io_writeback_20_bits_exceptionVec_22;
    rand bit         io_writeback_20_bits_exceptionVec_23;
    rand bit         io_writeback_20_bits_flushPipe;
    rand bit         io_writeback_20_bits_replay;
    rand bit         io_writeback_20_bits_lqIdx_flag;
    rand bit [6:0]   io_writeback_20_bits_lqIdx_value;
    rand bit [3:0]   io_writeback_20_bits_trigger;
    rand bit         io_writeback_20_bits_predecodeInfo_valid;
    rand bit         io_writeback_20_bits_predecodeInfo_isRVC;
    rand bit [1:0]   io_writeback_20_bits_predecodeInfo_brType;
    rand bit         io_writeback_20_bits_predecodeInfo_isCall;
    rand bit         io_writeback_20_bits_predecodeInfo_isRet;
    rand bit         io_writeback_20_bits_debug_isMMIO;
    rand bit         io_writeback_20_bits_debug_isNCIO;
    rand bit         io_writeback_20_bits_debug_isPerfCnt;
    rand bit [47:0]  io_writeback_20_bits_debug_paddr;
    rand bit [49:0]  io_writeback_20_bits_debug_vaddr;
    rand bit         io_writeback_20_bits_debugInfo_eliminatedMove;
    rand bit [63:0]  io_writeback_20_bits_debugInfo_renameTime;
    rand bit [63:0]  io_writeback_20_bits_debugInfo_dispatchTime;
    rand bit [63:0]  io_writeback_20_bits_debugInfo_enqRsTime;
    rand bit [63:0]  io_writeback_20_bits_debugInfo_selectTime;
    rand bit [63:0]  io_writeback_20_bits_debugInfo_issueTime;
    rand bit [63:0]  io_writeback_20_bits_debugInfo_writebackTime;
    rand bit [63:0]  io_writeback_20_bits_debugInfo_runahead_checkpoint_id;
    rand bit [63:0]  io_writeback_20_bits_debugInfo_tlbFirstReqTime;
    rand bit [63:0]  io_writeback_20_bits_debugInfo_tlbRespTime;
    rand bit [63:0]  io_writeback_20_bits_debug_seqNum;
    rand bit         io_writeback_19_valid;
    rand bit [63:0]  io_writeback_19_bits_data_0;
    rand bit [7:0]   io_writeback_19_bits_pdest;
    rand bit         io_writeback_19_bits_robIdx_flag;
    rand bit [7:0]   io_writeback_19_bits_robIdx_value;
    rand bit         io_writeback_19_bits_intWen;
    rand bit         io_writeback_19_bits_exceptionVec_0;
    rand bit         io_writeback_19_bits_exceptionVec_1;
    rand bit         io_writeback_19_bits_exceptionVec_2;
    rand bit         io_writeback_19_bits_exceptionVec_3;
    rand bit         io_writeback_19_bits_exceptionVec_4;
    rand bit         io_writeback_19_bits_exceptionVec_5;
    rand bit         io_writeback_19_bits_exceptionVec_6;
    rand bit         io_writeback_19_bits_exceptionVec_7;
    rand bit         io_writeback_19_bits_exceptionVec_8;
    rand bit         io_writeback_19_bits_exceptionVec_9;
    rand bit         io_writeback_19_bits_exceptionVec_10;
    rand bit         io_writeback_19_bits_exceptionVec_11;
    rand bit         io_writeback_19_bits_exceptionVec_12;
    rand bit         io_writeback_19_bits_exceptionVec_13;
    rand bit         io_writeback_19_bits_exceptionVec_14;
    rand bit         io_writeback_19_bits_exceptionVec_15;
    rand bit         io_writeback_19_bits_exceptionVec_16;
    rand bit         io_writeback_19_bits_exceptionVec_17;
    rand bit         io_writeback_19_bits_exceptionVec_18;
    rand bit         io_writeback_19_bits_exceptionVec_19;
    rand bit         io_writeback_19_bits_exceptionVec_20;
    rand bit         io_writeback_19_bits_exceptionVec_21;
    rand bit         io_writeback_19_bits_exceptionVec_22;
    rand bit         io_writeback_19_bits_exceptionVec_23;
    rand bit         io_writeback_19_bits_flushPipe;
    rand bit         io_writeback_19_bits_sqIdx_flag;
    rand bit [5:0]   io_writeback_19_bits_sqIdx_value;
    rand bit [3:0]   io_writeback_19_bits_trigger;
    rand bit         io_writeback_19_bits_debug_isMMIO;
    rand bit         io_writeback_19_bits_debug_isNCIO;
    rand bit         io_writeback_19_bits_debug_isPerfCnt;
    rand bit [47:0]  io_writeback_19_bits_debug_paddr;
    rand bit [49:0]  io_writeback_19_bits_debug_vaddr;
    rand bit         io_writeback_19_bits_debugInfo_eliminatedMove;
    rand bit [63:0]  io_writeback_19_bits_debugInfo_renameTime;
    rand bit [63:0]  io_writeback_19_bits_debugInfo_dispatchTime;
    rand bit [63:0]  io_writeback_19_bits_debugInfo_enqRsTime;
    rand bit [63:0]  io_writeback_19_bits_debugInfo_selectTime;
    rand bit [63:0]  io_writeback_19_bits_debugInfo_issueTime;
    rand bit [63:0]  io_writeback_19_bits_debugInfo_writebackTime;
    rand bit [63:0]  io_writeback_19_bits_debugInfo_runahead_checkpoint_id;
    rand bit [63:0]  io_writeback_19_bits_debugInfo_tlbFirstReqTime;
    rand bit [63:0]  io_writeback_19_bits_debugInfo_tlbRespTime;
    rand bit [63:0]  io_writeback_19_bits_debug_seqNum;
    rand bit         io_writeback_18_valid;
    rand bit [63:0]  io_writeback_18_bits_data_0;
    rand bit [7:0]   io_writeback_18_bits_pdest;
    rand bit         io_writeback_18_bits_robIdx_flag;
    rand bit [7:0]   io_writeback_18_bits_robIdx_value;
    rand bit         io_writeback_18_bits_intWen;
    rand bit         io_writeback_18_bits_exceptionVec_0;
    rand bit         io_writeback_18_bits_exceptionVec_1;
    rand bit         io_writeback_18_bits_exceptionVec_2;
    rand bit         io_writeback_18_bits_exceptionVec_3;
    rand bit         io_writeback_18_bits_exceptionVec_4;
    rand bit         io_writeback_18_bits_exceptionVec_5;
    rand bit         io_writeback_18_bits_exceptionVec_6;
    rand bit         io_writeback_18_bits_exceptionVec_7;
    rand bit         io_writeback_18_bits_exceptionVec_8;
    rand bit         io_writeback_18_bits_exceptionVec_9;
    rand bit         io_writeback_18_bits_exceptionVec_10;
    rand bit         io_writeback_18_bits_exceptionVec_11;
    rand bit         io_writeback_18_bits_exceptionVec_12;
    rand bit         io_writeback_18_bits_exceptionVec_13;
    rand bit         io_writeback_18_bits_exceptionVec_14;
    rand bit         io_writeback_18_bits_exceptionVec_15;
    rand bit         io_writeback_18_bits_exceptionVec_16;
    rand bit         io_writeback_18_bits_exceptionVec_17;
    rand bit         io_writeback_18_bits_exceptionVec_18;
    rand bit         io_writeback_18_bits_exceptionVec_19;
    rand bit         io_writeback_18_bits_exceptionVec_20;
    rand bit         io_writeback_18_bits_exceptionVec_21;
    rand bit         io_writeback_18_bits_exceptionVec_22;
    rand bit         io_writeback_18_bits_exceptionVec_23;
    rand bit         io_writeback_18_bits_flushPipe;
    rand bit         io_writeback_18_bits_sqIdx_flag;
    rand bit [5:0]   io_writeback_18_bits_sqIdx_value;
    rand bit [3:0]   io_writeback_18_bits_trigger;
    rand bit         io_writeback_18_bits_debug_isMMIO;
    rand bit         io_writeback_18_bits_debug_isNCIO;
    rand bit         io_writeback_18_bits_debug_isPerfCnt;
    rand bit [47:0]  io_writeback_18_bits_debug_paddr;
    rand bit [49:0]  io_writeback_18_bits_debug_vaddr;
    rand bit         io_writeback_18_bits_debugInfo_eliminatedMove;
    rand bit [63:0]  io_writeback_18_bits_debugInfo_renameTime;
    rand bit [63:0]  io_writeback_18_bits_debugInfo_dispatchTime;
    rand bit [63:0]  io_writeback_18_bits_debugInfo_enqRsTime;
    rand bit [63:0]  io_writeback_18_bits_debugInfo_selectTime;
    rand bit [63:0]  io_writeback_18_bits_debugInfo_issueTime;
    rand bit [63:0]  io_writeback_18_bits_debugInfo_writebackTime;
    rand bit [63:0]  io_writeback_18_bits_debugInfo_runahead_checkpoint_id;
    rand bit [63:0]  io_writeback_18_bits_debugInfo_tlbFirstReqTime;
    rand bit [63:0]  io_writeback_18_bits_debugInfo_tlbRespTime;
    rand bit [63:0]  io_writeback_18_bits_debug_seqNum;
    rand bit         io_writeback_17_valid;
    rand bit [127:0] io_writeback_17_bits_data_0;
    rand bit [127:0] io_writeback_17_bits_data_1;
    rand bit [127:0] io_writeback_17_bits_data_2;
    rand bit [6:0]   io_writeback_17_bits_pdest;
    rand bit         io_writeback_17_bits_robIdx_flag;
    rand bit [7:0]   io_writeback_17_bits_robIdx_value;
    rand bit         io_writeback_17_bits_vecWen;
    rand bit         io_writeback_17_bits_v0Wen;
    rand bit [4:0]   io_writeback_17_bits_fflags;
    rand bit         io_writeback_17_bits_wflags;
    rand bit         io_writeback_17_bits_debugInfo_eliminatedMove;
    rand bit [63:0]  io_writeback_17_bits_debugInfo_renameTime;
    rand bit [63:0]  io_writeback_17_bits_debugInfo_dispatchTime;
    rand bit [63:0]  io_writeback_17_bits_debugInfo_enqRsTime;
    rand bit [63:0]  io_writeback_17_bits_debugInfo_selectTime;
    rand bit [63:0]  io_writeback_17_bits_debugInfo_issueTime;
    rand bit [63:0]  io_writeback_17_bits_debugInfo_writebackTime;
    rand bit [63:0]  io_writeback_17_bits_debugInfo_runahead_checkpoint_id;
    rand bit [63:0]  io_writeback_17_bits_debugInfo_tlbFirstReqTime;
    rand bit [63:0]  io_writeback_17_bits_debugInfo_tlbRespTime;
    rand bit [63:0]  io_writeback_17_bits_debug_seqNum;
    rand bit         io_writeback_16_valid;
    rand bit [127:0] io_writeback_16_bits_data_0;
    rand bit [127:0] io_writeback_16_bits_data_1;
    rand bit [127:0] io_writeback_16_bits_data_2;
    rand bit [127:0] io_writeback_16_bits_data_3;
    rand bit [7:0]   io_writeback_16_bits_pdest;
    rand bit         io_writeback_16_bits_robIdx_flag;
    rand bit [7:0]   io_writeback_16_bits_robIdx_value;
    rand bit         io_writeback_16_bits_fpWen;
    rand bit         io_writeback_16_bits_vecWen;
    rand bit         io_writeback_16_bits_v0Wen;
    rand bit [4:0]   io_writeback_16_bits_fflags;
    rand bit         io_writeback_16_bits_wflags;
    rand bit         io_writeback_16_bits_debugInfo_eliminatedMove;
    rand bit [63:0]  io_writeback_16_bits_debugInfo_renameTime;
    rand bit [63:0]  io_writeback_16_bits_debugInfo_dispatchTime;
    rand bit [63:0]  io_writeback_16_bits_debugInfo_enqRsTime;
    rand bit [63:0]  io_writeback_16_bits_debugInfo_selectTime;
    rand bit [63:0]  io_writeback_16_bits_debugInfo_issueTime;
    rand bit [63:0]  io_writeback_16_bits_debugInfo_writebackTime;
    rand bit [63:0]  io_writeback_16_bits_debugInfo_runahead_checkpoint_id;
    rand bit [63:0]  io_writeback_16_bits_debugInfo_tlbFirstReqTime;
    rand bit [63:0]  io_writeback_16_bits_debugInfo_tlbRespTime;
    rand bit [63:0]  io_writeback_16_bits_debug_seqNum;
    rand bit         io_writeback_15_valid;
    rand bit [127:0] io_writeback_15_bits_data_0;
    rand bit [127:0] io_writeback_15_bits_data_1;
    rand bit [127:0] io_writeback_15_bits_data_2;
    rand bit [6:0]   io_writeback_15_bits_pdest;
    rand bit         io_writeback_15_bits_robIdx_flag;
    rand bit [7:0]   io_writeback_15_bits_robIdx_value;
    rand bit         io_writeback_15_bits_vecWen;
    rand bit         io_writeback_15_bits_v0Wen;
    rand bit [4:0]   io_writeback_15_bits_fflags;
    rand bit         io_writeback_15_bits_wflags;
    rand bit         io_writeback_15_bits_vxsat;
    rand bit         io_writeback_15_bits_debugInfo_eliminatedMove;
    rand bit [63:0]  io_writeback_15_bits_debugInfo_renameTime;
    rand bit [63:0]  io_writeback_15_bits_debugInfo_dispatchTime;
    rand bit [63:0]  io_writeback_15_bits_debugInfo_enqRsTime;
    rand bit [63:0]  io_writeback_15_bits_debugInfo_selectTime;
    rand bit [63:0]  io_writeback_15_bits_debugInfo_issueTime;
    rand bit [63:0]  io_writeback_15_bits_debugInfo_writebackTime;
    rand bit [63:0]  io_writeback_15_bits_debugInfo_runahead_checkpoint_id;
    rand bit [63:0]  io_writeback_15_bits_debugInfo_tlbFirstReqTime;
    rand bit [63:0]  io_writeback_15_bits_debugInfo_tlbRespTime;
    rand bit [63:0]  io_writeback_15_bits_debug_seqNum;
    rand bit         io_writeback_14_valid;
    rand bit [127:0] io_writeback_14_bits_data_0;
    rand bit [127:0] io_writeback_14_bits_data_1;
    rand bit [127:0] io_writeback_14_bits_data_2;
    rand bit [127:0] io_writeback_14_bits_data_3;
    rand bit [127:0] io_writeback_14_bits_data_4;
    rand bit [127:0] io_writeback_14_bits_data_5;
    rand bit [7:0]   io_writeback_14_bits_pdest;
    rand bit         io_writeback_14_bits_robIdx_flag;
    rand bit [7:0]   io_writeback_14_bits_robIdx_value;
    rand bit         io_writeback_14_bits_intWen;
    rand bit         io_writeback_14_bits_fpWen;
    rand bit         io_writeback_14_bits_vecWen;
    rand bit         io_writeback_14_bits_v0Wen;
    rand bit         io_writeback_14_bits_vlWen;
    rand bit [4:0]   io_writeback_14_bits_fflags;
    rand bit         io_writeback_14_bits_wflags;
    rand bit         io_writeback_14_bits_exceptionVec_2;
    rand bit         io_writeback_14_bits_debugInfo_eliminatedMove;
    rand bit [63:0]  io_writeback_14_bits_debugInfo_renameTime;
    rand bit [63:0]  io_writeback_14_bits_debugInfo_dispatchTime;
    rand bit [63:0]  io_writeback_14_bits_debugInfo_enqRsTime;
    rand bit [63:0]  io_writeback_14_bits_debugInfo_selectTime;
    rand bit [63:0]  io_writeback_14_bits_debugInfo_issueTime;
    rand bit [63:0]  io_writeback_14_bits_debugInfo_writebackTime;
    rand bit [63:0]  io_writeback_14_bits_debugInfo_runahead_checkpoint_id;
    rand bit [63:0]  io_writeback_14_bits_debugInfo_tlbFirstReqTime;
    rand bit [63:0]  io_writeback_14_bits_debugInfo_tlbRespTime;
    rand bit [63:0]  io_writeback_14_bits_debug_seqNum;
    rand bit         io_writeback_13_valid;
    rand bit [127:0] io_writeback_13_bits_data_0;
    rand bit [127:0] io_writeback_13_bits_data_1;
    rand bit [127:0] io_writeback_13_bits_data_2;
    rand bit [6:0]   io_writeback_13_bits_pdest;
    rand bit         io_writeback_13_bits_robIdx_flag;
    rand bit [7:0]   io_writeback_13_bits_robIdx_value;
    rand bit         io_writeback_13_bits_vecWen;
    rand bit         io_writeback_13_bits_v0Wen;
    rand bit [4:0]   io_writeback_13_bits_fflags;
    rand bit         io_writeback_13_bits_wflags;
    rand bit         io_writeback_13_bits_vxsat;
    rand bit         io_writeback_13_bits_exceptionVec_2;
    rand bit         io_writeback_13_bits_debugInfo_eliminatedMove;
    rand bit [63:0]  io_writeback_13_bits_debugInfo_renameTime;
    rand bit [63:0]  io_writeback_13_bits_debugInfo_dispatchTime;
    rand bit [63:0]  io_writeback_13_bits_debugInfo_enqRsTime;
    rand bit [63:0]  io_writeback_13_bits_debugInfo_selectTime;
    rand bit [63:0]  io_writeback_13_bits_debugInfo_issueTime;
    rand bit [63:0]  io_writeback_13_bits_debugInfo_writebackTime;
    rand bit [63:0]  io_writeback_13_bits_debugInfo_runahead_checkpoint_id;
    rand bit [63:0]  io_writeback_13_bits_debugInfo_tlbFirstReqTime;
    rand bit [63:0]  io_writeback_13_bits_debugInfo_tlbRespTime;
    rand bit [63:0]  io_writeback_13_bits_debug_seqNum;
    rand bit         io_writeback_7_valid;
    rand bit [63:0]  io_writeback_7_bits_data_0;
    rand bit [63:0]  io_writeback_7_bits_data_1;
    rand bit [7:0]   io_writeback_7_bits_pdest;
    rand bit         io_writeback_7_bits_robIdx_flag;
    rand bit [7:0]   io_writeback_7_bits_robIdx_value;
    rand bit         io_writeback_7_bits_intWen;
    rand bit         io_writeback_7_bits_redirect_valid;
    rand bit         io_writeback_7_bits_redirect_bits_isRVC;
    rand bit         io_writeback_7_bits_redirect_bits_robIdx_flag;
    rand bit [7:0]   io_writeback_7_bits_redirect_bits_robIdx_value;
    rand bit         io_writeback_7_bits_redirect_bits_ftqIdx_flag;
    rand bit [5:0]   io_writeback_7_bits_redirect_bits_ftqIdx_value;
    rand bit [3:0]   io_writeback_7_bits_redirect_bits_ftqOffset;
    rand bit         io_writeback_7_bits_redirect_bits_level;
    rand bit         io_writeback_7_bits_redirect_bits_interrupt;
    rand bit [49:0]  io_writeback_7_bits_redirect_bits_cfiUpdate_pc;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC;
    rand bit [1:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet;
    rand bit [3:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_ssp;
    rand bit [2:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_sctr;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag;
    rand bit [4:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag;
    rand bit [4:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag;
    rand bit [4:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value;
    rand bit [49:0]  io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr;
    rand bit [10:0]  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist;
    rand bit [10:0]  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist;
    rand bit [6:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist;
    rand bit [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist;
    rand bit [8:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist;
    rand bit [3:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist;
    rand bit [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist;
    rand bit [8:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist;
    rand bit [6:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist;
    rand bit [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist;
    rand bit [6:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist;
    rand bit [8:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist;
    rand bit [6:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist;
    rand bit [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist;
    rand bit [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist;
    rand bit [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist;
    rand bit [10:0]  io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist;
    rand bit [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3;
    rand bit [2:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH;
    rand bit [3:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_ghr;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag;
    rand bit [7:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value;
    rand bit [9:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0;
    rand bit [9:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken;
    rand bit [49:0]  io_writeback_7_bits_redirect_bits_cfiUpdate_target;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_taken;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred;
    rand bit [1:0]   io_writeback_7_bits_redirect_bits_cfiUpdate_shift;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF;
    rand bit         io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF;
    rand bit [63:0]  io_writeback_7_bits_redirect_bits_fullTarget;
    rand bit         io_writeback_7_bits_redirect_bits_stFtqIdx_flag;
    rand bit [5:0]   io_writeback_7_bits_redirect_bits_stFtqIdx_value;
    rand bit [3:0]   io_writeback_7_bits_redirect_bits_stFtqOffset;
    rand bit [63:0]  io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id;
    rand bit         io_writeback_7_bits_redirect_bits_debugIsCtrl;
    rand bit         io_writeback_7_bits_redirect_bits_debugIsMemVio;
    rand bit         io_writeback_7_bits_exceptionVec_2;
    rand bit         io_writeback_7_bits_exceptionVec_3;
    rand bit         io_writeback_7_bits_exceptionVec_8;
    rand bit         io_writeback_7_bits_exceptionVec_9;
    rand bit         io_writeback_7_bits_exceptionVec_10;
    rand bit         io_writeback_7_bits_exceptionVec_11;
    rand bit         io_writeback_7_bits_exceptionVec_22;
    rand bit         io_writeback_7_bits_flushPipe;
    rand bit         io_writeback_7_bits_predecodeInfo_valid;
    rand bit         io_writeback_7_bits_predecodeInfo_isRVC;
    rand bit [1:0]   io_writeback_7_bits_predecodeInfo_brType;
    rand bit         io_writeback_7_bits_predecodeInfo_isCall;
    rand bit         io_writeback_7_bits_predecodeInfo_isRet;
    rand bit         io_writeback_7_bits_debug_isPerfCnt;
    rand bit         io_writeback_7_bits_debugInfo_eliminatedMove;
    rand bit [63:0]  io_writeback_7_bits_debugInfo_renameTime;
    rand bit [63:0]  io_writeback_7_bits_debugInfo_dispatchTime;
    rand bit [63:0]  io_writeback_7_bits_debugInfo_enqRsTime;
    rand bit [63:0]  io_writeback_7_bits_debugInfo_selectTime;
    rand bit [63:0]  io_writeback_7_bits_debugInfo_issueTime;
    rand bit [63:0]  io_writeback_7_bits_debugInfo_writebackTime;
    rand bit [63:0]  io_writeback_7_bits_debugInfo_runahead_checkpoint_id;
    rand bit [63:0]  io_writeback_7_bits_debugInfo_tlbFirstReqTime;
    rand bit [63:0]  io_writeback_7_bits_debugInfo_tlbRespTime;
    rand bit [63:0]  io_writeback_7_bits_debug_seqNum;
    rand bit         io_writeback_5_valid;
    rand bit         io_writeback_5_bits_redirect_valid;
    rand bit         io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred;
    rand bit         io_writeback_3_valid;
    rand bit         io_writeback_3_bits_redirect_valid;
    rand bit         io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred;
    rand bit         io_writeback_1_valid;
    rand bit         io_writeback_1_bits_redirect_valid;
    rand bit         io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred;
    rand bit         io_exuWriteback_26_valid;
    rand bit [7:0]   io_exuWriteback_26_bits_robIdx_value;
    rand bit         io_exuWriteback_25_valid;
    rand bit [7:0]   io_exuWriteback_25_bits_robIdx_value;
    rand bit         io_exuWriteback_24_valid;
    rand bit [127:0] io_exuWriteback_24_bits_data_0;
    rand bit [6:0]   io_exuWriteback_24_bits_pdest;
    rand bit [7:0]   io_exuWriteback_24_bits_robIdx_value;
    rand bit         io_exuWriteback_24_bits_vecWen;
    rand bit         io_exuWriteback_24_bits_v0Wen;
    rand bit [2:0]   io_exuWriteback_24_bits_vls_vdIdx;
    rand bit         io_exuWriteback_24_bits_debug_isMMIO;
    rand bit         io_exuWriteback_24_bits_debug_isNCIO;
    rand bit         io_exuWriteback_24_bits_debug_isPerfCnt;
    rand bit [47:0]  io_exuWriteback_24_bits_debug_paddr;
    rand bit         io_exuWriteback_23_valid;
    rand bit [127:0] io_exuWriteback_23_bits_data_0;
    rand bit [6:0]   io_exuWriteback_23_bits_pdest;
    rand bit [7:0]   io_exuWriteback_23_bits_robIdx_value;
    rand bit         io_exuWriteback_23_bits_vecWen;
    rand bit         io_exuWriteback_23_bits_v0Wen;
    rand bit [2:0]   io_exuWriteback_23_bits_vls_vdIdx;
    rand bit         io_exuWriteback_23_bits_debug_isMMIO;
    rand bit         io_exuWriteback_23_bits_debug_isNCIO;
    rand bit         io_exuWriteback_23_bits_debug_isPerfCnt;
    rand bit [47:0]  io_exuWriteback_23_bits_debug_paddr;
    rand bit         io_exuWriteback_22_valid;
    rand bit [63:0]  io_exuWriteback_22_bits_data_0;
    rand bit [7:0]   io_exuWriteback_22_bits_robIdx_value;
    rand bit [6:0]   io_exuWriteback_22_bits_lqIdx_value;
    rand bit         io_exuWriteback_22_bits_debug_isMMIO;
    rand bit         io_exuWriteback_22_bits_debug_isNCIO;
    rand bit         io_exuWriteback_22_bits_debug_isPerfCnt;
    rand bit [47:0]  io_exuWriteback_22_bits_debug_paddr;
    rand bit         io_exuWriteback_21_valid;
    rand bit [63:0]  io_exuWriteback_21_bits_data_0;
    rand bit [7:0]   io_exuWriteback_21_bits_robIdx_value;
    rand bit [6:0]   io_exuWriteback_21_bits_lqIdx_value;
    rand bit         io_exuWriteback_21_bits_debug_isMMIO;
    rand bit         io_exuWriteback_21_bits_debug_isNCIO;
    rand bit         io_exuWriteback_21_bits_debug_isPerfCnt;
    rand bit [47:0]  io_exuWriteback_21_bits_debug_paddr;
    rand bit         io_exuWriteback_20_valid;
    rand bit [63:0]  io_exuWriteback_20_bits_data_0;
    rand bit [7:0]   io_exuWriteback_20_bits_robIdx_value;
    rand bit [6:0]   io_exuWriteback_20_bits_lqIdx_value;
    rand bit         io_exuWriteback_20_bits_debug_isMMIO;
    rand bit         io_exuWriteback_20_bits_debug_isNCIO;
    rand bit         io_exuWriteback_20_bits_debug_isPerfCnt;
    rand bit [47:0]  io_exuWriteback_20_bits_debug_paddr;
    rand bit         io_exuWriteback_19_valid;
    rand bit [63:0]  io_exuWriteback_19_bits_data_0;
    rand bit [7:0]   io_exuWriteback_19_bits_robIdx_value;
    rand bit [5:0]   io_exuWriteback_19_bits_sqIdx_value;
    rand bit         io_exuWriteback_19_bits_debug_isMMIO;
    rand bit         io_exuWriteback_19_bits_debug_isNCIO;
    rand bit         io_exuWriteback_19_bits_debug_isPerfCnt;
    rand bit [47:0]  io_exuWriteback_19_bits_debug_paddr;
    rand bit         io_exuWriteback_18_valid;
    rand bit [63:0]  io_exuWriteback_18_bits_data_0;
    rand bit [7:0]   io_exuWriteback_18_bits_robIdx_value;
    rand bit [5:0]   io_exuWriteback_18_bits_sqIdx_value;
    rand bit         io_exuWriteback_18_bits_debug_isMMIO;
    rand bit         io_exuWriteback_18_bits_debug_isNCIO;
    rand bit         io_exuWriteback_18_bits_debug_isPerfCnt;
    rand bit [47:0]  io_exuWriteback_18_bits_debug_paddr;
    rand bit         io_exuWriteback_17_valid;
    rand bit [127:0] io_exuWriteback_17_bits_data_0;
    rand bit [7:0]   io_exuWriteback_17_bits_robIdx_value;
    rand bit [4:0]   io_exuWriteback_17_bits_fflags;
    rand bit         io_exuWriteback_17_bits_wflags;
    rand bit         io_exuWriteback_16_valid;
    rand bit [127:0] io_exuWriteback_16_bits_data_0;
    rand bit [7:0]   io_exuWriteback_16_bits_robIdx_value;
    rand bit [4:0]   io_exuWriteback_16_bits_fflags;
    rand bit         io_exuWriteback_16_bits_wflags;
    rand bit         io_exuWriteback_15_valid;
    rand bit [127:0] io_exuWriteback_15_bits_data_0;
    rand bit [7:0]   io_exuWriteback_15_bits_robIdx_value;
    rand bit [4:0]   io_exuWriteback_15_bits_fflags;
    rand bit         io_exuWriteback_15_bits_wflags;
    rand bit         io_exuWriteback_15_bits_vxsat;
    rand bit         io_exuWriteback_14_valid;
    rand bit [127:0] io_exuWriteback_14_bits_data_0;
    rand bit [7:0]   io_exuWriteback_14_bits_robIdx_value;
    rand bit [4:0]   io_exuWriteback_14_bits_fflags;
    rand bit         io_exuWriteback_14_bits_wflags;
    rand bit         io_exuWriteback_13_valid;
    rand bit [127:0] io_exuWriteback_13_bits_data_0;
    rand bit [7:0]   io_exuWriteback_13_bits_robIdx_value;
    rand bit [4:0]   io_exuWriteback_13_bits_fflags;
    rand bit         io_exuWriteback_13_bits_wflags;
    rand bit         io_exuWriteback_13_bits_vxsat;
    rand bit         io_exuWriteback_12_valid;
    rand bit [63:0]  io_exuWriteback_12_bits_data_0;
    rand bit [7:0]   io_exuWriteback_12_bits_robIdx_value;
    rand bit [4:0]   io_exuWriteback_12_bits_fflags;
    rand bit         io_exuWriteback_12_bits_wflags;
    rand bit         io_exuWriteback_11_valid;
    rand bit [63:0]  io_exuWriteback_11_bits_data_0;
    rand bit [7:0]   io_exuWriteback_11_bits_robIdx_value;
    rand bit [4:0]   io_exuWriteback_11_bits_fflags;
    rand bit         io_exuWriteback_11_bits_wflags;
    rand bit         io_exuWriteback_10_valid;
    rand bit [63:0]  io_exuWriteback_10_bits_data_0;
    rand bit [7:0]   io_exuWriteback_10_bits_robIdx_value;
    rand bit [4:0]   io_exuWriteback_10_bits_fflags;
    rand bit         io_exuWriteback_10_bits_wflags;
    rand bit         io_exuWriteback_9_valid;
    rand bit [63:0]  io_exuWriteback_9_bits_data_0;
    rand bit [7:0]   io_exuWriteback_9_bits_robIdx_value;
    rand bit [4:0]   io_exuWriteback_9_bits_fflags;
    rand bit         io_exuWriteback_9_bits_wflags;
    rand bit         io_exuWriteback_8_valid;
    rand bit [127:0] io_exuWriteback_8_bits_data_0;
    rand bit [7:0]   io_exuWriteback_8_bits_robIdx_value;
    rand bit [4:0]   io_exuWriteback_8_bits_fflags;
    rand bit         io_exuWriteback_8_bits_wflags;
    rand bit         io_exuWriteback_7_valid;
    rand bit [63:0]  io_exuWriteback_7_bits_data_0;
    rand bit [7:0]   io_exuWriteback_7_bits_robIdx_value;
    rand bit         io_exuWriteback_7_bits_debug_isPerfCnt;
    rand bit         io_exuWriteback_6_valid;
    rand bit [63:0]  io_exuWriteback_6_bits_data_0;
    rand bit [7:0]   io_exuWriteback_6_bits_robIdx_value;
    rand bit         io_exuWriteback_5_valid;
    rand bit [127:0] io_exuWriteback_5_bits_data_0;
    rand bit [7:0]   io_exuWriteback_5_bits_robIdx_value;
    rand bit         io_exuWriteback_5_bits_redirect_valid;
    rand bit         io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken;
    rand bit [4:0]   io_exuWriteback_5_bits_fflags;
    rand bit         io_exuWriteback_5_bits_wflags;
    rand bit         io_exuWriteback_4_valid;
    rand bit [63:0]  io_exuWriteback_4_bits_data_0;
    rand bit [7:0]   io_exuWriteback_4_bits_robIdx_value;
    rand bit         io_exuWriteback_3_valid;
    rand bit [63:0]  io_exuWriteback_3_bits_data_0;
    rand bit [7:0]   io_exuWriteback_3_bits_robIdx_value;
    rand bit         io_exuWriteback_3_bits_redirect_valid;
    rand bit         io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken;
    rand bit         io_exuWriteback_2_valid;
    rand bit [63:0]  io_exuWriteback_2_bits_data_0;
    rand bit [7:0]   io_exuWriteback_2_bits_robIdx_value;
    rand bit         io_exuWriteback_1_valid;
    rand bit [63:0]  io_exuWriteback_1_bits_data_0;
    rand bit [7:0]   io_exuWriteback_1_bits_robIdx_value;
    rand bit         io_exuWriteback_1_bits_redirect_valid;
    rand bit         io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken;
    rand bit         io_exuWriteback_0_valid;
    rand bit [63:0]  io_exuWriteback_0_bits_data_0;
    rand bit [7:0]   io_exuWriteback_0_bits_robIdx_value;
    rand bit [4:0]   io_writebackNums_0_bits;
    rand bit [4:0]   io_writebackNums_1_bits;
    rand bit [4:0]   io_writebackNums_2_bits;
    rand bit [4:0]   io_writebackNums_3_bits;
    rand bit [4:0]   io_writebackNums_4_bits;
    rand bit [4:0]   io_writebackNums_5_bits;
    rand bit [4:0]   io_writebackNums_6_bits;
    rand bit [4:0]   io_writebackNums_7_bits;
    rand bit [4:0]   io_writebackNums_8_bits;
    rand bit [4:0]   io_writebackNums_9_bits;
    rand bit [4:0]   io_writebackNums_10_bits;
    rand bit [4:0]   io_writebackNums_11_bits;
    rand bit [4:0]   io_writebackNums_12_bits;
    rand bit [4:0]   io_writebackNums_13_bits;
    rand bit [4:0]   io_writebackNums_14_bits;
    rand bit [4:0]   io_writebackNums_15_bits;
    rand bit [4:0]   io_writebackNums_16_bits;
    rand bit [4:0]   io_writebackNums_17_bits;
    rand bit [4:0]   io_writebackNums_18_bits;
    rand bit [4:0]   io_writebackNums_19_bits;
    rand bit [4:0]   io_writebackNums_20_bits;
    rand bit [4:0]   io_writebackNums_21_bits;
    rand bit [4:0]   io_writebackNums_22_bits;
    rand bit [4:0]   io_writebackNums_23_bits;
    rand bit [4:0]   io_writebackNums_24_bits;
    rand bit         io_writebackNeedFlush_0;
    rand bit         io_writebackNeedFlush_1;
    rand bit         io_writebackNeedFlush_2;
    rand bit         io_writebackNeedFlush_6;
    rand bit         io_writebackNeedFlush_7;
    rand bit         io_writebackNeedFlush_8;
    rand bit         io_writebackNeedFlush_9;
    rand bit         io_writebackNeedFlush_10;
    rand bit         io_writebackNeedFlush_11;
    rand bit         io_writebackNeedFlush_12;

    extern constraint default_io_writeback_24_valid_cons;
    extern constraint default_io_writeback_24_bits_data_0_cons;
    extern constraint default_io_writeback_24_bits_pdest_cons;
    extern constraint default_io_writeback_24_bits_robIdx_flag_cons;
    extern constraint default_io_writeback_24_bits_robIdx_value_cons;
    extern constraint default_io_writeback_24_bits_vecWen_cons;
    extern constraint default_io_writeback_24_bits_v0Wen_cons;
    extern constraint default_io_writeback_24_bits_vlWen_cons;
    extern constraint default_io_writeback_24_bits_exceptionVec_0_cons;
    extern constraint default_io_writeback_24_bits_exceptionVec_1_cons;
    extern constraint default_io_writeback_24_bits_exceptionVec_2_cons;
    extern constraint default_io_writeback_24_bits_exceptionVec_3_cons;
    extern constraint default_io_writeback_24_bits_exceptionVec_4_cons;
    extern constraint default_io_writeback_24_bits_exceptionVec_5_cons;
    extern constraint default_io_writeback_24_bits_exceptionVec_6_cons;
    extern constraint default_io_writeback_24_bits_exceptionVec_7_cons;
    extern constraint default_io_writeback_24_bits_exceptionVec_8_cons;
    extern constraint default_io_writeback_24_bits_exceptionVec_9_cons;
    extern constraint default_io_writeback_24_bits_exceptionVec_10_cons;
    extern constraint default_io_writeback_24_bits_exceptionVec_11_cons;
    extern constraint default_io_writeback_24_bits_exceptionVec_12_cons;
    extern constraint default_io_writeback_24_bits_exceptionVec_13_cons;
    extern constraint default_io_writeback_24_bits_exceptionVec_14_cons;
    extern constraint default_io_writeback_24_bits_exceptionVec_15_cons;
    extern constraint default_io_writeback_24_bits_exceptionVec_16_cons;
    extern constraint default_io_writeback_24_bits_exceptionVec_17_cons;
    extern constraint default_io_writeback_24_bits_exceptionVec_18_cons;
    extern constraint default_io_writeback_24_bits_exceptionVec_19_cons;
    extern constraint default_io_writeback_24_bits_exceptionVec_20_cons;
    extern constraint default_io_writeback_24_bits_exceptionVec_21_cons;
    extern constraint default_io_writeback_24_bits_exceptionVec_22_cons;
    extern constraint default_io_writeback_24_bits_exceptionVec_23_cons;
    extern constraint default_io_writeback_24_bits_flushPipe_cons;
    extern constraint default_io_writeback_24_bits_replay_cons;
    extern constraint default_io_writeback_24_bits_trigger_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_vill_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_vma_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_vta_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_vsew_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_vlmul_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_specVill_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_specVma_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_specVta_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_specVsew_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_specVlmul_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_vm_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_vstart_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_frm_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_fpu_isFP32Instr_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_fpu_isFP64Instr_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_fpu_isReduction_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_vxrm_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_vuopIdx_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_lastUop_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_vmask_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_vl_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_nf_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_veew_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_isReverse_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_isExt_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_isNarrow_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_isDstMask_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_isOpMask_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_isMove_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_isDependOldVd_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_isWritePartVd_cons;
    extern constraint default_io_writeback_24_bits_vls_vpu_isVleff_cons;
    extern constraint default_io_writeback_24_bits_vls_oldVdPsrc_cons;
    extern constraint default_io_writeback_24_bits_vls_vdIdx_cons;
    extern constraint default_io_writeback_24_bits_vls_vdIdxInField_cons;
    extern constraint default_io_writeback_24_bits_vls_isIndexed_cons;
    extern constraint default_io_writeback_24_bits_vls_isMasked_cons;
    extern constraint default_io_writeback_24_bits_vls_isStrided_cons;
    extern constraint default_io_writeback_24_bits_vls_isWhole_cons;
    extern constraint default_io_writeback_24_bits_vls_isVecLoad_cons;
    extern constraint default_io_writeback_24_bits_vls_isVlm_cons;
    extern constraint default_io_writeback_24_bits_debug_isMMIO_cons;
    extern constraint default_io_writeback_24_bits_debug_isNCIO_cons;
    extern constraint default_io_writeback_24_bits_debug_isPerfCnt_cons;
    extern constraint default_io_writeback_24_bits_debug_paddr_cons;
    extern constraint default_io_writeback_24_bits_debug_vaddr_cons;
    extern constraint default_io_writeback_24_bits_debugInfo_eliminatedMove_cons;
    extern constraint default_io_writeback_24_bits_debugInfo_renameTime_cons;
    extern constraint default_io_writeback_24_bits_debugInfo_dispatchTime_cons;
    extern constraint default_io_writeback_24_bits_debugInfo_enqRsTime_cons;
    extern constraint default_io_writeback_24_bits_debugInfo_selectTime_cons;
    extern constraint default_io_writeback_24_bits_debugInfo_issueTime_cons;
    extern constraint default_io_writeback_24_bits_debugInfo_writebackTime_cons;
    extern constraint default_io_writeback_24_bits_debugInfo_runahead_checkpoint_id_cons;
    extern constraint default_io_writeback_24_bits_debugInfo_tlbFirstReqTime_cons;
    extern constraint default_io_writeback_24_bits_debugInfo_tlbRespTime_cons;
    extern constraint default_io_writeback_24_bits_debug_seqNum_cons;
    extern constraint default_io_writeback_23_valid_cons;
    extern constraint default_io_writeback_23_bits_data_0_cons;
    extern constraint default_io_writeback_23_bits_pdest_cons;
    extern constraint default_io_writeback_23_bits_robIdx_flag_cons;
    extern constraint default_io_writeback_23_bits_robIdx_value_cons;
    extern constraint default_io_writeback_23_bits_vecWen_cons;
    extern constraint default_io_writeback_23_bits_v0Wen_cons;
    extern constraint default_io_writeback_23_bits_vlWen_cons;
    extern constraint default_io_writeback_23_bits_exceptionVec_0_cons;
    extern constraint default_io_writeback_23_bits_exceptionVec_1_cons;
    extern constraint default_io_writeback_23_bits_exceptionVec_2_cons;
    extern constraint default_io_writeback_23_bits_exceptionVec_3_cons;
    extern constraint default_io_writeback_23_bits_exceptionVec_4_cons;
    extern constraint default_io_writeback_23_bits_exceptionVec_5_cons;
    extern constraint default_io_writeback_23_bits_exceptionVec_6_cons;
    extern constraint default_io_writeback_23_bits_exceptionVec_7_cons;
    extern constraint default_io_writeback_23_bits_exceptionVec_8_cons;
    extern constraint default_io_writeback_23_bits_exceptionVec_9_cons;
    extern constraint default_io_writeback_23_bits_exceptionVec_10_cons;
    extern constraint default_io_writeback_23_bits_exceptionVec_11_cons;
    extern constraint default_io_writeback_23_bits_exceptionVec_12_cons;
    extern constraint default_io_writeback_23_bits_exceptionVec_13_cons;
    extern constraint default_io_writeback_23_bits_exceptionVec_14_cons;
    extern constraint default_io_writeback_23_bits_exceptionVec_15_cons;
    extern constraint default_io_writeback_23_bits_exceptionVec_16_cons;
    extern constraint default_io_writeback_23_bits_exceptionVec_17_cons;
    extern constraint default_io_writeback_23_bits_exceptionVec_18_cons;
    extern constraint default_io_writeback_23_bits_exceptionVec_19_cons;
    extern constraint default_io_writeback_23_bits_exceptionVec_20_cons;
    extern constraint default_io_writeback_23_bits_exceptionVec_21_cons;
    extern constraint default_io_writeback_23_bits_exceptionVec_22_cons;
    extern constraint default_io_writeback_23_bits_exceptionVec_23_cons;
    extern constraint default_io_writeback_23_bits_flushPipe_cons;
    extern constraint default_io_writeback_23_bits_replay_cons;
    extern constraint default_io_writeback_23_bits_trigger_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_vill_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_vma_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_vta_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_vsew_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_vlmul_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_specVill_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_specVma_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_specVta_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_specVsew_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_specVlmul_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_vm_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_vstart_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_frm_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_fpu_isFP32Instr_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_fpu_isFP64Instr_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_fpu_isReduction_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_vxrm_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_vuopIdx_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_lastUop_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_vmask_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_vl_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_nf_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_veew_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_isReverse_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_isExt_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_isNarrow_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_isDstMask_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_isOpMask_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_isMove_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_isDependOldVd_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_isWritePartVd_cons;
    extern constraint default_io_writeback_23_bits_vls_vpu_isVleff_cons;
    extern constraint default_io_writeback_23_bits_vls_oldVdPsrc_cons;
    extern constraint default_io_writeback_23_bits_vls_vdIdx_cons;
    extern constraint default_io_writeback_23_bits_vls_vdIdxInField_cons;
    extern constraint default_io_writeback_23_bits_vls_isIndexed_cons;
    extern constraint default_io_writeback_23_bits_vls_isMasked_cons;
    extern constraint default_io_writeback_23_bits_vls_isStrided_cons;
    extern constraint default_io_writeback_23_bits_vls_isWhole_cons;
    extern constraint default_io_writeback_23_bits_vls_isVecLoad_cons;
    extern constraint default_io_writeback_23_bits_vls_isVlm_cons;
    extern constraint default_io_writeback_23_bits_debug_isMMIO_cons;
    extern constraint default_io_writeback_23_bits_debug_isNCIO_cons;
    extern constraint default_io_writeback_23_bits_debug_isPerfCnt_cons;
    extern constraint default_io_writeback_23_bits_debug_paddr_cons;
    extern constraint default_io_writeback_23_bits_debug_vaddr_cons;
    extern constraint default_io_writeback_23_bits_debugInfo_eliminatedMove_cons;
    extern constraint default_io_writeback_23_bits_debugInfo_renameTime_cons;
    extern constraint default_io_writeback_23_bits_debugInfo_dispatchTime_cons;
    extern constraint default_io_writeback_23_bits_debugInfo_enqRsTime_cons;
    extern constraint default_io_writeback_23_bits_debugInfo_selectTime_cons;
    extern constraint default_io_writeback_23_bits_debugInfo_issueTime_cons;
    extern constraint default_io_writeback_23_bits_debugInfo_writebackTime_cons;
    extern constraint default_io_writeback_23_bits_debugInfo_runahead_checkpoint_id_cons;
    extern constraint default_io_writeback_23_bits_debugInfo_tlbFirstReqTime_cons;
    extern constraint default_io_writeback_23_bits_debugInfo_tlbRespTime_cons;
    extern constraint default_io_writeback_23_bits_debug_seqNum_cons;
    extern constraint default_io_writeback_22_valid_cons;
    extern constraint default_io_writeback_22_bits_data_0_cons;
    extern constraint default_io_writeback_22_bits_pdest_cons;
    extern constraint default_io_writeback_22_bits_robIdx_flag_cons;
    extern constraint default_io_writeback_22_bits_robIdx_value_cons;
    extern constraint default_io_writeback_22_bits_intWen_cons;
    extern constraint default_io_writeback_22_bits_fpWen_cons;
    extern constraint default_io_writeback_22_bits_exceptionVec_0_cons;
    extern constraint default_io_writeback_22_bits_exceptionVec_1_cons;
    extern constraint default_io_writeback_22_bits_exceptionVec_2_cons;
    extern constraint default_io_writeback_22_bits_exceptionVec_3_cons;
    extern constraint default_io_writeback_22_bits_exceptionVec_4_cons;
    extern constraint default_io_writeback_22_bits_exceptionVec_5_cons;
    extern constraint default_io_writeback_22_bits_exceptionVec_6_cons;
    extern constraint default_io_writeback_22_bits_exceptionVec_7_cons;
    extern constraint default_io_writeback_22_bits_exceptionVec_8_cons;
    extern constraint default_io_writeback_22_bits_exceptionVec_9_cons;
    extern constraint default_io_writeback_22_bits_exceptionVec_10_cons;
    extern constraint default_io_writeback_22_bits_exceptionVec_11_cons;
    extern constraint default_io_writeback_22_bits_exceptionVec_12_cons;
    extern constraint default_io_writeback_22_bits_exceptionVec_13_cons;
    extern constraint default_io_writeback_22_bits_exceptionVec_14_cons;
    extern constraint default_io_writeback_22_bits_exceptionVec_15_cons;
    extern constraint default_io_writeback_22_bits_exceptionVec_16_cons;
    extern constraint default_io_writeback_22_bits_exceptionVec_17_cons;
    extern constraint default_io_writeback_22_bits_exceptionVec_18_cons;
    extern constraint default_io_writeback_22_bits_exceptionVec_19_cons;
    extern constraint default_io_writeback_22_bits_exceptionVec_20_cons;
    extern constraint default_io_writeback_22_bits_exceptionVec_21_cons;
    extern constraint default_io_writeback_22_bits_exceptionVec_22_cons;
    extern constraint default_io_writeback_22_bits_exceptionVec_23_cons;
    extern constraint default_io_writeback_22_bits_flushPipe_cons;
    extern constraint default_io_writeback_22_bits_replay_cons;
    extern constraint default_io_writeback_22_bits_lqIdx_flag_cons;
    extern constraint default_io_writeback_22_bits_lqIdx_value_cons;
    extern constraint default_io_writeback_22_bits_trigger_cons;
    extern constraint default_io_writeback_22_bits_predecodeInfo_valid_cons;
    extern constraint default_io_writeback_22_bits_predecodeInfo_isRVC_cons;
    extern constraint default_io_writeback_22_bits_predecodeInfo_brType_cons;
    extern constraint default_io_writeback_22_bits_predecodeInfo_isCall_cons;
    extern constraint default_io_writeback_22_bits_predecodeInfo_isRet_cons;
    extern constraint default_io_writeback_22_bits_debug_isMMIO_cons;
    extern constraint default_io_writeback_22_bits_debug_isNCIO_cons;
    extern constraint default_io_writeback_22_bits_debug_isPerfCnt_cons;
    extern constraint default_io_writeback_22_bits_debug_paddr_cons;
    extern constraint default_io_writeback_22_bits_debug_vaddr_cons;
    extern constraint default_io_writeback_22_bits_debugInfo_eliminatedMove_cons;
    extern constraint default_io_writeback_22_bits_debugInfo_renameTime_cons;
    extern constraint default_io_writeback_22_bits_debugInfo_dispatchTime_cons;
    extern constraint default_io_writeback_22_bits_debugInfo_enqRsTime_cons;
    extern constraint default_io_writeback_22_bits_debugInfo_selectTime_cons;
    extern constraint default_io_writeback_22_bits_debugInfo_issueTime_cons;
    extern constraint default_io_writeback_22_bits_debugInfo_writebackTime_cons;
    extern constraint default_io_writeback_22_bits_debugInfo_runahead_checkpoint_id_cons;
    extern constraint default_io_writeback_22_bits_debugInfo_tlbFirstReqTime_cons;
    extern constraint default_io_writeback_22_bits_debugInfo_tlbRespTime_cons;
    extern constraint default_io_writeback_22_bits_debug_seqNum_cons;
    extern constraint default_io_writeback_21_valid_cons;
    extern constraint default_io_writeback_21_bits_data_0_cons;
    extern constraint default_io_writeback_21_bits_pdest_cons;
    extern constraint default_io_writeback_21_bits_robIdx_flag_cons;
    extern constraint default_io_writeback_21_bits_robIdx_value_cons;
    extern constraint default_io_writeback_21_bits_intWen_cons;
    extern constraint default_io_writeback_21_bits_fpWen_cons;
    extern constraint default_io_writeback_21_bits_exceptionVec_0_cons;
    extern constraint default_io_writeback_21_bits_exceptionVec_1_cons;
    extern constraint default_io_writeback_21_bits_exceptionVec_2_cons;
    extern constraint default_io_writeback_21_bits_exceptionVec_3_cons;
    extern constraint default_io_writeback_21_bits_exceptionVec_4_cons;
    extern constraint default_io_writeback_21_bits_exceptionVec_5_cons;
    extern constraint default_io_writeback_21_bits_exceptionVec_6_cons;
    extern constraint default_io_writeback_21_bits_exceptionVec_7_cons;
    extern constraint default_io_writeback_21_bits_exceptionVec_8_cons;
    extern constraint default_io_writeback_21_bits_exceptionVec_9_cons;
    extern constraint default_io_writeback_21_bits_exceptionVec_10_cons;
    extern constraint default_io_writeback_21_bits_exceptionVec_11_cons;
    extern constraint default_io_writeback_21_bits_exceptionVec_12_cons;
    extern constraint default_io_writeback_21_bits_exceptionVec_13_cons;
    extern constraint default_io_writeback_21_bits_exceptionVec_14_cons;
    extern constraint default_io_writeback_21_bits_exceptionVec_15_cons;
    extern constraint default_io_writeback_21_bits_exceptionVec_16_cons;
    extern constraint default_io_writeback_21_bits_exceptionVec_17_cons;
    extern constraint default_io_writeback_21_bits_exceptionVec_18_cons;
    extern constraint default_io_writeback_21_bits_exceptionVec_19_cons;
    extern constraint default_io_writeback_21_bits_exceptionVec_20_cons;
    extern constraint default_io_writeback_21_bits_exceptionVec_21_cons;
    extern constraint default_io_writeback_21_bits_exceptionVec_22_cons;
    extern constraint default_io_writeback_21_bits_exceptionVec_23_cons;
    extern constraint default_io_writeback_21_bits_flushPipe_cons;
    extern constraint default_io_writeback_21_bits_replay_cons;
    extern constraint default_io_writeback_21_bits_lqIdx_flag_cons;
    extern constraint default_io_writeback_21_bits_lqIdx_value_cons;
    extern constraint default_io_writeback_21_bits_trigger_cons;
    extern constraint default_io_writeback_21_bits_predecodeInfo_valid_cons;
    extern constraint default_io_writeback_21_bits_predecodeInfo_isRVC_cons;
    extern constraint default_io_writeback_21_bits_predecodeInfo_brType_cons;
    extern constraint default_io_writeback_21_bits_predecodeInfo_isCall_cons;
    extern constraint default_io_writeback_21_bits_predecodeInfo_isRet_cons;
    extern constraint default_io_writeback_21_bits_debug_isMMIO_cons;
    extern constraint default_io_writeback_21_bits_debug_isNCIO_cons;
    extern constraint default_io_writeback_21_bits_debug_isPerfCnt_cons;
    extern constraint default_io_writeback_21_bits_debug_paddr_cons;
    extern constraint default_io_writeback_21_bits_debug_vaddr_cons;
    extern constraint default_io_writeback_21_bits_debugInfo_eliminatedMove_cons;
    extern constraint default_io_writeback_21_bits_debugInfo_renameTime_cons;
    extern constraint default_io_writeback_21_bits_debugInfo_dispatchTime_cons;
    extern constraint default_io_writeback_21_bits_debugInfo_enqRsTime_cons;
    extern constraint default_io_writeback_21_bits_debugInfo_selectTime_cons;
    extern constraint default_io_writeback_21_bits_debugInfo_issueTime_cons;
    extern constraint default_io_writeback_21_bits_debugInfo_writebackTime_cons;
    extern constraint default_io_writeback_21_bits_debugInfo_runahead_checkpoint_id_cons;
    extern constraint default_io_writeback_21_bits_debugInfo_tlbFirstReqTime_cons;
    extern constraint default_io_writeback_21_bits_debugInfo_tlbRespTime_cons;
    extern constraint default_io_writeback_21_bits_debug_seqNum_cons;
    extern constraint default_io_writeback_20_valid_cons;
    extern constraint default_io_writeback_20_bits_data_0_cons;
    extern constraint default_io_writeback_20_bits_pdest_cons;
    extern constraint default_io_writeback_20_bits_robIdx_flag_cons;
    extern constraint default_io_writeback_20_bits_robIdx_value_cons;
    extern constraint default_io_writeback_20_bits_intWen_cons;
    extern constraint default_io_writeback_20_bits_fpWen_cons;
    extern constraint default_io_writeback_20_bits_exceptionVec_0_cons;
    extern constraint default_io_writeback_20_bits_exceptionVec_1_cons;
    extern constraint default_io_writeback_20_bits_exceptionVec_2_cons;
    extern constraint default_io_writeback_20_bits_exceptionVec_3_cons;
    extern constraint default_io_writeback_20_bits_exceptionVec_4_cons;
    extern constraint default_io_writeback_20_bits_exceptionVec_5_cons;
    extern constraint default_io_writeback_20_bits_exceptionVec_6_cons;
    extern constraint default_io_writeback_20_bits_exceptionVec_7_cons;
    extern constraint default_io_writeback_20_bits_exceptionVec_8_cons;
    extern constraint default_io_writeback_20_bits_exceptionVec_9_cons;
    extern constraint default_io_writeback_20_bits_exceptionVec_10_cons;
    extern constraint default_io_writeback_20_bits_exceptionVec_11_cons;
    extern constraint default_io_writeback_20_bits_exceptionVec_12_cons;
    extern constraint default_io_writeback_20_bits_exceptionVec_13_cons;
    extern constraint default_io_writeback_20_bits_exceptionVec_14_cons;
    extern constraint default_io_writeback_20_bits_exceptionVec_15_cons;
    extern constraint default_io_writeback_20_bits_exceptionVec_16_cons;
    extern constraint default_io_writeback_20_bits_exceptionVec_17_cons;
    extern constraint default_io_writeback_20_bits_exceptionVec_18_cons;
    extern constraint default_io_writeback_20_bits_exceptionVec_19_cons;
    extern constraint default_io_writeback_20_bits_exceptionVec_20_cons;
    extern constraint default_io_writeback_20_bits_exceptionVec_21_cons;
    extern constraint default_io_writeback_20_bits_exceptionVec_22_cons;
    extern constraint default_io_writeback_20_bits_exceptionVec_23_cons;
    extern constraint default_io_writeback_20_bits_flushPipe_cons;
    extern constraint default_io_writeback_20_bits_replay_cons;
    extern constraint default_io_writeback_20_bits_lqIdx_flag_cons;
    extern constraint default_io_writeback_20_bits_lqIdx_value_cons;
    extern constraint default_io_writeback_20_bits_trigger_cons;
    extern constraint default_io_writeback_20_bits_predecodeInfo_valid_cons;
    extern constraint default_io_writeback_20_bits_predecodeInfo_isRVC_cons;
    extern constraint default_io_writeback_20_bits_predecodeInfo_brType_cons;
    extern constraint default_io_writeback_20_bits_predecodeInfo_isCall_cons;
    extern constraint default_io_writeback_20_bits_predecodeInfo_isRet_cons;
    extern constraint default_io_writeback_20_bits_debug_isMMIO_cons;
    extern constraint default_io_writeback_20_bits_debug_isNCIO_cons;
    extern constraint default_io_writeback_20_bits_debug_isPerfCnt_cons;
    extern constraint default_io_writeback_20_bits_debug_paddr_cons;
    extern constraint default_io_writeback_20_bits_debug_vaddr_cons;
    extern constraint default_io_writeback_20_bits_debugInfo_eliminatedMove_cons;
    extern constraint default_io_writeback_20_bits_debugInfo_renameTime_cons;
    extern constraint default_io_writeback_20_bits_debugInfo_dispatchTime_cons;
    extern constraint default_io_writeback_20_bits_debugInfo_enqRsTime_cons;
    extern constraint default_io_writeback_20_bits_debugInfo_selectTime_cons;
    extern constraint default_io_writeback_20_bits_debugInfo_issueTime_cons;
    extern constraint default_io_writeback_20_bits_debugInfo_writebackTime_cons;
    extern constraint default_io_writeback_20_bits_debugInfo_runahead_checkpoint_id_cons;
    extern constraint default_io_writeback_20_bits_debugInfo_tlbFirstReqTime_cons;
    extern constraint default_io_writeback_20_bits_debugInfo_tlbRespTime_cons;
    extern constraint default_io_writeback_20_bits_debug_seqNum_cons;
    extern constraint default_io_writeback_19_valid_cons;
    extern constraint default_io_writeback_19_bits_data_0_cons;
    extern constraint default_io_writeback_19_bits_pdest_cons;
    extern constraint default_io_writeback_19_bits_robIdx_flag_cons;
    extern constraint default_io_writeback_19_bits_robIdx_value_cons;
    extern constraint default_io_writeback_19_bits_intWen_cons;
    extern constraint default_io_writeback_19_bits_exceptionVec_0_cons;
    extern constraint default_io_writeback_19_bits_exceptionVec_1_cons;
    extern constraint default_io_writeback_19_bits_exceptionVec_2_cons;
    extern constraint default_io_writeback_19_bits_exceptionVec_3_cons;
    extern constraint default_io_writeback_19_bits_exceptionVec_4_cons;
    extern constraint default_io_writeback_19_bits_exceptionVec_5_cons;
    extern constraint default_io_writeback_19_bits_exceptionVec_6_cons;
    extern constraint default_io_writeback_19_bits_exceptionVec_7_cons;
    extern constraint default_io_writeback_19_bits_exceptionVec_8_cons;
    extern constraint default_io_writeback_19_bits_exceptionVec_9_cons;
    extern constraint default_io_writeback_19_bits_exceptionVec_10_cons;
    extern constraint default_io_writeback_19_bits_exceptionVec_11_cons;
    extern constraint default_io_writeback_19_bits_exceptionVec_12_cons;
    extern constraint default_io_writeback_19_bits_exceptionVec_13_cons;
    extern constraint default_io_writeback_19_bits_exceptionVec_14_cons;
    extern constraint default_io_writeback_19_bits_exceptionVec_15_cons;
    extern constraint default_io_writeback_19_bits_exceptionVec_16_cons;
    extern constraint default_io_writeback_19_bits_exceptionVec_17_cons;
    extern constraint default_io_writeback_19_bits_exceptionVec_18_cons;
    extern constraint default_io_writeback_19_bits_exceptionVec_19_cons;
    extern constraint default_io_writeback_19_bits_exceptionVec_20_cons;
    extern constraint default_io_writeback_19_bits_exceptionVec_21_cons;
    extern constraint default_io_writeback_19_bits_exceptionVec_22_cons;
    extern constraint default_io_writeback_19_bits_exceptionVec_23_cons;
    extern constraint default_io_writeback_19_bits_flushPipe_cons;
    extern constraint default_io_writeback_19_bits_sqIdx_flag_cons;
    extern constraint default_io_writeback_19_bits_sqIdx_value_cons;
    extern constraint default_io_writeback_19_bits_trigger_cons;
    extern constraint default_io_writeback_19_bits_debug_isMMIO_cons;
    extern constraint default_io_writeback_19_bits_debug_isNCIO_cons;
    extern constraint default_io_writeback_19_bits_debug_isPerfCnt_cons;
    extern constraint default_io_writeback_19_bits_debug_paddr_cons;
    extern constraint default_io_writeback_19_bits_debug_vaddr_cons;
    extern constraint default_io_writeback_19_bits_debugInfo_eliminatedMove_cons;
    extern constraint default_io_writeback_19_bits_debugInfo_renameTime_cons;
    extern constraint default_io_writeback_19_bits_debugInfo_dispatchTime_cons;
    extern constraint default_io_writeback_19_bits_debugInfo_enqRsTime_cons;
    extern constraint default_io_writeback_19_bits_debugInfo_selectTime_cons;
    extern constraint default_io_writeback_19_bits_debugInfo_issueTime_cons;
    extern constraint default_io_writeback_19_bits_debugInfo_writebackTime_cons;
    extern constraint default_io_writeback_19_bits_debugInfo_runahead_checkpoint_id_cons;
    extern constraint default_io_writeback_19_bits_debugInfo_tlbFirstReqTime_cons;
    extern constraint default_io_writeback_19_bits_debugInfo_tlbRespTime_cons;
    extern constraint default_io_writeback_19_bits_debug_seqNum_cons;
    extern constraint default_io_writeback_18_valid_cons;
    extern constraint default_io_writeback_18_bits_data_0_cons;
    extern constraint default_io_writeback_18_bits_pdest_cons;
    extern constraint default_io_writeback_18_bits_robIdx_flag_cons;
    extern constraint default_io_writeback_18_bits_robIdx_value_cons;
    extern constraint default_io_writeback_18_bits_intWen_cons;
    extern constraint default_io_writeback_18_bits_exceptionVec_0_cons;
    extern constraint default_io_writeback_18_bits_exceptionVec_1_cons;
    extern constraint default_io_writeback_18_bits_exceptionVec_2_cons;
    extern constraint default_io_writeback_18_bits_exceptionVec_3_cons;
    extern constraint default_io_writeback_18_bits_exceptionVec_4_cons;
    extern constraint default_io_writeback_18_bits_exceptionVec_5_cons;
    extern constraint default_io_writeback_18_bits_exceptionVec_6_cons;
    extern constraint default_io_writeback_18_bits_exceptionVec_7_cons;
    extern constraint default_io_writeback_18_bits_exceptionVec_8_cons;
    extern constraint default_io_writeback_18_bits_exceptionVec_9_cons;
    extern constraint default_io_writeback_18_bits_exceptionVec_10_cons;
    extern constraint default_io_writeback_18_bits_exceptionVec_11_cons;
    extern constraint default_io_writeback_18_bits_exceptionVec_12_cons;
    extern constraint default_io_writeback_18_bits_exceptionVec_13_cons;
    extern constraint default_io_writeback_18_bits_exceptionVec_14_cons;
    extern constraint default_io_writeback_18_bits_exceptionVec_15_cons;
    extern constraint default_io_writeback_18_bits_exceptionVec_16_cons;
    extern constraint default_io_writeback_18_bits_exceptionVec_17_cons;
    extern constraint default_io_writeback_18_bits_exceptionVec_18_cons;
    extern constraint default_io_writeback_18_bits_exceptionVec_19_cons;
    extern constraint default_io_writeback_18_bits_exceptionVec_20_cons;
    extern constraint default_io_writeback_18_bits_exceptionVec_21_cons;
    extern constraint default_io_writeback_18_bits_exceptionVec_22_cons;
    extern constraint default_io_writeback_18_bits_exceptionVec_23_cons;
    extern constraint default_io_writeback_18_bits_flushPipe_cons;
    extern constraint default_io_writeback_18_bits_sqIdx_flag_cons;
    extern constraint default_io_writeback_18_bits_sqIdx_value_cons;
    extern constraint default_io_writeback_18_bits_trigger_cons;
    extern constraint default_io_writeback_18_bits_debug_isMMIO_cons;
    extern constraint default_io_writeback_18_bits_debug_isNCIO_cons;
    extern constraint default_io_writeback_18_bits_debug_isPerfCnt_cons;
    extern constraint default_io_writeback_18_bits_debug_paddr_cons;
    extern constraint default_io_writeback_18_bits_debug_vaddr_cons;
    extern constraint default_io_writeback_18_bits_debugInfo_eliminatedMove_cons;
    extern constraint default_io_writeback_18_bits_debugInfo_renameTime_cons;
    extern constraint default_io_writeback_18_bits_debugInfo_dispatchTime_cons;
    extern constraint default_io_writeback_18_bits_debugInfo_enqRsTime_cons;
    extern constraint default_io_writeback_18_bits_debugInfo_selectTime_cons;
    extern constraint default_io_writeback_18_bits_debugInfo_issueTime_cons;
    extern constraint default_io_writeback_18_bits_debugInfo_writebackTime_cons;
    extern constraint default_io_writeback_18_bits_debugInfo_runahead_checkpoint_id_cons;
    extern constraint default_io_writeback_18_bits_debugInfo_tlbFirstReqTime_cons;
    extern constraint default_io_writeback_18_bits_debugInfo_tlbRespTime_cons;
    extern constraint default_io_writeback_18_bits_debug_seqNum_cons;
    extern constraint default_io_writeback_17_valid_cons;
    extern constraint default_io_writeback_17_bits_data_0_cons;
    extern constraint default_io_writeback_17_bits_data_1_cons;
    extern constraint default_io_writeback_17_bits_data_2_cons;
    extern constraint default_io_writeback_17_bits_pdest_cons;
    extern constraint default_io_writeback_17_bits_robIdx_flag_cons;
    extern constraint default_io_writeback_17_bits_robIdx_value_cons;
    extern constraint default_io_writeback_17_bits_vecWen_cons;
    extern constraint default_io_writeback_17_bits_v0Wen_cons;
    extern constraint default_io_writeback_17_bits_fflags_cons;
    extern constraint default_io_writeback_17_bits_wflags_cons;
    extern constraint default_io_writeback_17_bits_debugInfo_eliminatedMove_cons;
    extern constraint default_io_writeback_17_bits_debugInfo_renameTime_cons;
    extern constraint default_io_writeback_17_bits_debugInfo_dispatchTime_cons;
    extern constraint default_io_writeback_17_bits_debugInfo_enqRsTime_cons;
    extern constraint default_io_writeback_17_bits_debugInfo_selectTime_cons;
    extern constraint default_io_writeback_17_bits_debugInfo_issueTime_cons;
    extern constraint default_io_writeback_17_bits_debugInfo_writebackTime_cons;
    extern constraint default_io_writeback_17_bits_debugInfo_runahead_checkpoint_id_cons;
    extern constraint default_io_writeback_17_bits_debugInfo_tlbFirstReqTime_cons;
    extern constraint default_io_writeback_17_bits_debugInfo_tlbRespTime_cons;
    extern constraint default_io_writeback_17_bits_debug_seqNum_cons;
    extern constraint default_io_writeback_16_valid_cons;
    extern constraint default_io_writeback_16_bits_data_0_cons;
    extern constraint default_io_writeback_16_bits_data_1_cons;
    extern constraint default_io_writeback_16_bits_data_2_cons;
    extern constraint default_io_writeback_16_bits_data_3_cons;
    extern constraint default_io_writeback_16_bits_pdest_cons;
    extern constraint default_io_writeback_16_bits_robIdx_flag_cons;
    extern constraint default_io_writeback_16_bits_robIdx_value_cons;
    extern constraint default_io_writeback_16_bits_fpWen_cons;
    extern constraint default_io_writeback_16_bits_vecWen_cons;
    extern constraint default_io_writeback_16_bits_v0Wen_cons;
    extern constraint default_io_writeback_16_bits_fflags_cons;
    extern constraint default_io_writeback_16_bits_wflags_cons;
    extern constraint default_io_writeback_16_bits_debugInfo_eliminatedMove_cons;
    extern constraint default_io_writeback_16_bits_debugInfo_renameTime_cons;
    extern constraint default_io_writeback_16_bits_debugInfo_dispatchTime_cons;
    extern constraint default_io_writeback_16_bits_debugInfo_enqRsTime_cons;
    extern constraint default_io_writeback_16_bits_debugInfo_selectTime_cons;
    extern constraint default_io_writeback_16_bits_debugInfo_issueTime_cons;
    extern constraint default_io_writeback_16_bits_debugInfo_writebackTime_cons;
    extern constraint default_io_writeback_16_bits_debugInfo_runahead_checkpoint_id_cons;
    extern constraint default_io_writeback_16_bits_debugInfo_tlbFirstReqTime_cons;
    extern constraint default_io_writeback_16_bits_debugInfo_tlbRespTime_cons;
    extern constraint default_io_writeback_16_bits_debug_seqNum_cons;
    extern constraint default_io_writeback_15_valid_cons;
    extern constraint default_io_writeback_15_bits_data_0_cons;
    extern constraint default_io_writeback_15_bits_data_1_cons;
    extern constraint default_io_writeback_15_bits_data_2_cons;
    extern constraint default_io_writeback_15_bits_pdest_cons;
    extern constraint default_io_writeback_15_bits_robIdx_flag_cons;
    extern constraint default_io_writeback_15_bits_robIdx_value_cons;
    extern constraint default_io_writeback_15_bits_vecWen_cons;
    extern constraint default_io_writeback_15_bits_v0Wen_cons;
    extern constraint default_io_writeback_15_bits_fflags_cons;
    extern constraint default_io_writeback_15_bits_wflags_cons;
    extern constraint default_io_writeback_15_bits_vxsat_cons;
    extern constraint default_io_writeback_15_bits_debugInfo_eliminatedMove_cons;
    extern constraint default_io_writeback_15_bits_debugInfo_renameTime_cons;
    extern constraint default_io_writeback_15_bits_debugInfo_dispatchTime_cons;
    extern constraint default_io_writeback_15_bits_debugInfo_enqRsTime_cons;
    extern constraint default_io_writeback_15_bits_debugInfo_selectTime_cons;
    extern constraint default_io_writeback_15_bits_debugInfo_issueTime_cons;
    extern constraint default_io_writeback_15_bits_debugInfo_writebackTime_cons;
    extern constraint default_io_writeback_15_bits_debugInfo_runahead_checkpoint_id_cons;
    extern constraint default_io_writeback_15_bits_debugInfo_tlbFirstReqTime_cons;
    extern constraint default_io_writeback_15_bits_debugInfo_tlbRespTime_cons;
    extern constraint default_io_writeback_15_bits_debug_seqNum_cons;
    extern constraint default_io_writeback_14_valid_cons;
    extern constraint default_io_writeback_14_bits_data_0_cons;
    extern constraint default_io_writeback_14_bits_data_1_cons;
    extern constraint default_io_writeback_14_bits_data_2_cons;
    extern constraint default_io_writeback_14_bits_data_3_cons;
    extern constraint default_io_writeback_14_bits_data_4_cons;
    extern constraint default_io_writeback_14_bits_data_5_cons;
    extern constraint default_io_writeback_14_bits_pdest_cons;
    extern constraint default_io_writeback_14_bits_robIdx_flag_cons;
    extern constraint default_io_writeback_14_bits_robIdx_value_cons;
    extern constraint default_io_writeback_14_bits_intWen_cons;
    extern constraint default_io_writeback_14_bits_fpWen_cons;
    extern constraint default_io_writeback_14_bits_vecWen_cons;
    extern constraint default_io_writeback_14_bits_v0Wen_cons;
    extern constraint default_io_writeback_14_bits_vlWen_cons;
    extern constraint default_io_writeback_14_bits_fflags_cons;
    extern constraint default_io_writeback_14_bits_wflags_cons;
    extern constraint default_io_writeback_14_bits_exceptionVec_2_cons;
    extern constraint default_io_writeback_14_bits_debugInfo_eliminatedMove_cons;
    extern constraint default_io_writeback_14_bits_debugInfo_renameTime_cons;
    extern constraint default_io_writeback_14_bits_debugInfo_dispatchTime_cons;
    extern constraint default_io_writeback_14_bits_debugInfo_enqRsTime_cons;
    extern constraint default_io_writeback_14_bits_debugInfo_selectTime_cons;
    extern constraint default_io_writeback_14_bits_debugInfo_issueTime_cons;
    extern constraint default_io_writeback_14_bits_debugInfo_writebackTime_cons;
    extern constraint default_io_writeback_14_bits_debugInfo_runahead_checkpoint_id_cons;
    extern constraint default_io_writeback_14_bits_debugInfo_tlbFirstReqTime_cons;
    extern constraint default_io_writeback_14_bits_debugInfo_tlbRespTime_cons;
    extern constraint default_io_writeback_14_bits_debug_seqNum_cons;
    extern constraint default_io_writeback_13_valid_cons;
    extern constraint default_io_writeback_13_bits_data_0_cons;
    extern constraint default_io_writeback_13_bits_data_1_cons;
    extern constraint default_io_writeback_13_bits_data_2_cons;
    extern constraint default_io_writeback_13_bits_pdest_cons;
    extern constraint default_io_writeback_13_bits_robIdx_flag_cons;
    extern constraint default_io_writeback_13_bits_robIdx_value_cons;
    extern constraint default_io_writeback_13_bits_vecWen_cons;
    extern constraint default_io_writeback_13_bits_v0Wen_cons;
    extern constraint default_io_writeback_13_bits_fflags_cons;
    extern constraint default_io_writeback_13_bits_wflags_cons;
    extern constraint default_io_writeback_13_bits_vxsat_cons;
    extern constraint default_io_writeback_13_bits_exceptionVec_2_cons;
    extern constraint default_io_writeback_13_bits_debugInfo_eliminatedMove_cons;
    extern constraint default_io_writeback_13_bits_debugInfo_renameTime_cons;
    extern constraint default_io_writeback_13_bits_debugInfo_dispatchTime_cons;
    extern constraint default_io_writeback_13_bits_debugInfo_enqRsTime_cons;
    extern constraint default_io_writeback_13_bits_debugInfo_selectTime_cons;
    extern constraint default_io_writeback_13_bits_debugInfo_issueTime_cons;
    extern constraint default_io_writeback_13_bits_debugInfo_writebackTime_cons;
    extern constraint default_io_writeback_13_bits_debugInfo_runahead_checkpoint_id_cons;
    extern constraint default_io_writeback_13_bits_debugInfo_tlbFirstReqTime_cons;
    extern constraint default_io_writeback_13_bits_debugInfo_tlbRespTime_cons;
    extern constraint default_io_writeback_13_bits_debug_seqNum_cons;
    extern constraint default_io_writeback_7_valid_cons;
    extern constraint default_io_writeback_7_bits_data_0_cons;
    extern constraint default_io_writeback_7_bits_data_1_cons;
    extern constraint default_io_writeback_7_bits_pdest_cons;
    extern constraint default_io_writeback_7_bits_robIdx_flag_cons;
    extern constraint default_io_writeback_7_bits_robIdx_value_cons;
    extern constraint default_io_writeback_7_bits_intWen_cons;
    extern constraint default_io_writeback_7_bits_redirect_valid_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_isRVC_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_robIdx_flag_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_robIdx_value_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_ftqIdx_flag_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_ftqIdx_value_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_ftqOffset_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_level_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_interrupt_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_pc_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_ssp_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_sctr_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_ghr_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_target_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_taken_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_shift_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_fullTarget_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_stFtqIdx_flag_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_stFtqIdx_value_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_stFtqOffset_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_debugIsCtrl_cons;
    extern constraint default_io_writeback_7_bits_redirect_bits_debugIsMemVio_cons;
    extern constraint default_io_writeback_7_bits_exceptionVec_2_cons;
    extern constraint default_io_writeback_7_bits_exceptionVec_3_cons;
    extern constraint default_io_writeback_7_bits_exceptionVec_8_cons;
    extern constraint default_io_writeback_7_bits_exceptionVec_9_cons;
    extern constraint default_io_writeback_7_bits_exceptionVec_10_cons;
    extern constraint default_io_writeback_7_bits_exceptionVec_11_cons;
    extern constraint default_io_writeback_7_bits_exceptionVec_22_cons;
    extern constraint default_io_writeback_7_bits_flushPipe_cons;
    extern constraint default_io_writeback_7_bits_predecodeInfo_valid_cons;
    extern constraint default_io_writeback_7_bits_predecodeInfo_isRVC_cons;
    extern constraint default_io_writeback_7_bits_predecodeInfo_brType_cons;
    extern constraint default_io_writeback_7_bits_predecodeInfo_isCall_cons;
    extern constraint default_io_writeback_7_bits_predecodeInfo_isRet_cons;
    extern constraint default_io_writeback_7_bits_debug_isPerfCnt_cons;
    extern constraint default_io_writeback_7_bits_debugInfo_eliminatedMove_cons;
    extern constraint default_io_writeback_7_bits_debugInfo_renameTime_cons;
    extern constraint default_io_writeback_7_bits_debugInfo_dispatchTime_cons;
    extern constraint default_io_writeback_7_bits_debugInfo_enqRsTime_cons;
    extern constraint default_io_writeback_7_bits_debugInfo_selectTime_cons;
    extern constraint default_io_writeback_7_bits_debugInfo_issueTime_cons;
    extern constraint default_io_writeback_7_bits_debugInfo_writebackTime_cons;
    extern constraint default_io_writeback_7_bits_debugInfo_runahead_checkpoint_id_cons;
    extern constraint default_io_writeback_7_bits_debugInfo_tlbFirstReqTime_cons;
    extern constraint default_io_writeback_7_bits_debugInfo_tlbRespTime_cons;
    extern constraint default_io_writeback_7_bits_debug_seqNum_cons;
    extern constraint default_io_writeback_5_valid_cons;
    extern constraint default_io_writeback_5_bits_redirect_valid_cons;
    extern constraint default_io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred_cons;
    extern constraint default_io_writeback_3_valid_cons;
    extern constraint default_io_writeback_3_bits_redirect_valid_cons;
    extern constraint default_io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred_cons;
    extern constraint default_io_writeback_1_valid_cons;
    extern constraint default_io_writeback_1_bits_redirect_valid_cons;
    extern constraint default_io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred_cons;
    extern constraint default_io_exuWriteback_26_valid_cons;
    extern constraint default_io_exuWriteback_26_bits_robIdx_value_cons;
    extern constraint default_io_exuWriteback_25_valid_cons;
    extern constraint default_io_exuWriteback_25_bits_robIdx_value_cons;
    extern constraint default_io_exuWriteback_24_valid_cons;
    extern constraint default_io_exuWriteback_24_bits_data_0_cons;
    extern constraint default_io_exuWriteback_24_bits_pdest_cons;
    extern constraint default_io_exuWriteback_24_bits_robIdx_value_cons;
    extern constraint default_io_exuWriteback_24_bits_vecWen_cons;
    extern constraint default_io_exuWriteback_24_bits_v0Wen_cons;
    extern constraint default_io_exuWriteback_24_bits_vls_vdIdx_cons;
    extern constraint default_io_exuWriteback_24_bits_debug_isMMIO_cons;
    extern constraint default_io_exuWriteback_24_bits_debug_isNCIO_cons;
    extern constraint default_io_exuWriteback_24_bits_debug_isPerfCnt_cons;
    extern constraint default_io_exuWriteback_24_bits_debug_paddr_cons;
    extern constraint default_io_exuWriteback_23_valid_cons;
    extern constraint default_io_exuWriteback_23_bits_data_0_cons;
    extern constraint default_io_exuWriteback_23_bits_pdest_cons;
    extern constraint default_io_exuWriteback_23_bits_robIdx_value_cons;
    extern constraint default_io_exuWriteback_23_bits_vecWen_cons;
    extern constraint default_io_exuWriteback_23_bits_v0Wen_cons;
    extern constraint default_io_exuWriteback_23_bits_vls_vdIdx_cons;
    extern constraint default_io_exuWriteback_23_bits_debug_isMMIO_cons;
    extern constraint default_io_exuWriteback_23_bits_debug_isNCIO_cons;
    extern constraint default_io_exuWriteback_23_bits_debug_isPerfCnt_cons;
    extern constraint default_io_exuWriteback_23_bits_debug_paddr_cons;
    extern constraint default_io_exuWriteback_22_valid_cons;
    extern constraint default_io_exuWriteback_22_bits_data_0_cons;
    extern constraint default_io_exuWriteback_22_bits_robIdx_value_cons;
    extern constraint default_io_exuWriteback_22_bits_lqIdx_value_cons;
    extern constraint default_io_exuWriteback_22_bits_debug_isMMIO_cons;
    extern constraint default_io_exuWriteback_22_bits_debug_isNCIO_cons;
    extern constraint default_io_exuWriteback_22_bits_debug_isPerfCnt_cons;
    extern constraint default_io_exuWriteback_22_bits_debug_paddr_cons;
    extern constraint default_io_exuWriteback_21_valid_cons;
    extern constraint default_io_exuWriteback_21_bits_data_0_cons;
    extern constraint default_io_exuWriteback_21_bits_robIdx_value_cons;
    extern constraint default_io_exuWriteback_21_bits_lqIdx_value_cons;
    extern constraint default_io_exuWriteback_21_bits_debug_isMMIO_cons;
    extern constraint default_io_exuWriteback_21_bits_debug_isNCIO_cons;
    extern constraint default_io_exuWriteback_21_bits_debug_isPerfCnt_cons;
    extern constraint default_io_exuWriteback_21_bits_debug_paddr_cons;
    extern constraint default_io_exuWriteback_20_valid_cons;
    extern constraint default_io_exuWriteback_20_bits_data_0_cons;
    extern constraint default_io_exuWriteback_20_bits_robIdx_value_cons;
    extern constraint default_io_exuWriteback_20_bits_lqIdx_value_cons;
    extern constraint default_io_exuWriteback_20_bits_debug_isMMIO_cons;
    extern constraint default_io_exuWriteback_20_bits_debug_isNCIO_cons;
    extern constraint default_io_exuWriteback_20_bits_debug_isPerfCnt_cons;
    extern constraint default_io_exuWriteback_20_bits_debug_paddr_cons;
    extern constraint default_io_exuWriteback_19_valid_cons;
    extern constraint default_io_exuWriteback_19_bits_data_0_cons;
    extern constraint default_io_exuWriteback_19_bits_robIdx_value_cons;
    extern constraint default_io_exuWriteback_19_bits_sqIdx_value_cons;
    extern constraint default_io_exuWriteback_19_bits_debug_isMMIO_cons;
    extern constraint default_io_exuWriteback_19_bits_debug_isNCIO_cons;
    extern constraint default_io_exuWriteback_19_bits_debug_isPerfCnt_cons;
    extern constraint default_io_exuWriteback_19_bits_debug_paddr_cons;
    extern constraint default_io_exuWriteback_18_valid_cons;
    extern constraint default_io_exuWriteback_18_bits_data_0_cons;
    extern constraint default_io_exuWriteback_18_bits_robIdx_value_cons;
    extern constraint default_io_exuWriteback_18_bits_sqIdx_value_cons;
    extern constraint default_io_exuWriteback_18_bits_debug_isMMIO_cons;
    extern constraint default_io_exuWriteback_18_bits_debug_isNCIO_cons;
    extern constraint default_io_exuWriteback_18_bits_debug_isPerfCnt_cons;
    extern constraint default_io_exuWriteback_18_bits_debug_paddr_cons;
    extern constraint default_io_exuWriteback_17_valid_cons;
    extern constraint default_io_exuWriteback_17_bits_data_0_cons;
    extern constraint default_io_exuWriteback_17_bits_robIdx_value_cons;
    extern constraint default_io_exuWriteback_17_bits_fflags_cons;
    extern constraint default_io_exuWriteback_17_bits_wflags_cons;
    extern constraint default_io_exuWriteback_16_valid_cons;
    extern constraint default_io_exuWriteback_16_bits_data_0_cons;
    extern constraint default_io_exuWriteback_16_bits_robIdx_value_cons;
    extern constraint default_io_exuWriteback_16_bits_fflags_cons;
    extern constraint default_io_exuWriteback_16_bits_wflags_cons;
    extern constraint default_io_exuWriteback_15_valid_cons;
    extern constraint default_io_exuWriteback_15_bits_data_0_cons;
    extern constraint default_io_exuWriteback_15_bits_robIdx_value_cons;
    extern constraint default_io_exuWriteback_15_bits_fflags_cons;
    extern constraint default_io_exuWriteback_15_bits_wflags_cons;
    extern constraint default_io_exuWriteback_15_bits_vxsat_cons;
    extern constraint default_io_exuWriteback_14_valid_cons;
    extern constraint default_io_exuWriteback_14_bits_data_0_cons;
    extern constraint default_io_exuWriteback_14_bits_robIdx_value_cons;
    extern constraint default_io_exuWriteback_14_bits_fflags_cons;
    extern constraint default_io_exuWriteback_14_bits_wflags_cons;
    extern constraint default_io_exuWriteback_13_valid_cons;
    extern constraint default_io_exuWriteback_13_bits_data_0_cons;
    extern constraint default_io_exuWriteback_13_bits_robIdx_value_cons;
    extern constraint default_io_exuWriteback_13_bits_fflags_cons;
    extern constraint default_io_exuWriteback_13_bits_wflags_cons;
    extern constraint default_io_exuWriteback_13_bits_vxsat_cons;
    extern constraint default_io_exuWriteback_12_valid_cons;
    extern constraint default_io_exuWriteback_12_bits_data_0_cons;
    extern constraint default_io_exuWriteback_12_bits_robIdx_value_cons;
    extern constraint default_io_exuWriteback_12_bits_fflags_cons;
    extern constraint default_io_exuWriteback_12_bits_wflags_cons;
    extern constraint default_io_exuWriteback_11_valid_cons;
    extern constraint default_io_exuWriteback_11_bits_data_0_cons;
    extern constraint default_io_exuWriteback_11_bits_robIdx_value_cons;
    extern constraint default_io_exuWriteback_11_bits_fflags_cons;
    extern constraint default_io_exuWriteback_11_bits_wflags_cons;
    extern constraint default_io_exuWriteback_10_valid_cons;
    extern constraint default_io_exuWriteback_10_bits_data_0_cons;
    extern constraint default_io_exuWriteback_10_bits_robIdx_value_cons;
    extern constraint default_io_exuWriteback_10_bits_fflags_cons;
    extern constraint default_io_exuWriteback_10_bits_wflags_cons;
    extern constraint default_io_exuWriteback_9_valid_cons;
    extern constraint default_io_exuWriteback_9_bits_data_0_cons;
    extern constraint default_io_exuWriteback_9_bits_robIdx_value_cons;
    extern constraint default_io_exuWriteback_9_bits_fflags_cons;
    extern constraint default_io_exuWriteback_9_bits_wflags_cons;
    extern constraint default_io_exuWriteback_8_valid_cons;
    extern constraint default_io_exuWriteback_8_bits_data_0_cons;
    extern constraint default_io_exuWriteback_8_bits_robIdx_value_cons;
    extern constraint default_io_exuWriteback_8_bits_fflags_cons;
    extern constraint default_io_exuWriteback_8_bits_wflags_cons;
    extern constraint default_io_exuWriteback_7_valid_cons;
    extern constraint default_io_exuWriteback_7_bits_data_0_cons;
    extern constraint default_io_exuWriteback_7_bits_robIdx_value_cons;
    extern constraint default_io_exuWriteback_7_bits_debug_isPerfCnt_cons;
    extern constraint default_io_exuWriteback_6_valid_cons;
    extern constraint default_io_exuWriteback_6_bits_data_0_cons;
    extern constraint default_io_exuWriteback_6_bits_robIdx_value_cons;
    extern constraint default_io_exuWriteback_5_valid_cons;
    extern constraint default_io_exuWriteback_5_bits_data_0_cons;
    extern constraint default_io_exuWriteback_5_bits_robIdx_value_cons;
    extern constraint default_io_exuWriteback_5_bits_redirect_valid_cons;
    extern constraint default_io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken_cons;
    extern constraint default_io_exuWriteback_5_bits_fflags_cons;
    extern constraint default_io_exuWriteback_5_bits_wflags_cons;
    extern constraint default_io_exuWriteback_4_valid_cons;
    extern constraint default_io_exuWriteback_4_bits_data_0_cons;
    extern constraint default_io_exuWriteback_4_bits_robIdx_value_cons;
    extern constraint default_io_exuWriteback_3_valid_cons;
    extern constraint default_io_exuWriteback_3_bits_data_0_cons;
    extern constraint default_io_exuWriteback_3_bits_robIdx_value_cons;
    extern constraint default_io_exuWriteback_3_bits_redirect_valid_cons;
    extern constraint default_io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken_cons;
    extern constraint default_io_exuWriteback_2_valid_cons;
    extern constraint default_io_exuWriteback_2_bits_data_0_cons;
    extern constraint default_io_exuWriteback_2_bits_robIdx_value_cons;
    extern constraint default_io_exuWriteback_1_valid_cons;
    extern constraint default_io_exuWriteback_1_bits_data_0_cons;
    extern constraint default_io_exuWriteback_1_bits_robIdx_value_cons;
    extern constraint default_io_exuWriteback_1_bits_redirect_valid_cons;
    extern constraint default_io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken_cons;
    extern constraint default_io_exuWriteback_0_valid_cons;
    extern constraint default_io_exuWriteback_0_bits_data_0_cons;
    extern constraint default_io_exuWriteback_0_bits_robIdx_value_cons;
    extern constraint default_io_writebackNums_0_bits_cons;
    extern constraint default_io_writebackNums_1_bits_cons;
    extern constraint default_io_writebackNums_2_bits_cons;
    extern constraint default_io_writebackNums_3_bits_cons;
    extern constraint default_io_writebackNums_4_bits_cons;
    extern constraint default_io_writebackNums_5_bits_cons;
    extern constraint default_io_writebackNums_6_bits_cons;
    extern constraint default_io_writebackNums_7_bits_cons;
    extern constraint default_io_writebackNums_8_bits_cons;
    extern constraint default_io_writebackNums_9_bits_cons;
    extern constraint default_io_writebackNums_10_bits_cons;
    extern constraint default_io_writebackNums_11_bits_cons;
    extern constraint default_io_writebackNums_12_bits_cons;
    extern constraint default_io_writebackNums_13_bits_cons;
    extern constraint default_io_writebackNums_14_bits_cons;
    extern constraint default_io_writebackNums_15_bits_cons;
    extern constraint default_io_writebackNums_16_bits_cons;
    extern constraint default_io_writebackNums_17_bits_cons;
    extern constraint default_io_writebackNums_18_bits_cons;
    extern constraint default_io_writebackNums_19_bits_cons;
    extern constraint default_io_writebackNums_20_bits_cons;
    extern constraint default_io_writebackNums_21_bits_cons;
    extern constraint default_io_writebackNums_22_bits_cons;
    extern constraint default_io_writebackNums_23_bits_cons;
    extern constraint default_io_writebackNums_24_bits_cons;
    extern constraint default_io_writebackNeedFlush_0_cons;
    extern constraint default_io_writebackNeedFlush_1_cons;
    extern constraint default_io_writebackNeedFlush_2_cons;
    extern constraint default_io_writebackNeedFlush_6_cons;
    extern constraint default_io_writebackNeedFlush_7_cons;
    extern constraint default_io_writebackNeedFlush_8_cons;
    extern constraint default_io_writebackNeedFlush_9_cons;
    extern constraint default_io_writebackNeedFlush_10_cons;
    extern constraint default_io_writebackNeedFlush_11_cons;
    extern constraint default_io_writebackNeedFlush_12_cons;

    extern function new(string name="WriteBack_in_agent_xaction");
    extern function void pack();
    extern function void unpack();
    extern function void pre_randomize();
    extern function void post_randomize();
    extern function string psdisplay(string prefix = "");
    extern function bit compare(uvm_object rhs, uvm_comparer comparer=null);

    `uvm_object_utils_begin(WriteBack_in_agent_xaction)
        `uvm_field_int(io_writeback_24_valid, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_pdest, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_robIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_exceptionVec_0, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_exceptionVec_1, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_exceptionVec_2, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_exceptionVec_3, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_exceptionVec_4, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_exceptionVec_5, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_exceptionVec_6, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_exceptionVec_7, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_exceptionVec_8, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_exceptionVec_9, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_exceptionVec_10, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_exceptionVec_11, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_exceptionVec_12, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_exceptionVec_13, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_exceptionVec_14, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_exceptionVec_15, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_exceptionVec_16, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_exceptionVec_17, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_exceptionVec_18, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_exceptionVec_19, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_exceptionVec_20, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_exceptionVec_21, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_exceptionVec_22, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_exceptionVec_23, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_flushPipe, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_replay, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_trigger, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_vill, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_vma, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_vta, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_vsew, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_vlmul, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_specVill, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_specVma, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_specVta, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_specVsew, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_specVlmul, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_vm, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_vstart, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_frm, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_fpu_isFP32Instr, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_fpu_isFP64Instr, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_fpu_isReduction, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_vxrm, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_vuopIdx, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_lastUop, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_vmask, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_vl, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_nf, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_veew, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_isReverse, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_isExt, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_isNarrow, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_isDstMask, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_isOpMask, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_isMove, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_isDependOldVd, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_isWritePartVd, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vpu_isVleff, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_oldVdPsrc, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vdIdx, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_vdIdxInField, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_isIndexed, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_isMasked, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_isStrided, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_isWhole, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_isVecLoad, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_vls_isVlm, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_debug_isMMIO, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_debug_isNCIO, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_debug_isPerfCnt, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_debug_paddr, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_debug_vaddr, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_debugInfo_eliminatedMove, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_debugInfo_renameTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_debugInfo_dispatchTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_debugInfo_enqRsTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_debugInfo_selectTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_debugInfo_issueTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_debugInfo_writebackTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_debugInfo_runahead_checkpoint_id, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_debugInfo_tlbFirstReqTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_debugInfo_tlbRespTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_24_bits_debug_seqNum, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_valid, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_pdest, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_robIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_exceptionVec_0, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_exceptionVec_1, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_exceptionVec_2, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_exceptionVec_3, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_exceptionVec_4, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_exceptionVec_5, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_exceptionVec_6, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_exceptionVec_7, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_exceptionVec_8, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_exceptionVec_9, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_exceptionVec_10, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_exceptionVec_11, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_exceptionVec_12, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_exceptionVec_13, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_exceptionVec_14, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_exceptionVec_15, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_exceptionVec_16, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_exceptionVec_17, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_exceptionVec_18, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_exceptionVec_19, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_exceptionVec_20, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_exceptionVec_21, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_exceptionVec_22, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_exceptionVec_23, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_flushPipe, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_replay, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_trigger, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_vill, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_vma, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_vta, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_vsew, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_vlmul, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_specVill, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_specVma, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_specVta, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_specVsew, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_specVlmul, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_vm, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_vstart, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_frm, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_fpu_isFP32Instr, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_fpu_isFP64Instr, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_fpu_isReduction, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_vxrm, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_vuopIdx, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_lastUop, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_vmask, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_vl, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_nf, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_veew, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_isReverse, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_isExt, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_isNarrow, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_isDstMask, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_isOpMask, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_isMove, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_isDependOldVd, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_isWritePartVd, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vpu_isVleff, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_oldVdPsrc, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vdIdx, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_vdIdxInField, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_isIndexed, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_isMasked, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_isStrided, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_isWhole, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_isVecLoad, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_vls_isVlm, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_debug_isMMIO, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_debug_isNCIO, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_debug_isPerfCnt, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_debug_paddr, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_debug_vaddr, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_debugInfo_eliminatedMove, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_debugInfo_renameTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_debugInfo_dispatchTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_debugInfo_enqRsTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_debugInfo_selectTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_debugInfo_issueTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_debugInfo_writebackTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_debugInfo_runahead_checkpoint_id, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_debugInfo_tlbFirstReqTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_debugInfo_tlbRespTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_23_bits_debug_seqNum, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_valid, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_pdest, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_robIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_intWen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_exceptionVec_0, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_exceptionVec_1, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_exceptionVec_2, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_exceptionVec_3, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_exceptionVec_4, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_exceptionVec_5, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_exceptionVec_6, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_exceptionVec_7, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_exceptionVec_8, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_exceptionVec_9, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_exceptionVec_10, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_exceptionVec_11, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_exceptionVec_12, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_exceptionVec_13, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_exceptionVec_14, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_exceptionVec_15, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_exceptionVec_16, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_exceptionVec_17, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_exceptionVec_18, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_exceptionVec_19, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_exceptionVec_20, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_exceptionVec_21, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_exceptionVec_22, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_exceptionVec_23, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_flushPipe, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_replay, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_lqIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_lqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_trigger, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_predecodeInfo_valid, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_predecodeInfo_isRVC, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_predecodeInfo_brType, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_predecodeInfo_isCall, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_predecodeInfo_isRet, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_debug_isMMIO, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_debug_isNCIO, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_debug_isPerfCnt, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_debug_paddr, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_debug_vaddr, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_debugInfo_eliminatedMove, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_debugInfo_renameTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_debugInfo_dispatchTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_debugInfo_enqRsTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_debugInfo_selectTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_debugInfo_issueTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_debugInfo_writebackTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_debugInfo_runahead_checkpoint_id, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_debugInfo_tlbFirstReqTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_debugInfo_tlbRespTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_22_bits_debug_seqNum, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_valid, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_pdest, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_robIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_intWen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_exceptionVec_0, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_exceptionVec_1, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_exceptionVec_2, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_exceptionVec_3, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_exceptionVec_4, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_exceptionVec_5, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_exceptionVec_6, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_exceptionVec_7, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_exceptionVec_8, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_exceptionVec_9, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_exceptionVec_10, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_exceptionVec_11, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_exceptionVec_12, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_exceptionVec_13, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_exceptionVec_14, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_exceptionVec_15, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_exceptionVec_16, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_exceptionVec_17, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_exceptionVec_18, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_exceptionVec_19, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_exceptionVec_20, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_exceptionVec_21, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_exceptionVec_22, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_exceptionVec_23, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_flushPipe, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_replay, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_lqIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_lqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_trigger, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_predecodeInfo_valid, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_predecodeInfo_isRVC, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_predecodeInfo_brType, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_predecodeInfo_isCall, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_predecodeInfo_isRet, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_debug_isMMIO, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_debug_isNCIO, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_debug_isPerfCnt, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_debug_paddr, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_debug_vaddr, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_debugInfo_eliminatedMove, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_debugInfo_renameTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_debugInfo_dispatchTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_debugInfo_enqRsTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_debugInfo_selectTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_debugInfo_issueTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_debugInfo_writebackTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_debugInfo_runahead_checkpoint_id, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_debugInfo_tlbFirstReqTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_debugInfo_tlbRespTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_21_bits_debug_seqNum, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_valid, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_pdest, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_robIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_intWen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_exceptionVec_0, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_exceptionVec_1, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_exceptionVec_2, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_exceptionVec_3, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_exceptionVec_4, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_exceptionVec_5, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_exceptionVec_6, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_exceptionVec_7, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_exceptionVec_8, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_exceptionVec_9, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_exceptionVec_10, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_exceptionVec_11, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_exceptionVec_12, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_exceptionVec_13, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_exceptionVec_14, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_exceptionVec_15, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_exceptionVec_16, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_exceptionVec_17, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_exceptionVec_18, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_exceptionVec_19, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_exceptionVec_20, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_exceptionVec_21, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_exceptionVec_22, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_exceptionVec_23, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_flushPipe, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_replay, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_lqIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_lqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_trigger, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_predecodeInfo_valid, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_predecodeInfo_isRVC, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_predecodeInfo_brType, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_predecodeInfo_isCall, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_predecodeInfo_isRet, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_debug_isMMIO, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_debug_isNCIO, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_debug_isPerfCnt, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_debug_paddr, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_debug_vaddr, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_debugInfo_eliminatedMove, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_debugInfo_renameTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_debugInfo_dispatchTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_debugInfo_enqRsTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_debugInfo_selectTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_debugInfo_issueTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_debugInfo_writebackTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_debugInfo_runahead_checkpoint_id, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_debugInfo_tlbFirstReqTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_debugInfo_tlbRespTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_20_bits_debug_seqNum, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_valid, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_pdest, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_robIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_intWen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_exceptionVec_0, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_exceptionVec_1, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_exceptionVec_2, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_exceptionVec_3, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_exceptionVec_4, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_exceptionVec_5, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_exceptionVec_6, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_exceptionVec_7, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_exceptionVec_8, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_exceptionVec_9, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_exceptionVec_10, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_exceptionVec_11, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_exceptionVec_12, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_exceptionVec_13, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_exceptionVec_14, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_exceptionVec_15, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_exceptionVec_16, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_exceptionVec_17, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_exceptionVec_18, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_exceptionVec_19, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_exceptionVec_20, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_exceptionVec_21, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_exceptionVec_22, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_exceptionVec_23, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_flushPipe, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_sqIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_sqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_trigger, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_debug_isMMIO, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_debug_isNCIO, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_debug_isPerfCnt, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_debug_paddr, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_debug_vaddr, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_debugInfo_eliminatedMove, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_debugInfo_renameTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_debugInfo_dispatchTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_debugInfo_enqRsTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_debugInfo_selectTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_debugInfo_issueTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_debugInfo_writebackTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_debugInfo_runahead_checkpoint_id, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_debugInfo_tlbFirstReqTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_debugInfo_tlbRespTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_19_bits_debug_seqNum, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_valid, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_pdest, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_robIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_intWen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_exceptionVec_0, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_exceptionVec_1, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_exceptionVec_2, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_exceptionVec_3, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_exceptionVec_4, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_exceptionVec_5, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_exceptionVec_6, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_exceptionVec_7, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_exceptionVec_8, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_exceptionVec_9, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_exceptionVec_10, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_exceptionVec_11, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_exceptionVec_12, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_exceptionVec_13, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_exceptionVec_14, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_exceptionVec_15, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_exceptionVec_16, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_exceptionVec_17, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_exceptionVec_18, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_exceptionVec_19, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_exceptionVec_20, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_exceptionVec_21, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_exceptionVec_22, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_exceptionVec_23, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_flushPipe, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_sqIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_sqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_trigger, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_debug_isMMIO, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_debug_isNCIO, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_debug_isPerfCnt, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_debug_paddr, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_debug_vaddr, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_debugInfo_eliminatedMove, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_debugInfo_renameTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_debugInfo_dispatchTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_debugInfo_enqRsTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_debugInfo_selectTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_debugInfo_issueTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_debugInfo_writebackTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_debugInfo_runahead_checkpoint_id, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_debugInfo_tlbFirstReqTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_debugInfo_tlbRespTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_18_bits_debug_seqNum, UVM_ALL_ON);
        `uvm_field_int(io_writeback_17_valid, UVM_ALL_ON);
        `uvm_field_int(io_writeback_17_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_writeback_17_bits_data_1, UVM_ALL_ON);
        `uvm_field_int(io_writeback_17_bits_data_2, UVM_ALL_ON);
        `uvm_field_int(io_writeback_17_bits_pdest, UVM_ALL_ON);
        `uvm_field_int(io_writeback_17_bits_robIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_writeback_17_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_writeback_17_bits_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_17_bits_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_17_bits_fflags, UVM_ALL_ON);
        `uvm_field_int(io_writeback_17_bits_wflags, UVM_ALL_ON);
        `uvm_field_int(io_writeback_17_bits_debugInfo_eliminatedMove, UVM_ALL_ON);
        `uvm_field_int(io_writeback_17_bits_debugInfo_renameTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_17_bits_debugInfo_dispatchTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_17_bits_debugInfo_enqRsTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_17_bits_debugInfo_selectTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_17_bits_debugInfo_issueTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_17_bits_debugInfo_writebackTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_17_bits_debugInfo_runahead_checkpoint_id, UVM_ALL_ON);
        `uvm_field_int(io_writeback_17_bits_debugInfo_tlbFirstReqTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_17_bits_debugInfo_tlbRespTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_17_bits_debug_seqNum, UVM_ALL_ON);
        `uvm_field_int(io_writeback_16_valid, UVM_ALL_ON);
        `uvm_field_int(io_writeback_16_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_writeback_16_bits_data_1, UVM_ALL_ON);
        `uvm_field_int(io_writeback_16_bits_data_2, UVM_ALL_ON);
        `uvm_field_int(io_writeback_16_bits_data_3, UVM_ALL_ON);
        `uvm_field_int(io_writeback_16_bits_pdest, UVM_ALL_ON);
        `uvm_field_int(io_writeback_16_bits_robIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_writeback_16_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_writeback_16_bits_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_16_bits_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_16_bits_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_16_bits_fflags, UVM_ALL_ON);
        `uvm_field_int(io_writeback_16_bits_wflags, UVM_ALL_ON);
        `uvm_field_int(io_writeback_16_bits_debugInfo_eliminatedMove, UVM_ALL_ON);
        `uvm_field_int(io_writeback_16_bits_debugInfo_renameTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_16_bits_debugInfo_dispatchTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_16_bits_debugInfo_enqRsTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_16_bits_debugInfo_selectTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_16_bits_debugInfo_issueTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_16_bits_debugInfo_writebackTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_16_bits_debugInfo_runahead_checkpoint_id, UVM_ALL_ON);
        `uvm_field_int(io_writeback_16_bits_debugInfo_tlbFirstReqTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_16_bits_debugInfo_tlbRespTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_16_bits_debug_seqNum, UVM_ALL_ON);
        `uvm_field_int(io_writeback_15_valid, UVM_ALL_ON);
        `uvm_field_int(io_writeback_15_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_writeback_15_bits_data_1, UVM_ALL_ON);
        `uvm_field_int(io_writeback_15_bits_data_2, UVM_ALL_ON);
        `uvm_field_int(io_writeback_15_bits_pdest, UVM_ALL_ON);
        `uvm_field_int(io_writeback_15_bits_robIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_writeback_15_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_writeback_15_bits_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_15_bits_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_15_bits_fflags, UVM_ALL_ON);
        `uvm_field_int(io_writeback_15_bits_wflags, UVM_ALL_ON);
        `uvm_field_int(io_writeback_15_bits_vxsat, UVM_ALL_ON);
        `uvm_field_int(io_writeback_15_bits_debugInfo_eliminatedMove, UVM_ALL_ON);
        `uvm_field_int(io_writeback_15_bits_debugInfo_renameTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_15_bits_debugInfo_dispatchTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_15_bits_debugInfo_enqRsTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_15_bits_debugInfo_selectTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_15_bits_debugInfo_issueTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_15_bits_debugInfo_writebackTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_15_bits_debugInfo_runahead_checkpoint_id, UVM_ALL_ON);
        `uvm_field_int(io_writeback_15_bits_debugInfo_tlbFirstReqTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_15_bits_debugInfo_tlbRespTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_15_bits_debug_seqNum, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_valid, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_bits_data_1, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_bits_data_2, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_bits_data_3, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_bits_data_4, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_bits_data_5, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_bits_pdest, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_bits_robIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_bits_intWen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_bits_fpWen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_bits_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_bits_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_bits_vlWen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_bits_fflags, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_bits_wflags, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_bits_exceptionVec_2, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_bits_debugInfo_eliminatedMove, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_bits_debugInfo_renameTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_bits_debugInfo_dispatchTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_bits_debugInfo_enqRsTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_bits_debugInfo_selectTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_bits_debugInfo_issueTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_bits_debugInfo_writebackTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_bits_debugInfo_runahead_checkpoint_id, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_bits_debugInfo_tlbFirstReqTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_bits_debugInfo_tlbRespTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_14_bits_debug_seqNum, UVM_ALL_ON);
        `uvm_field_int(io_writeback_13_valid, UVM_ALL_ON);
        `uvm_field_int(io_writeback_13_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_writeback_13_bits_data_1, UVM_ALL_ON);
        `uvm_field_int(io_writeback_13_bits_data_2, UVM_ALL_ON);
        `uvm_field_int(io_writeback_13_bits_pdest, UVM_ALL_ON);
        `uvm_field_int(io_writeback_13_bits_robIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_writeback_13_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_writeback_13_bits_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_13_bits_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_13_bits_fflags, UVM_ALL_ON);
        `uvm_field_int(io_writeback_13_bits_wflags, UVM_ALL_ON);
        `uvm_field_int(io_writeback_13_bits_vxsat, UVM_ALL_ON);
        `uvm_field_int(io_writeback_13_bits_exceptionVec_2, UVM_ALL_ON);
        `uvm_field_int(io_writeback_13_bits_debugInfo_eliminatedMove, UVM_ALL_ON);
        `uvm_field_int(io_writeback_13_bits_debugInfo_renameTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_13_bits_debugInfo_dispatchTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_13_bits_debugInfo_enqRsTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_13_bits_debugInfo_selectTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_13_bits_debugInfo_issueTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_13_bits_debugInfo_writebackTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_13_bits_debugInfo_runahead_checkpoint_id, UVM_ALL_ON);
        `uvm_field_int(io_writeback_13_bits_debugInfo_tlbFirstReqTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_13_bits_debugInfo_tlbRespTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_13_bits_debug_seqNum, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_valid, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_data_1, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_pdest, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_robIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_intWen, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_valid, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_isRVC, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_robIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_ftqIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_ftqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_ftqOffset, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_level, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_interrupt, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_pc, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_ssp, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_sctr, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_ghr, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_target, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_taken, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_shift, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_fullTarget, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_stFtqIdx_flag, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_stFtqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_stFtqOffset, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_debugIsCtrl, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_redirect_bits_debugIsMemVio, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_exceptionVec_2, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_exceptionVec_3, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_exceptionVec_8, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_exceptionVec_9, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_exceptionVec_10, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_exceptionVec_11, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_exceptionVec_22, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_flushPipe, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_predecodeInfo_valid, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_predecodeInfo_isRVC, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_predecodeInfo_brType, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_predecodeInfo_isCall, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_predecodeInfo_isRet, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_debug_isPerfCnt, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_debugInfo_eliminatedMove, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_debugInfo_renameTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_debugInfo_dispatchTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_debugInfo_enqRsTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_debugInfo_selectTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_debugInfo_issueTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_debugInfo_writebackTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_debugInfo_runahead_checkpoint_id, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_debugInfo_tlbFirstReqTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_debugInfo_tlbRespTime, UVM_ALL_ON);
        `uvm_field_int(io_writeback_7_bits_debug_seqNum, UVM_ALL_ON);
        `uvm_field_int(io_writeback_5_valid, UVM_ALL_ON);
        `uvm_field_int(io_writeback_5_bits_redirect_valid, UVM_ALL_ON);
        `uvm_field_int(io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred, UVM_ALL_ON);
        `uvm_field_int(io_writeback_3_valid, UVM_ALL_ON);
        `uvm_field_int(io_writeback_3_bits_redirect_valid, UVM_ALL_ON);
        `uvm_field_int(io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred, UVM_ALL_ON);
        `uvm_field_int(io_writeback_1_valid, UVM_ALL_ON);
        `uvm_field_int(io_writeback_1_bits_redirect_valid, UVM_ALL_ON);
        `uvm_field_int(io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_26_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_26_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_25_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_25_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_24_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_24_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_24_bits_pdest, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_24_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_24_bits_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_24_bits_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_24_bits_vls_vdIdx, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_24_bits_debug_isMMIO, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_24_bits_debug_isNCIO, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_24_bits_debug_isPerfCnt, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_24_bits_debug_paddr, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_23_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_23_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_23_bits_pdest, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_23_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_23_bits_vecWen, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_23_bits_v0Wen, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_23_bits_vls_vdIdx, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_23_bits_debug_isMMIO, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_23_bits_debug_isNCIO, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_23_bits_debug_isPerfCnt, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_23_bits_debug_paddr, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_22_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_22_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_22_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_22_bits_lqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_22_bits_debug_isMMIO, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_22_bits_debug_isNCIO, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_22_bits_debug_isPerfCnt, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_22_bits_debug_paddr, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_21_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_21_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_21_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_21_bits_lqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_21_bits_debug_isMMIO, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_21_bits_debug_isNCIO, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_21_bits_debug_isPerfCnt, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_21_bits_debug_paddr, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_20_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_20_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_20_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_20_bits_lqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_20_bits_debug_isMMIO, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_20_bits_debug_isNCIO, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_20_bits_debug_isPerfCnt, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_20_bits_debug_paddr, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_19_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_19_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_19_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_19_bits_sqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_19_bits_debug_isMMIO, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_19_bits_debug_isNCIO, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_19_bits_debug_isPerfCnt, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_19_bits_debug_paddr, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_18_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_18_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_18_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_18_bits_sqIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_18_bits_debug_isMMIO, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_18_bits_debug_isNCIO, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_18_bits_debug_isPerfCnt, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_18_bits_debug_paddr, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_17_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_17_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_17_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_17_bits_fflags, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_17_bits_wflags, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_16_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_16_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_16_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_16_bits_fflags, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_16_bits_wflags, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_15_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_15_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_15_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_15_bits_fflags, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_15_bits_wflags, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_15_bits_vxsat, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_14_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_14_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_14_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_14_bits_fflags, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_14_bits_wflags, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_13_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_13_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_13_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_13_bits_fflags, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_13_bits_wflags, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_13_bits_vxsat, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_12_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_12_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_12_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_12_bits_fflags, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_12_bits_wflags, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_11_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_11_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_11_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_11_bits_fflags, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_11_bits_wflags, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_10_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_10_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_10_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_10_bits_fflags, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_10_bits_wflags, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_9_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_9_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_9_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_9_bits_fflags, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_9_bits_wflags, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_8_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_8_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_8_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_8_bits_fflags, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_8_bits_wflags, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_7_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_7_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_7_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_7_bits_debug_isPerfCnt, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_6_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_6_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_6_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_5_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_5_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_5_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_5_bits_redirect_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_5_bits_fflags, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_5_bits_wflags, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_4_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_4_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_4_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_3_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_3_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_3_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_3_bits_redirect_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_2_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_2_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_2_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_1_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_1_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_1_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_1_bits_redirect_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_0_valid, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_0_bits_data_0, UVM_ALL_ON);
        `uvm_field_int(io_exuWriteback_0_bits_robIdx_value, UVM_ALL_ON);
        `uvm_field_int(io_writebackNums_0_bits, UVM_ALL_ON);
        `uvm_field_int(io_writebackNums_1_bits, UVM_ALL_ON);
        `uvm_field_int(io_writebackNums_2_bits, UVM_ALL_ON);
        `uvm_field_int(io_writebackNums_3_bits, UVM_ALL_ON);
        `uvm_field_int(io_writebackNums_4_bits, UVM_ALL_ON);
        `uvm_field_int(io_writebackNums_5_bits, UVM_ALL_ON);
        `uvm_field_int(io_writebackNums_6_bits, UVM_ALL_ON);
        `uvm_field_int(io_writebackNums_7_bits, UVM_ALL_ON);
        `uvm_field_int(io_writebackNums_8_bits, UVM_ALL_ON);
        `uvm_field_int(io_writebackNums_9_bits, UVM_ALL_ON);
        `uvm_field_int(io_writebackNums_10_bits, UVM_ALL_ON);
        `uvm_field_int(io_writebackNums_11_bits, UVM_ALL_ON);
        `uvm_field_int(io_writebackNums_12_bits, UVM_ALL_ON);
        `uvm_field_int(io_writebackNums_13_bits, UVM_ALL_ON);
        `uvm_field_int(io_writebackNums_14_bits, UVM_ALL_ON);
        `uvm_field_int(io_writebackNums_15_bits, UVM_ALL_ON);
        `uvm_field_int(io_writebackNums_16_bits, UVM_ALL_ON);
        `uvm_field_int(io_writebackNums_17_bits, UVM_ALL_ON);
        `uvm_field_int(io_writebackNums_18_bits, UVM_ALL_ON);
        `uvm_field_int(io_writebackNums_19_bits, UVM_ALL_ON);
        `uvm_field_int(io_writebackNums_20_bits, UVM_ALL_ON);
        `uvm_field_int(io_writebackNums_21_bits, UVM_ALL_ON);
        `uvm_field_int(io_writebackNums_22_bits, UVM_ALL_ON);
        `uvm_field_int(io_writebackNums_23_bits, UVM_ALL_ON);
        `uvm_field_int(io_writebackNums_24_bits, UVM_ALL_ON);
        `uvm_field_int(io_writebackNeedFlush_0, UVM_ALL_ON);
        `uvm_field_int(io_writebackNeedFlush_1, UVM_ALL_ON);
        `uvm_field_int(io_writebackNeedFlush_2, UVM_ALL_ON);
        `uvm_field_int(io_writebackNeedFlush_6, UVM_ALL_ON);
        `uvm_field_int(io_writebackNeedFlush_7, UVM_ALL_ON);
        `uvm_field_int(io_writebackNeedFlush_8, UVM_ALL_ON);
        `uvm_field_int(io_writebackNeedFlush_9, UVM_ALL_ON);
        `uvm_field_int(io_writebackNeedFlush_10, UVM_ALL_ON);
        `uvm_field_int(io_writebackNeedFlush_11, UVM_ALL_ON);
        `uvm_field_int(io_writebackNeedFlush_12, UVM_ALL_ON);

    `uvm_object_utils_end

endclass:WriteBack_in_agent_xaction

constraint WriteBack_in_agent_xaction::default_io_writeback_24_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_pdest_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_robIdx_flag_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vecWen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_v0Wen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vlWen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_exceptionVec_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_exceptionVec_1_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_exceptionVec_2_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_exceptionVec_3_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_exceptionVec_4_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_exceptionVec_5_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_exceptionVec_6_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_exceptionVec_7_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_exceptionVec_8_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_exceptionVec_9_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_exceptionVec_10_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_exceptionVec_11_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_exceptionVec_12_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_exceptionVec_13_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_exceptionVec_14_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_exceptionVec_15_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_exceptionVec_16_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_exceptionVec_17_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_exceptionVec_18_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_exceptionVec_19_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_exceptionVec_20_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_exceptionVec_21_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_exceptionVec_22_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_exceptionVec_23_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_flushPipe_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_replay_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_trigger_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_vill_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_vma_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_vta_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_vsew_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_vlmul_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_specVill_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_specVma_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_specVta_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_specVsew_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_specVlmul_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_vm_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_vstart_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_frm_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_fpu_isFP32Instr_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_fpu_isFP64Instr_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_fpu_isReduction_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_vxrm_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_vuopIdx_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_lastUop_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_vmask_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_vl_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_nf_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_veew_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_isReverse_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_isExt_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_isNarrow_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_isDstMask_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_isOpMask_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_isMove_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_isDependOldVd_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_isWritePartVd_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vpu_isVleff_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_oldVdPsrc_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vdIdx_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_vdIdxInField_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_isIndexed_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_isMasked_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_isStrided_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_isWhole_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_isVecLoad_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_vls_isVlm_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_debug_isMMIO_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_debug_isNCIO_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_debug_isPerfCnt_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_debug_paddr_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_debug_vaddr_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_debugInfo_eliminatedMove_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_debugInfo_renameTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_debugInfo_dispatchTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_debugInfo_enqRsTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_debugInfo_selectTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_debugInfo_issueTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_debugInfo_writebackTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_debugInfo_runahead_checkpoint_id_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_debugInfo_tlbFirstReqTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_debugInfo_tlbRespTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_24_bits_debug_seqNum_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_pdest_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_robIdx_flag_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vecWen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_v0Wen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vlWen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_exceptionVec_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_exceptionVec_1_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_exceptionVec_2_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_exceptionVec_3_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_exceptionVec_4_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_exceptionVec_5_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_exceptionVec_6_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_exceptionVec_7_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_exceptionVec_8_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_exceptionVec_9_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_exceptionVec_10_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_exceptionVec_11_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_exceptionVec_12_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_exceptionVec_13_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_exceptionVec_14_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_exceptionVec_15_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_exceptionVec_16_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_exceptionVec_17_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_exceptionVec_18_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_exceptionVec_19_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_exceptionVec_20_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_exceptionVec_21_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_exceptionVec_22_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_exceptionVec_23_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_flushPipe_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_replay_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_trigger_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_vill_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_vma_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_vta_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_vsew_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_vlmul_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_specVill_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_specVma_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_specVta_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_specVsew_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_specVlmul_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_vm_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_vstart_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_frm_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_fpu_isFP32Instr_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_fpu_isFP64Instr_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_fpu_isReduction_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_vxrm_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_vuopIdx_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_lastUop_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_vmask_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_vl_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_nf_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_veew_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_isReverse_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_isExt_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_isNarrow_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_isDstMask_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_isOpMask_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_isMove_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_isDependOldVd_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_isWritePartVd_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vpu_isVleff_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_oldVdPsrc_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vdIdx_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_vdIdxInField_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_isIndexed_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_isMasked_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_isStrided_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_isWhole_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_isVecLoad_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_vls_isVlm_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_debug_isMMIO_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_debug_isNCIO_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_debug_isPerfCnt_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_debug_paddr_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_debug_vaddr_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_debugInfo_eliminatedMove_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_debugInfo_renameTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_debugInfo_dispatchTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_debugInfo_enqRsTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_debugInfo_selectTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_debugInfo_issueTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_debugInfo_writebackTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_debugInfo_runahead_checkpoint_id_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_debugInfo_tlbFirstReqTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_debugInfo_tlbRespTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_23_bits_debug_seqNum_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_pdest_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_robIdx_flag_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_intWen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_fpWen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_exceptionVec_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_exceptionVec_1_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_exceptionVec_2_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_exceptionVec_3_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_exceptionVec_4_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_exceptionVec_5_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_exceptionVec_6_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_exceptionVec_7_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_exceptionVec_8_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_exceptionVec_9_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_exceptionVec_10_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_exceptionVec_11_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_exceptionVec_12_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_exceptionVec_13_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_exceptionVec_14_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_exceptionVec_15_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_exceptionVec_16_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_exceptionVec_17_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_exceptionVec_18_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_exceptionVec_19_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_exceptionVec_20_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_exceptionVec_21_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_exceptionVec_22_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_exceptionVec_23_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_flushPipe_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_replay_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_lqIdx_flag_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_lqIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_trigger_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_predecodeInfo_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_predecodeInfo_isRVC_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_predecodeInfo_brType_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_predecodeInfo_isCall_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_predecodeInfo_isRet_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_debug_isMMIO_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_debug_isNCIO_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_debug_isPerfCnt_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_debug_paddr_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_debug_vaddr_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_debugInfo_eliminatedMove_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_debugInfo_renameTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_debugInfo_dispatchTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_debugInfo_enqRsTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_debugInfo_selectTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_debugInfo_issueTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_debugInfo_writebackTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_debugInfo_runahead_checkpoint_id_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_debugInfo_tlbFirstReqTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_debugInfo_tlbRespTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_22_bits_debug_seqNum_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_pdest_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_robIdx_flag_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_intWen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_fpWen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_exceptionVec_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_exceptionVec_1_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_exceptionVec_2_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_exceptionVec_3_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_exceptionVec_4_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_exceptionVec_5_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_exceptionVec_6_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_exceptionVec_7_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_exceptionVec_8_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_exceptionVec_9_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_exceptionVec_10_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_exceptionVec_11_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_exceptionVec_12_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_exceptionVec_13_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_exceptionVec_14_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_exceptionVec_15_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_exceptionVec_16_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_exceptionVec_17_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_exceptionVec_18_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_exceptionVec_19_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_exceptionVec_20_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_exceptionVec_21_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_exceptionVec_22_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_exceptionVec_23_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_flushPipe_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_replay_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_lqIdx_flag_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_lqIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_trigger_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_predecodeInfo_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_predecodeInfo_isRVC_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_predecodeInfo_brType_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_predecodeInfo_isCall_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_predecodeInfo_isRet_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_debug_isMMIO_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_debug_isNCIO_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_debug_isPerfCnt_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_debug_paddr_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_debug_vaddr_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_debugInfo_eliminatedMove_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_debugInfo_renameTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_debugInfo_dispatchTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_debugInfo_enqRsTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_debugInfo_selectTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_debugInfo_issueTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_debugInfo_writebackTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_debugInfo_runahead_checkpoint_id_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_debugInfo_tlbFirstReqTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_debugInfo_tlbRespTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_21_bits_debug_seqNum_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_pdest_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_robIdx_flag_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_intWen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_fpWen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_exceptionVec_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_exceptionVec_1_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_exceptionVec_2_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_exceptionVec_3_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_exceptionVec_4_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_exceptionVec_5_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_exceptionVec_6_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_exceptionVec_7_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_exceptionVec_8_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_exceptionVec_9_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_exceptionVec_10_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_exceptionVec_11_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_exceptionVec_12_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_exceptionVec_13_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_exceptionVec_14_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_exceptionVec_15_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_exceptionVec_16_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_exceptionVec_17_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_exceptionVec_18_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_exceptionVec_19_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_exceptionVec_20_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_exceptionVec_21_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_exceptionVec_22_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_exceptionVec_23_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_flushPipe_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_replay_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_lqIdx_flag_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_lqIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_trigger_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_predecodeInfo_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_predecodeInfo_isRVC_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_predecodeInfo_brType_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_predecodeInfo_isCall_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_predecodeInfo_isRet_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_debug_isMMIO_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_debug_isNCIO_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_debug_isPerfCnt_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_debug_paddr_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_debug_vaddr_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_debugInfo_eliminatedMove_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_debugInfo_renameTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_debugInfo_dispatchTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_debugInfo_enqRsTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_debugInfo_selectTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_debugInfo_issueTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_debugInfo_writebackTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_debugInfo_runahead_checkpoint_id_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_debugInfo_tlbFirstReqTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_debugInfo_tlbRespTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_20_bits_debug_seqNum_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_pdest_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_robIdx_flag_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_intWen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_exceptionVec_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_exceptionVec_1_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_exceptionVec_2_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_exceptionVec_3_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_exceptionVec_4_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_exceptionVec_5_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_exceptionVec_6_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_exceptionVec_7_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_exceptionVec_8_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_exceptionVec_9_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_exceptionVec_10_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_exceptionVec_11_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_exceptionVec_12_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_exceptionVec_13_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_exceptionVec_14_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_exceptionVec_15_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_exceptionVec_16_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_exceptionVec_17_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_exceptionVec_18_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_exceptionVec_19_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_exceptionVec_20_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_exceptionVec_21_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_exceptionVec_22_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_exceptionVec_23_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_flushPipe_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_sqIdx_flag_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_sqIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_trigger_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_debug_isMMIO_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_debug_isNCIO_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_debug_isPerfCnt_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_debug_paddr_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_debug_vaddr_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_debugInfo_eliminatedMove_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_debugInfo_renameTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_debugInfo_dispatchTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_debugInfo_enqRsTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_debugInfo_selectTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_debugInfo_issueTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_debugInfo_writebackTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_debugInfo_runahead_checkpoint_id_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_debugInfo_tlbFirstReqTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_debugInfo_tlbRespTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_19_bits_debug_seqNum_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_pdest_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_robIdx_flag_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_intWen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_exceptionVec_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_exceptionVec_1_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_exceptionVec_2_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_exceptionVec_3_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_exceptionVec_4_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_exceptionVec_5_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_exceptionVec_6_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_exceptionVec_7_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_exceptionVec_8_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_exceptionVec_9_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_exceptionVec_10_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_exceptionVec_11_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_exceptionVec_12_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_exceptionVec_13_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_exceptionVec_14_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_exceptionVec_15_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_exceptionVec_16_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_exceptionVec_17_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_exceptionVec_18_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_exceptionVec_19_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_exceptionVec_20_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_exceptionVec_21_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_exceptionVec_22_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_exceptionVec_23_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_flushPipe_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_sqIdx_flag_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_sqIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_trigger_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_debug_isMMIO_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_debug_isNCIO_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_debug_isPerfCnt_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_debug_paddr_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_debug_vaddr_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_debugInfo_eliminatedMove_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_debugInfo_renameTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_debugInfo_dispatchTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_debugInfo_enqRsTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_debugInfo_selectTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_debugInfo_issueTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_debugInfo_writebackTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_debugInfo_runahead_checkpoint_id_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_debugInfo_tlbFirstReqTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_debugInfo_tlbRespTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_18_bits_debug_seqNum_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_17_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_17_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_17_bits_data_1_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_17_bits_data_2_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_17_bits_pdest_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_17_bits_robIdx_flag_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_17_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_17_bits_vecWen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_17_bits_v0Wen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_17_bits_fflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_17_bits_wflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_17_bits_debugInfo_eliminatedMove_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_17_bits_debugInfo_renameTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_17_bits_debugInfo_dispatchTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_17_bits_debugInfo_enqRsTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_17_bits_debugInfo_selectTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_17_bits_debugInfo_issueTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_17_bits_debugInfo_writebackTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_17_bits_debugInfo_runahead_checkpoint_id_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_17_bits_debugInfo_tlbFirstReqTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_17_bits_debugInfo_tlbRespTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_17_bits_debug_seqNum_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_16_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_16_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_16_bits_data_1_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_16_bits_data_2_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_16_bits_data_3_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_16_bits_pdest_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_16_bits_robIdx_flag_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_16_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_16_bits_fpWen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_16_bits_vecWen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_16_bits_v0Wen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_16_bits_fflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_16_bits_wflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_16_bits_debugInfo_eliminatedMove_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_16_bits_debugInfo_renameTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_16_bits_debugInfo_dispatchTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_16_bits_debugInfo_enqRsTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_16_bits_debugInfo_selectTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_16_bits_debugInfo_issueTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_16_bits_debugInfo_writebackTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_16_bits_debugInfo_runahead_checkpoint_id_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_16_bits_debugInfo_tlbFirstReqTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_16_bits_debugInfo_tlbRespTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_16_bits_debug_seqNum_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_15_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_15_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_15_bits_data_1_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_15_bits_data_2_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_15_bits_pdest_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_15_bits_robIdx_flag_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_15_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_15_bits_vecWen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_15_bits_v0Wen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_15_bits_fflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_15_bits_wflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_15_bits_vxsat_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_15_bits_debugInfo_eliminatedMove_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_15_bits_debugInfo_renameTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_15_bits_debugInfo_dispatchTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_15_bits_debugInfo_enqRsTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_15_bits_debugInfo_selectTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_15_bits_debugInfo_issueTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_15_bits_debugInfo_writebackTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_15_bits_debugInfo_runahead_checkpoint_id_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_15_bits_debugInfo_tlbFirstReqTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_15_bits_debugInfo_tlbRespTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_15_bits_debug_seqNum_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_bits_data_1_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_bits_data_2_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_bits_data_3_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_bits_data_4_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_bits_data_5_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_bits_pdest_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_bits_robIdx_flag_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_bits_intWen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_bits_fpWen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_bits_vecWen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_bits_v0Wen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_bits_vlWen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_bits_fflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_bits_wflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_bits_exceptionVec_2_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_bits_debugInfo_eliminatedMove_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_bits_debugInfo_renameTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_bits_debugInfo_dispatchTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_bits_debugInfo_enqRsTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_bits_debugInfo_selectTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_bits_debugInfo_issueTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_bits_debugInfo_writebackTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_bits_debugInfo_runahead_checkpoint_id_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_bits_debugInfo_tlbFirstReqTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_bits_debugInfo_tlbRespTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_14_bits_debug_seqNum_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_13_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_13_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_13_bits_data_1_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_13_bits_data_2_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_13_bits_pdest_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_13_bits_robIdx_flag_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_13_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_13_bits_vecWen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_13_bits_v0Wen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_13_bits_fflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_13_bits_wflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_13_bits_vxsat_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_13_bits_exceptionVec_2_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_13_bits_debugInfo_eliminatedMove_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_13_bits_debugInfo_renameTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_13_bits_debugInfo_dispatchTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_13_bits_debugInfo_enqRsTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_13_bits_debugInfo_selectTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_13_bits_debugInfo_issueTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_13_bits_debugInfo_writebackTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_13_bits_debugInfo_runahead_checkpoint_id_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_13_bits_debugInfo_tlbFirstReqTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_13_bits_debugInfo_tlbRespTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_13_bits_debug_seqNum_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_data_1_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_pdest_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_robIdx_flag_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_intWen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_isRVC_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_robIdx_flag_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_ftqIdx_flag_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_ftqIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_ftqOffset_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_level_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_interrupt_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_pc_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_ssp_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_sctr_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_ghr_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_target_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_taken_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_shift_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_fullTarget_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_stFtqIdx_flag_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_stFtqIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_stFtqOffset_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_debugIsCtrl_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_redirect_bits_debugIsMemVio_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_exceptionVec_2_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_exceptionVec_3_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_exceptionVec_8_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_exceptionVec_9_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_exceptionVec_10_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_exceptionVec_11_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_exceptionVec_22_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_flushPipe_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_predecodeInfo_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_predecodeInfo_isRVC_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_predecodeInfo_brType_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_predecodeInfo_isCall_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_predecodeInfo_isRet_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_debug_isPerfCnt_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_debugInfo_eliminatedMove_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_debugInfo_renameTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_debugInfo_dispatchTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_debugInfo_enqRsTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_debugInfo_selectTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_debugInfo_issueTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_debugInfo_writebackTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_debugInfo_runahead_checkpoint_id_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_debugInfo_tlbFirstReqTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_debugInfo_tlbRespTime_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_7_bits_debug_seqNum_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_5_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_5_bits_redirect_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_3_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_3_bits_redirect_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_1_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_1_bits_redirect_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_26_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_26_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_25_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_25_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_24_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_24_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_24_bits_pdest_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_24_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_24_bits_vecWen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_24_bits_v0Wen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_24_bits_vls_vdIdx_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_24_bits_debug_isMMIO_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_24_bits_debug_isNCIO_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_24_bits_debug_isPerfCnt_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_24_bits_debug_paddr_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_23_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_23_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_23_bits_pdest_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_23_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_23_bits_vecWen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_23_bits_v0Wen_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_23_bits_vls_vdIdx_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_23_bits_debug_isMMIO_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_23_bits_debug_isNCIO_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_23_bits_debug_isPerfCnt_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_23_bits_debug_paddr_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_22_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_22_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_22_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_22_bits_lqIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_22_bits_debug_isMMIO_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_22_bits_debug_isNCIO_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_22_bits_debug_isPerfCnt_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_22_bits_debug_paddr_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_21_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_21_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_21_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_21_bits_lqIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_21_bits_debug_isMMIO_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_21_bits_debug_isNCIO_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_21_bits_debug_isPerfCnt_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_21_bits_debug_paddr_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_20_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_20_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_20_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_20_bits_lqIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_20_bits_debug_isMMIO_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_20_bits_debug_isNCIO_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_20_bits_debug_isPerfCnt_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_20_bits_debug_paddr_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_19_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_19_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_19_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_19_bits_sqIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_19_bits_debug_isMMIO_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_19_bits_debug_isNCIO_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_19_bits_debug_isPerfCnt_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_19_bits_debug_paddr_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_18_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_18_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_18_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_18_bits_sqIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_18_bits_debug_isMMIO_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_18_bits_debug_isNCIO_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_18_bits_debug_isPerfCnt_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_18_bits_debug_paddr_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_17_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_17_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_17_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_17_bits_fflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_17_bits_wflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_16_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_16_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_16_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_16_bits_fflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_16_bits_wflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_15_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_15_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_15_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_15_bits_fflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_15_bits_wflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_15_bits_vxsat_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_14_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_14_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_14_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_14_bits_fflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_14_bits_wflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_13_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_13_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_13_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_13_bits_fflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_13_bits_wflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_13_bits_vxsat_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_12_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_12_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_12_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_12_bits_fflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_12_bits_wflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_11_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_11_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_11_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_11_bits_fflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_11_bits_wflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_10_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_10_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_10_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_10_bits_fflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_10_bits_wflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_9_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_9_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_9_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_9_bits_fflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_9_bits_wflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_8_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_8_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_8_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_8_bits_fflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_8_bits_wflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_7_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_7_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_7_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_7_bits_debug_isPerfCnt_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_6_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_6_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_6_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_5_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_5_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_5_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_5_bits_redirect_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_5_bits_fflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_5_bits_wflags_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_4_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_4_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_4_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_3_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_3_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_3_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_3_bits_redirect_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_2_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_2_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_2_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_1_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_1_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_1_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_1_bits_redirect_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_0_valid_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_0_bits_data_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_exuWriteback_0_bits_robIdx_value_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNums_0_bits_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNums_1_bits_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNums_2_bits_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNums_3_bits_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNums_4_bits_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNums_5_bits_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNums_6_bits_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNums_7_bits_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNums_8_bits_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNums_9_bits_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNums_10_bits_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNums_11_bits_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNums_12_bits_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNums_13_bits_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNums_14_bits_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNums_15_bits_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNums_16_bits_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNums_17_bits_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNums_18_bits_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNums_19_bits_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNums_20_bits_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNums_21_bits_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNums_22_bits_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNums_23_bits_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNums_24_bits_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNeedFlush_0_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNeedFlush_1_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNeedFlush_2_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNeedFlush_6_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNeedFlush_7_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNeedFlush_8_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNeedFlush_9_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNeedFlush_10_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNeedFlush_11_cons{

}

constraint WriteBack_in_agent_xaction::default_io_writebackNeedFlush_12_cons{

}

function WriteBack_in_agent_xaction::new(string name = "WriteBack_in_agent_xaction");
    super.new();
endfunction:new

function void WriteBack_in_agent_xaction::pack();
    super.pack();
endfunction:pack
function void WriteBack_in_agent_xaction::unpack();
    super.unpack();
endfunction:unpack
function void WriteBack_in_agent_xaction::pre_randomize();
    super.pre_randomize();
endfunction:pre_randomize
function void WriteBack_in_agent_xaction::post_randomize();
    super.post_randomize();
    //this.pack();
endfunction:post_randomize

function string WriteBack_in_agent_xaction::psdisplay(string prefix = "");
    string pkt_str;
    pkt_str = $sformatf("%s for packet[%0d] >>>>",prefix,this.pkt_index);
    pkt_str = $sformatf("%schannel_id=%0d ",pkt_str,this.channel_id);
    pkt_str = $sformatf("%sstart=%0f finish=%0f >>>>\n",pkt_str,this.start,this.finish);
    //foreach(this.pload_q[i]) begin
    //    pkt_str = $sformatf("%spload_q[%0d]=0x%2h  ",pkt_str,i,this.pload_q[i]);
    //end
    pkt_str = $sformatf("%sio_writeback_24_valid = 0x%0h ",pkt_str,this.io_writeback_24_valid);
    pkt_str = $sformatf("%sio_writeback_24_bits_data_0 = 0x%0h ",pkt_str,this.io_writeback_24_bits_data_0);
    pkt_str = $sformatf("%sio_writeback_24_bits_pdest = 0x%0h ",pkt_str,this.io_writeback_24_bits_pdest);
    pkt_str = $sformatf("%sio_writeback_24_bits_robIdx_flag = 0x%0h ",pkt_str,this.io_writeback_24_bits_robIdx_flag);
    pkt_str = $sformatf("%sio_writeback_24_bits_robIdx_value = 0x%0h ",pkt_str,this.io_writeback_24_bits_robIdx_value);
    pkt_str = $sformatf("%sio_writeback_24_bits_vecWen = 0x%0h ",pkt_str,this.io_writeback_24_bits_vecWen);
    pkt_str = $sformatf("%sio_writeback_24_bits_v0Wen = 0x%0h ",pkt_str,this.io_writeback_24_bits_v0Wen);
    pkt_str = $sformatf("%sio_writeback_24_bits_vlWen = 0x%0h ",pkt_str,this.io_writeback_24_bits_vlWen);
    pkt_str = $sformatf("%sio_writeback_24_bits_exceptionVec_0 = 0x%0h ",pkt_str,this.io_writeback_24_bits_exceptionVec_0);
    pkt_str = $sformatf("%sio_writeback_24_bits_exceptionVec_1 = 0x%0h ",pkt_str,this.io_writeback_24_bits_exceptionVec_1);
    pkt_str = $sformatf("%sio_writeback_24_bits_exceptionVec_2 = 0x%0h ",pkt_str,this.io_writeback_24_bits_exceptionVec_2);
    pkt_str = $sformatf("%sio_writeback_24_bits_exceptionVec_3 = 0x%0h ",pkt_str,this.io_writeback_24_bits_exceptionVec_3);
    pkt_str = $sformatf("%sio_writeback_24_bits_exceptionVec_4 = 0x%0h ",pkt_str,this.io_writeback_24_bits_exceptionVec_4);
    pkt_str = $sformatf("%sio_writeback_24_bits_exceptionVec_5 = 0x%0h ",pkt_str,this.io_writeback_24_bits_exceptionVec_5);
    pkt_str = $sformatf("%sio_writeback_24_bits_exceptionVec_6 = 0x%0h ",pkt_str,this.io_writeback_24_bits_exceptionVec_6);
    pkt_str = $sformatf("%sio_writeback_24_bits_exceptionVec_7 = 0x%0h ",pkt_str,this.io_writeback_24_bits_exceptionVec_7);
    pkt_str = $sformatf("%sio_writeback_24_bits_exceptionVec_8 = 0x%0h ",pkt_str,this.io_writeback_24_bits_exceptionVec_8);
    pkt_str = $sformatf("%sio_writeback_24_bits_exceptionVec_9 = 0x%0h ",pkt_str,this.io_writeback_24_bits_exceptionVec_9);
    pkt_str = $sformatf("%sio_writeback_24_bits_exceptionVec_10 = 0x%0h ",pkt_str,this.io_writeback_24_bits_exceptionVec_10);
    pkt_str = $sformatf("%sio_writeback_24_bits_exceptionVec_11 = 0x%0h ",pkt_str,this.io_writeback_24_bits_exceptionVec_11);
    pkt_str = $sformatf("%sio_writeback_24_bits_exceptionVec_12 = 0x%0h ",pkt_str,this.io_writeback_24_bits_exceptionVec_12);
    pkt_str = $sformatf("%sio_writeback_24_bits_exceptionVec_13 = 0x%0h ",pkt_str,this.io_writeback_24_bits_exceptionVec_13);
    pkt_str = $sformatf("%sio_writeback_24_bits_exceptionVec_14 = 0x%0h ",pkt_str,this.io_writeback_24_bits_exceptionVec_14);
    pkt_str = $sformatf("%sio_writeback_24_bits_exceptionVec_15 = 0x%0h ",pkt_str,this.io_writeback_24_bits_exceptionVec_15);
    pkt_str = $sformatf("%sio_writeback_24_bits_exceptionVec_16 = 0x%0h ",pkt_str,this.io_writeback_24_bits_exceptionVec_16);
    pkt_str = $sformatf("%sio_writeback_24_bits_exceptionVec_17 = 0x%0h ",pkt_str,this.io_writeback_24_bits_exceptionVec_17);
    pkt_str = $sformatf("%sio_writeback_24_bits_exceptionVec_18 = 0x%0h ",pkt_str,this.io_writeback_24_bits_exceptionVec_18);
    pkt_str = $sformatf("%sio_writeback_24_bits_exceptionVec_19 = 0x%0h ",pkt_str,this.io_writeback_24_bits_exceptionVec_19);
    pkt_str = $sformatf("%sio_writeback_24_bits_exceptionVec_20 = 0x%0h ",pkt_str,this.io_writeback_24_bits_exceptionVec_20);
    pkt_str = $sformatf("%sio_writeback_24_bits_exceptionVec_21 = 0x%0h ",pkt_str,this.io_writeback_24_bits_exceptionVec_21);
    pkt_str = $sformatf("%sio_writeback_24_bits_exceptionVec_22 = 0x%0h ",pkt_str,this.io_writeback_24_bits_exceptionVec_22);
    pkt_str = $sformatf("%sio_writeback_24_bits_exceptionVec_23 = 0x%0h ",pkt_str,this.io_writeback_24_bits_exceptionVec_23);
    pkt_str = $sformatf("%sio_writeback_24_bits_flushPipe = 0x%0h ",pkt_str,this.io_writeback_24_bits_flushPipe);
    pkt_str = $sformatf("%sio_writeback_24_bits_replay = 0x%0h ",pkt_str,this.io_writeback_24_bits_replay);
    pkt_str = $sformatf("%sio_writeback_24_bits_trigger = 0x%0h ",pkt_str,this.io_writeback_24_bits_trigger);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_vill = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_vill);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_vma = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_vma);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_vta = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_vta);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_vsew = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_vsew);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_vlmul = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_vlmul);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_specVill = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_specVill);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_specVma = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_specVma);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_specVta = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_specVta);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_specVsew = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_specVsew);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_specVlmul = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_specVlmul);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_vm = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_vm);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_vstart = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_vstart);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_frm = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_frm);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_fpu_isFpToVecInst = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_fpu_isFP32Instr = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_fpu_isFP32Instr);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_fpu_isFP64Instr = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_fpu_isFP64Instr);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_fpu_isReduction = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_fpu_isReduction);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2 = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4 = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8 = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_vxrm = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_vxrm);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_vuopIdx = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_vuopIdx);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_lastUop = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_lastUop);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_vmask = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_vmask);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_vl = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_vl);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_nf = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_nf);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_veew = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_veew);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_isReverse = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_isReverse);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_isExt = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_isExt);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_isNarrow = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_isNarrow);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_isDstMask = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_isDstMask);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_isOpMask = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_isOpMask);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_isMove = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_isMove);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_isDependOldVd = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_isDependOldVd);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_isWritePartVd = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_isWritePartVd);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vpu_isVleff = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vpu_isVleff);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_oldVdPsrc = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_oldVdPsrc);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vdIdx = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vdIdx);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_vdIdxInField = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_vdIdxInField);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_isIndexed = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_isIndexed);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_isMasked = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_isMasked);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_isStrided = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_isStrided);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_isWhole = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_isWhole);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_isVecLoad = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_isVecLoad);
    pkt_str = $sformatf("%sio_writeback_24_bits_vls_isVlm = 0x%0h ",pkt_str,this.io_writeback_24_bits_vls_isVlm);
    pkt_str = $sformatf("%sio_writeback_24_bits_debug_isMMIO = 0x%0h ",pkt_str,this.io_writeback_24_bits_debug_isMMIO);
    pkt_str = $sformatf("%sio_writeback_24_bits_debug_isNCIO = 0x%0h ",pkt_str,this.io_writeback_24_bits_debug_isNCIO);
    pkt_str = $sformatf("%sio_writeback_24_bits_debug_isPerfCnt = 0x%0h ",pkt_str,this.io_writeback_24_bits_debug_isPerfCnt);
    pkt_str = $sformatf("%sio_writeback_24_bits_debug_paddr = 0x%0h ",pkt_str,this.io_writeback_24_bits_debug_paddr);
    pkt_str = $sformatf("%sio_writeback_24_bits_debug_vaddr = 0x%0h ",pkt_str,this.io_writeback_24_bits_debug_vaddr);
    pkt_str = $sformatf("%sio_writeback_24_bits_debugInfo_eliminatedMove = 0x%0h ",pkt_str,this.io_writeback_24_bits_debugInfo_eliminatedMove);
    pkt_str = $sformatf("%sio_writeback_24_bits_debugInfo_renameTime = 0x%0h ",pkt_str,this.io_writeback_24_bits_debugInfo_renameTime);
    pkt_str = $sformatf("%sio_writeback_24_bits_debugInfo_dispatchTime = 0x%0h ",pkt_str,this.io_writeback_24_bits_debugInfo_dispatchTime);
    pkt_str = $sformatf("%sio_writeback_24_bits_debugInfo_enqRsTime = 0x%0h ",pkt_str,this.io_writeback_24_bits_debugInfo_enqRsTime);
    pkt_str = $sformatf("%sio_writeback_24_bits_debugInfo_selectTime = 0x%0h ",pkt_str,this.io_writeback_24_bits_debugInfo_selectTime);
    pkt_str = $sformatf("%sio_writeback_24_bits_debugInfo_issueTime = 0x%0h ",pkt_str,this.io_writeback_24_bits_debugInfo_issueTime);
    pkt_str = $sformatf("%sio_writeback_24_bits_debugInfo_writebackTime = 0x%0h ",pkt_str,this.io_writeback_24_bits_debugInfo_writebackTime);
    pkt_str = $sformatf("%sio_writeback_24_bits_debugInfo_runahead_checkpoint_id = 0x%0h ",pkt_str,this.io_writeback_24_bits_debugInfo_runahead_checkpoint_id);
    pkt_str = $sformatf("%sio_writeback_24_bits_debugInfo_tlbFirstReqTime = 0x%0h ",pkt_str,this.io_writeback_24_bits_debugInfo_tlbFirstReqTime);
    pkt_str = $sformatf("%sio_writeback_24_bits_debugInfo_tlbRespTime = 0x%0h ",pkt_str,this.io_writeback_24_bits_debugInfo_tlbRespTime);
    pkt_str = $sformatf("%sio_writeback_24_bits_debug_seqNum = 0x%0h ",pkt_str,this.io_writeback_24_bits_debug_seqNum);
    pkt_str = $sformatf("%sio_writeback_23_valid = 0x%0h ",pkt_str,this.io_writeback_23_valid);
    pkt_str = $sformatf("%sio_writeback_23_bits_data_0 = 0x%0h ",pkt_str,this.io_writeback_23_bits_data_0);
    pkt_str = $sformatf("%sio_writeback_23_bits_pdest = 0x%0h ",pkt_str,this.io_writeback_23_bits_pdest);
    pkt_str = $sformatf("%sio_writeback_23_bits_robIdx_flag = 0x%0h ",pkt_str,this.io_writeback_23_bits_robIdx_flag);
    pkt_str = $sformatf("%sio_writeback_23_bits_robIdx_value = 0x%0h ",pkt_str,this.io_writeback_23_bits_robIdx_value);
    pkt_str = $sformatf("%sio_writeback_23_bits_vecWen = 0x%0h ",pkt_str,this.io_writeback_23_bits_vecWen);
    pkt_str = $sformatf("%sio_writeback_23_bits_v0Wen = 0x%0h ",pkt_str,this.io_writeback_23_bits_v0Wen);
    pkt_str = $sformatf("%sio_writeback_23_bits_vlWen = 0x%0h ",pkt_str,this.io_writeback_23_bits_vlWen);
    pkt_str = $sformatf("%sio_writeback_23_bits_exceptionVec_0 = 0x%0h ",pkt_str,this.io_writeback_23_bits_exceptionVec_0);
    pkt_str = $sformatf("%sio_writeback_23_bits_exceptionVec_1 = 0x%0h ",pkt_str,this.io_writeback_23_bits_exceptionVec_1);
    pkt_str = $sformatf("%sio_writeback_23_bits_exceptionVec_2 = 0x%0h ",pkt_str,this.io_writeback_23_bits_exceptionVec_2);
    pkt_str = $sformatf("%sio_writeback_23_bits_exceptionVec_3 = 0x%0h ",pkt_str,this.io_writeback_23_bits_exceptionVec_3);
    pkt_str = $sformatf("%sio_writeback_23_bits_exceptionVec_4 = 0x%0h ",pkt_str,this.io_writeback_23_bits_exceptionVec_4);
    pkt_str = $sformatf("%sio_writeback_23_bits_exceptionVec_5 = 0x%0h ",pkt_str,this.io_writeback_23_bits_exceptionVec_5);
    pkt_str = $sformatf("%sio_writeback_23_bits_exceptionVec_6 = 0x%0h ",pkt_str,this.io_writeback_23_bits_exceptionVec_6);
    pkt_str = $sformatf("%sio_writeback_23_bits_exceptionVec_7 = 0x%0h ",pkt_str,this.io_writeback_23_bits_exceptionVec_7);
    pkt_str = $sformatf("%sio_writeback_23_bits_exceptionVec_8 = 0x%0h ",pkt_str,this.io_writeback_23_bits_exceptionVec_8);
    pkt_str = $sformatf("%sio_writeback_23_bits_exceptionVec_9 = 0x%0h ",pkt_str,this.io_writeback_23_bits_exceptionVec_9);
    pkt_str = $sformatf("%sio_writeback_23_bits_exceptionVec_10 = 0x%0h ",pkt_str,this.io_writeback_23_bits_exceptionVec_10);
    pkt_str = $sformatf("%sio_writeback_23_bits_exceptionVec_11 = 0x%0h ",pkt_str,this.io_writeback_23_bits_exceptionVec_11);
    pkt_str = $sformatf("%sio_writeback_23_bits_exceptionVec_12 = 0x%0h ",pkt_str,this.io_writeback_23_bits_exceptionVec_12);
    pkt_str = $sformatf("%sio_writeback_23_bits_exceptionVec_13 = 0x%0h ",pkt_str,this.io_writeback_23_bits_exceptionVec_13);
    pkt_str = $sformatf("%sio_writeback_23_bits_exceptionVec_14 = 0x%0h ",pkt_str,this.io_writeback_23_bits_exceptionVec_14);
    pkt_str = $sformatf("%sio_writeback_23_bits_exceptionVec_15 = 0x%0h ",pkt_str,this.io_writeback_23_bits_exceptionVec_15);
    pkt_str = $sformatf("%sio_writeback_23_bits_exceptionVec_16 = 0x%0h ",pkt_str,this.io_writeback_23_bits_exceptionVec_16);
    pkt_str = $sformatf("%sio_writeback_23_bits_exceptionVec_17 = 0x%0h ",pkt_str,this.io_writeback_23_bits_exceptionVec_17);
    pkt_str = $sformatf("%sio_writeback_23_bits_exceptionVec_18 = 0x%0h ",pkt_str,this.io_writeback_23_bits_exceptionVec_18);
    pkt_str = $sformatf("%sio_writeback_23_bits_exceptionVec_19 = 0x%0h ",pkt_str,this.io_writeback_23_bits_exceptionVec_19);
    pkt_str = $sformatf("%sio_writeback_23_bits_exceptionVec_20 = 0x%0h ",pkt_str,this.io_writeback_23_bits_exceptionVec_20);
    pkt_str = $sformatf("%sio_writeback_23_bits_exceptionVec_21 = 0x%0h ",pkt_str,this.io_writeback_23_bits_exceptionVec_21);
    pkt_str = $sformatf("%sio_writeback_23_bits_exceptionVec_22 = 0x%0h ",pkt_str,this.io_writeback_23_bits_exceptionVec_22);
    pkt_str = $sformatf("%sio_writeback_23_bits_exceptionVec_23 = 0x%0h ",pkt_str,this.io_writeback_23_bits_exceptionVec_23);
    pkt_str = $sformatf("%sio_writeback_23_bits_flushPipe = 0x%0h ",pkt_str,this.io_writeback_23_bits_flushPipe);
    pkt_str = $sformatf("%sio_writeback_23_bits_replay = 0x%0h ",pkt_str,this.io_writeback_23_bits_replay);
    pkt_str = $sformatf("%sio_writeback_23_bits_trigger = 0x%0h ",pkt_str,this.io_writeback_23_bits_trigger);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_vill = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_vill);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_vma = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_vma);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_vta = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_vta);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_vsew = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_vsew);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_vlmul = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_vlmul);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_specVill = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_specVill);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_specVma = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_specVma);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_specVta = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_specVta);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_specVsew = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_specVsew);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_specVlmul = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_specVlmul);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_vm = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_vm);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_vstart = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_vstart);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_frm = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_frm);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_fpu_isFpToVecInst = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_fpu_isFP32Instr = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_fpu_isFP32Instr);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_fpu_isFP64Instr = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_fpu_isFP64Instr);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_fpu_isReduction = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_fpu_isReduction);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2 = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4 = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8 = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_vxrm = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_vxrm);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_vuopIdx = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_vuopIdx);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_lastUop = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_lastUop);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_vmask = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_vmask);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_vl = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_vl);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_nf = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_nf);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_veew = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_veew);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_isReverse = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_isReverse);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_isExt = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_isExt);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_isNarrow = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_isNarrow);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_isDstMask = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_isDstMask);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_isOpMask = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_isOpMask);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_isMove = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_isMove);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_isDependOldVd = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_isDependOldVd);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_isWritePartVd = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_isWritePartVd);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vpu_isVleff = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vpu_isVleff);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_oldVdPsrc = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_oldVdPsrc);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vdIdx = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vdIdx);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_vdIdxInField = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_vdIdxInField);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_isIndexed = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_isIndexed);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_isMasked = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_isMasked);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_isStrided = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_isStrided);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_isWhole = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_isWhole);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_isVecLoad = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_isVecLoad);
    pkt_str = $sformatf("%sio_writeback_23_bits_vls_isVlm = 0x%0h ",pkt_str,this.io_writeback_23_bits_vls_isVlm);
    pkt_str = $sformatf("%sio_writeback_23_bits_debug_isMMIO = 0x%0h ",pkt_str,this.io_writeback_23_bits_debug_isMMIO);
    pkt_str = $sformatf("%sio_writeback_23_bits_debug_isNCIO = 0x%0h ",pkt_str,this.io_writeback_23_bits_debug_isNCIO);
    pkt_str = $sformatf("%sio_writeback_23_bits_debug_isPerfCnt = 0x%0h ",pkt_str,this.io_writeback_23_bits_debug_isPerfCnt);
    pkt_str = $sformatf("%sio_writeback_23_bits_debug_paddr = 0x%0h ",pkt_str,this.io_writeback_23_bits_debug_paddr);
    pkt_str = $sformatf("%sio_writeback_23_bits_debug_vaddr = 0x%0h ",pkt_str,this.io_writeback_23_bits_debug_vaddr);
    pkt_str = $sformatf("%sio_writeback_23_bits_debugInfo_eliminatedMove = 0x%0h ",pkt_str,this.io_writeback_23_bits_debugInfo_eliminatedMove);
    pkt_str = $sformatf("%sio_writeback_23_bits_debugInfo_renameTime = 0x%0h ",pkt_str,this.io_writeback_23_bits_debugInfo_renameTime);
    pkt_str = $sformatf("%sio_writeback_23_bits_debugInfo_dispatchTime = 0x%0h ",pkt_str,this.io_writeback_23_bits_debugInfo_dispatchTime);
    pkt_str = $sformatf("%sio_writeback_23_bits_debugInfo_enqRsTime = 0x%0h ",pkt_str,this.io_writeback_23_bits_debugInfo_enqRsTime);
    pkt_str = $sformatf("%sio_writeback_23_bits_debugInfo_selectTime = 0x%0h ",pkt_str,this.io_writeback_23_bits_debugInfo_selectTime);
    pkt_str = $sformatf("%sio_writeback_23_bits_debugInfo_issueTime = 0x%0h ",pkt_str,this.io_writeback_23_bits_debugInfo_issueTime);
    pkt_str = $sformatf("%sio_writeback_23_bits_debugInfo_writebackTime = 0x%0h ",pkt_str,this.io_writeback_23_bits_debugInfo_writebackTime);
    pkt_str = $sformatf("%sio_writeback_23_bits_debugInfo_runahead_checkpoint_id = 0x%0h ",pkt_str,this.io_writeback_23_bits_debugInfo_runahead_checkpoint_id);
    pkt_str = $sformatf("%sio_writeback_23_bits_debugInfo_tlbFirstReqTime = 0x%0h ",pkt_str,this.io_writeback_23_bits_debugInfo_tlbFirstReqTime);
    pkt_str = $sformatf("%sio_writeback_23_bits_debugInfo_tlbRespTime = 0x%0h ",pkt_str,this.io_writeback_23_bits_debugInfo_tlbRespTime);
    pkt_str = $sformatf("%sio_writeback_23_bits_debug_seqNum = 0x%0h ",pkt_str,this.io_writeback_23_bits_debug_seqNum);
    pkt_str = $sformatf("%sio_writeback_22_valid = 0x%0h ",pkt_str,this.io_writeback_22_valid);
    pkt_str = $sformatf("%sio_writeback_22_bits_data_0 = 0x%0h ",pkt_str,this.io_writeback_22_bits_data_0);
    pkt_str = $sformatf("%sio_writeback_22_bits_pdest = 0x%0h ",pkt_str,this.io_writeback_22_bits_pdest);
    pkt_str = $sformatf("%sio_writeback_22_bits_robIdx_flag = 0x%0h ",pkt_str,this.io_writeback_22_bits_robIdx_flag);
    pkt_str = $sformatf("%sio_writeback_22_bits_robIdx_value = 0x%0h ",pkt_str,this.io_writeback_22_bits_robIdx_value);
    pkt_str = $sformatf("%sio_writeback_22_bits_intWen = 0x%0h ",pkt_str,this.io_writeback_22_bits_intWen);
    pkt_str = $sformatf("%sio_writeback_22_bits_fpWen = 0x%0h ",pkt_str,this.io_writeback_22_bits_fpWen);
    pkt_str = $sformatf("%sio_writeback_22_bits_exceptionVec_0 = 0x%0h ",pkt_str,this.io_writeback_22_bits_exceptionVec_0);
    pkt_str = $sformatf("%sio_writeback_22_bits_exceptionVec_1 = 0x%0h ",pkt_str,this.io_writeback_22_bits_exceptionVec_1);
    pkt_str = $sformatf("%sio_writeback_22_bits_exceptionVec_2 = 0x%0h ",pkt_str,this.io_writeback_22_bits_exceptionVec_2);
    pkt_str = $sformatf("%sio_writeback_22_bits_exceptionVec_3 = 0x%0h ",pkt_str,this.io_writeback_22_bits_exceptionVec_3);
    pkt_str = $sformatf("%sio_writeback_22_bits_exceptionVec_4 = 0x%0h ",pkt_str,this.io_writeback_22_bits_exceptionVec_4);
    pkt_str = $sformatf("%sio_writeback_22_bits_exceptionVec_5 = 0x%0h ",pkt_str,this.io_writeback_22_bits_exceptionVec_5);
    pkt_str = $sformatf("%sio_writeback_22_bits_exceptionVec_6 = 0x%0h ",pkt_str,this.io_writeback_22_bits_exceptionVec_6);
    pkt_str = $sformatf("%sio_writeback_22_bits_exceptionVec_7 = 0x%0h ",pkt_str,this.io_writeback_22_bits_exceptionVec_7);
    pkt_str = $sformatf("%sio_writeback_22_bits_exceptionVec_8 = 0x%0h ",pkt_str,this.io_writeback_22_bits_exceptionVec_8);
    pkt_str = $sformatf("%sio_writeback_22_bits_exceptionVec_9 = 0x%0h ",pkt_str,this.io_writeback_22_bits_exceptionVec_9);
    pkt_str = $sformatf("%sio_writeback_22_bits_exceptionVec_10 = 0x%0h ",pkt_str,this.io_writeback_22_bits_exceptionVec_10);
    pkt_str = $sformatf("%sio_writeback_22_bits_exceptionVec_11 = 0x%0h ",pkt_str,this.io_writeback_22_bits_exceptionVec_11);
    pkt_str = $sformatf("%sio_writeback_22_bits_exceptionVec_12 = 0x%0h ",pkt_str,this.io_writeback_22_bits_exceptionVec_12);
    pkt_str = $sformatf("%sio_writeback_22_bits_exceptionVec_13 = 0x%0h ",pkt_str,this.io_writeback_22_bits_exceptionVec_13);
    pkt_str = $sformatf("%sio_writeback_22_bits_exceptionVec_14 = 0x%0h ",pkt_str,this.io_writeback_22_bits_exceptionVec_14);
    pkt_str = $sformatf("%sio_writeback_22_bits_exceptionVec_15 = 0x%0h ",pkt_str,this.io_writeback_22_bits_exceptionVec_15);
    pkt_str = $sformatf("%sio_writeback_22_bits_exceptionVec_16 = 0x%0h ",pkt_str,this.io_writeback_22_bits_exceptionVec_16);
    pkt_str = $sformatf("%sio_writeback_22_bits_exceptionVec_17 = 0x%0h ",pkt_str,this.io_writeback_22_bits_exceptionVec_17);
    pkt_str = $sformatf("%sio_writeback_22_bits_exceptionVec_18 = 0x%0h ",pkt_str,this.io_writeback_22_bits_exceptionVec_18);
    pkt_str = $sformatf("%sio_writeback_22_bits_exceptionVec_19 = 0x%0h ",pkt_str,this.io_writeback_22_bits_exceptionVec_19);
    pkt_str = $sformatf("%sio_writeback_22_bits_exceptionVec_20 = 0x%0h ",pkt_str,this.io_writeback_22_bits_exceptionVec_20);
    pkt_str = $sformatf("%sio_writeback_22_bits_exceptionVec_21 = 0x%0h ",pkt_str,this.io_writeback_22_bits_exceptionVec_21);
    pkt_str = $sformatf("%sio_writeback_22_bits_exceptionVec_22 = 0x%0h ",pkt_str,this.io_writeback_22_bits_exceptionVec_22);
    pkt_str = $sformatf("%sio_writeback_22_bits_exceptionVec_23 = 0x%0h ",pkt_str,this.io_writeback_22_bits_exceptionVec_23);
    pkt_str = $sformatf("%sio_writeback_22_bits_flushPipe = 0x%0h ",pkt_str,this.io_writeback_22_bits_flushPipe);
    pkt_str = $sformatf("%sio_writeback_22_bits_replay = 0x%0h ",pkt_str,this.io_writeback_22_bits_replay);
    pkt_str = $sformatf("%sio_writeback_22_bits_lqIdx_flag = 0x%0h ",pkt_str,this.io_writeback_22_bits_lqIdx_flag);
    pkt_str = $sformatf("%sio_writeback_22_bits_lqIdx_value = 0x%0h ",pkt_str,this.io_writeback_22_bits_lqIdx_value);
    pkt_str = $sformatf("%sio_writeback_22_bits_trigger = 0x%0h ",pkt_str,this.io_writeback_22_bits_trigger);
    pkt_str = $sformatf("%sio_writeback_22_bits_predecodeInfo_valid = 0x%0h ",pkt_str,this.io_writeback_22_bits_predecodeInfo_valid);
    pkt_str = $sformatf("%sio_writeback_22_bits_predecodeInfo_isRVC = 0x%0h ",pkt_str,this.io_writeback_22_bits_predecodeInfo_isRVC);
    pkt_str = $sformatf("%sio_writeback_22_bits_predecodeInfo_brType = 0x%0h ",pkt_str,this.io_writeback_22_bits_predecodeInfo_brType);
    pkt_str = $sformatf("%sio_writeback_22_bits_predecodeInfo_isCall = 0x%0h ",pkt_str,this.io_writeback_22_bits_predecodeInfo_isCall);
    pkt_str = $sformatf("%sio_writeback_22_bits_predecodeInfo_isRet = 0x%0h ",pkt_str,this.io_writeback_22_bits_predecodeInfo_isRet);
    pkt_str = $sformatf("%sio_writeback_22_bits_debug_isMMIO = 0x%0h ",pkt_str,this.io_writeback_22_bits_debug_isMMIO);
    pkt_str = $sformatf("%sio_writeback_22_bits_debug_isNCIO = 0x%0h ",pkt_str,this.io_writeback_22_bits_debug_isNCIO);
    pkt_str = $sformatf("%sio_writeback_22_bits_debug_isPerfCnt = 0x%0h ",pkt_str,this.io_writeback_22_bits_debug_isPerfCnt);
    pkt_str = $sformatf("%sio_writeback_22_bits_debug_paddr = 0x%0h ",pkt_str,this.io_writeback_22_bits_debug_paddr);
    pkt_str = $sformatf("%sio_writeback_22_bits_debug_vaddr = 0x%0h ",pkt_str,this.io_writeback_22_bits_debug_vaddr);
    pkt_str = $sformatf("%sio_writeback_22_bits_debugInfo_eliminatedMove = 0x%0h ",pkt_str,this.io_writeback_22_bits_debugInfo_eliminatedMove);
    pkt_str = $sformatf("%sio_writeback_22_bits_debugInfo_renameTime = 0x%0h ",pkt_str,this.io_writeback_22_bits_debugInfo_renameTime);
    pkt_str = $sformatf("%sio_writeback_22_bits_debugInfo_dispatchTime = 0x%0h ",pkt_str,this.io_writeback_22_bits_debugInfo_dispatchTime);
    pkt_str = $sformatf("%sio_writeback_22_bits_debugInfo_enqRsTime = 0x%0h ",pkt_str,this.io_writeback_22_bits_debugInfo_enqRsTime);
    pkt_str = $sformatf("%sio_writeback_22_bits_debugInfo_selectTime = 0x%0h ",pkt_str,this.io_writeback_22_bits_debugInfo_selectTime);
    pkt_str = $sformatf("%sio_writeback_22_bits_debugInfo_issueTime = 0x%0h ",pkt_str,this.io_writeback_22_bits_debugInfo_issueTime);
    pkt_str = $sformatf("%sio_writeback_22_bits_debugInfo_writebackTime = 0x%0h ",pkt_str,this.io_writeback_22_bits_debugInfo_writebackTime);
    pkt_str = $sformatf("%sio_writeback_22_bits_debugInfo_runahead_checkpoint_id = 0x%0h ",pkt_str,this.io_writeback_22_bits_debugInfo_runahead_checkpoint_id);
    pkt_str = $sformatf("%sio_writeback_22_bits_debugInfo_tlbFirstReqTime = 0x%0h ",pkt_str,this.io_writeback_22_bits_debugInfo_tlbFirstReqTime);
    pkt_str = $sformatf("%sio_writeback_22_bits_debugInfo_tlbRespTime = 0x%0h ",pkt_str,this.io_writeback_22_bits_debugInfo_tlbRespTime);
    pkt_str = $sformatf("%sio_writeback_22_bits_debug_seqNum = 0x%0h ",pkt_str,this.io_writeback_22_bits_debug_seqNum);
    pkt_str = $sformatf("%sio_writeback_21_valid = 0x%0h ",pkt_str,this.io_writeback_21_valid);
    pkt_str = $sformatf("%sio_writeback_21_bits_data_0 = 0x%0h ",pkt_str,this.io_writeback_21_bits_data_0);
    pkt_str = $sformatf("%sio_writeback_21_bits_pdest = 0x%0h ",pkt_str,this.io_writeback_21_bits_pdest);
    pkt_str = $sformatf("%sio_writeback_21_bits_robIdx_flag = 0x%0h ",pkt_str,this.io_writeback_21_bits_robIdx_flag);
    pkt_str = $sformatf("%sio_writeback_21_bits_robIdx_value = 0x%0h ",pkt_str,this.io_writeback_21_bits_robIdx_value);
    pkt_str = $sformatf("%sio_writeback_21_bits_intWen = 0x%0h ",pkt_str,this.io_writeback_21_bits_intWen);
    pkt_str = $sformatf("%sio_writeback_21_bits_fpWen = 0x%0h ",pkt_str,this.io_writeback_21_bits_fpWen);
    pkt_str = $sformatf("%sio_writeback_21_bits_exceptionVec_0 = 0x%0h ",pkt_str,this.io_writeback_21_bits_exceptionVec_0);
    pkt_str = $sformatf("%sio_writeback_21_bits_exceptionVec_1 = 0x%0h ",pkt_str,this.io_writeback_21_bits_exceptionVec_1);
    pkt_str = $sformatf("%sio_writeback_21_bits_exceptionVec_2 = 0x%0h ",pkt_str,this.io_writeback_21_bits_exceptionVec_2);
    pkt_str = $sformatf("%sio_writeback_21_bits_exceptionVec_3 = 0x%0h ",pkt_str,this.io_writeback_21_bits_exceptionVec_3);
    pkt_str = $sformatf("%sio_writeback_21_bits_exceptionVec_4 = 0x%0h ",pkt_str,this.io_writeback_21_bits_exceptionVec_4);
    pkt_str = $sformatf("%sio_writeback_21_bits_exceptionVec_5 = 0x%0h ",pkt_str,this.io_writeback_21_bits_exceptionVec_5);
    pkt_str = $sformatf("%sio_writeback_21_bits_exceptionVec_6 = 0x%0h ",pkt_str,this.io_writeback_21_bits_exceptionVec_6);
    pkt_str = $sformatf("%sio_writeback_21_bits_exceptionVec_7 = 0x%0h ",pkt_str,this.io_writeback_21_bits_exceptionVec_7);
    pkt_str = $sformatf("%sio_writeback_21_bits_exceptionVec_8 = 0x%0h ",pkt_str,this.io_writeback_21_bits_exceptionVec_8);
    pkt_str = $sformatf("%sio_writeback_21_bits_exceptionVec_9 = 0x%0h ",pkt_str,this.io_writeback_21_bits_exceptionVec_9);
    pkt_str = $sformatf("%sio_writeback_21_bits_exceptionVec_10 = 0x%0h ",pkt_str,this.io_writeback_21_bits_exceptionVec_10);
    pkt_str = $sformatf("%sio_writeback_21_bits_exceptionVec_11 = 0x%0h ",pkt_str,this.io_writeback_21_bits_exceptionVec_11);
    pkt_str = $sformatf("%sio_writeback_21_bits_exceptionVec_12 = 0x%0h ",pkt_str,this.io_writeback_21_bits_exceptionVec_12);
    pkt_str = $sformatf("%sio_writeback_21_bits_exceptionVec_13 = 0x%0h ",pkt_str,this.io_writeback_21_bits_exceptionVec_13);
    pkt_str = $sformatf("%sio_writeback_21_bits_exceptionVec_14 = 0x%0h ",pkt_str,this.io_writeback_21_bits_exceptionVec_14);
    pkt_str = $sformatf("%sio_writeback_21_bits_exceptionVec_15 = 0x%0h ",pkt_str,this.io_writeback_21_bits_exceptionVec_15);
    pkt_str = $sformatf("%sio_writeback_21_bits_exceptionVec_16 = 0x%0h ",pkt_str,this.io_writeback_21_bits_exceptionVec_16);
    pkt_str = $sformatf("%sio_writeback_21_bits_exceptionVec_17 = 0x%0h ",pkt_str,this.io_writeback_21_bits_exceptionVec_17);
    pkt_str = $sformatf("%sio_writeback_21_bits_exceptionVec_18 = 0x%0h ",pkt_str,this.io_writeback_21_bits_exceptionVec_18);
    pkt_str = $sformatf("%sio_writeback_21_bits_exceptionVec_19 = 0x%0h ",pkt_str,this.io_writeback_21_bits_exceptionVec_19);
    pkt_str = $sformatf("%sio_writeback_21_bits_exceptionVec_20 = 0x%0h ",pkt_str,this.io_writeback_21_bits_exceptionVec_20);
    pkt_str = $sformatf("%sio_writeback_21_bits_exceptionVec_21 = 0x%0h ",pkt_str,this.io_writeback_21_bits_exceptionVec_21);
    pkt_str = $sformatf("%sio_writeback_21_bits_exceptionVec_22 = 0x%0h ",pkt_str,this.io_writeback_21_bits_exceptionVec_22);
    pkt_str = $sformatf("%sio_writeback_21_bits_exceptionVec_23 = 0x%0h ",pkt_str,this.io_writeback_21_bits_exceptionVec_23);
    pkt_str = $sformatf("%sio_writeback_21_bits_flushPipe = 0x%0h ",pkt_str,this.io_writeback_21_bits_flushPipe);
    pkt_str = $sformatf("%sio_writeback_21_bits_replay = 0x%0h ",pkt_str,this.io_writeback_21_bits_replay);
    pkt_str = $sformatf("%sio_writeback_21_bits_lqIdx_flag = 0x%0h ",pkt_str,this.io_writeback_21_bits_lqIdx_flag);
    pkt_str = $sformatf("%sio_writeback_21_bits_lqIdx_value = 0x%0h ",pkt_str,this.io_writeback_21_bits_lqIdx_value);
    pkt_str = $sformatf("%sio_writeback_21_bits_trigger = 0x%0h ",pkt_str,this.io_writeback_21_bits_trigger);
    pkt_str = $sformatf("%sio_writeback_21_bits_predecodeInfo_valid = 0x%0h ",pkt_str,this.io_writeback_21_bits_predecodeInfo_valid);
    pkt_str = $sformatf("%sio_writeback_21_bits_predecodeInfo_isRVC = 0x%0h ",pkt_str,this.io_writeback_21_bits_predecodeInfo_isRVC);
    pkt_str = $sformatf("%sio_writeback_21_bits_predecodeInfo_brType = 0x%0h ",pkt_str,this.io_writeback_21_bits_predecodeInfo_brType);
    pkt_str = $sformatf("%sio_writeback_21_bits_predecodeInfo_isCall = 0x%0h ",pkt_str,this.io_writeback_21_bits_predecodeInfo_isCall);
    pkt_str = $sformatf("%sio_writeback_21_bits_predecodeInfo_isRet = 0x%0h ",pkt_str,this.io_writeback_21_bits_predecodeInfo_isRet);
    pkt_str = $sformatf("%sio_writeback_21_bits_debug_isMMIO = 0x%0h ",pkt_str,this.io_writeback_21_bits_debug_isMMIO);
    pkt_str = $sformatf("%sio_writeback_21_bits_debug_isNCIO = 0x%0h ",pkt_str,this.io_writeback_21_bits_debug_isNCIO);
    pkt_str = $sformatf("%sio_writeback_21_bits_debug_isPerfCnt = 0x%0h ",pkt_str,this.io_writeback_21_bits_debug_isPerfCnt);
    pkt_str = $sformatf("%sio_writeback_21_bits_debug_paddr = 0x%0h ",pkt_str,this.io_writeback_21_bits_debug_paddr);
    pkt_str = $sformatf("%sio_writeback_21_bits_debug_vaddr = 0x%0h ",pkt_str,this.io_writeback_21_bits_debug_vaddr);
    pkt_str = $sformatf("%sio_writeback_21_bits_debugInfo_eliminatedMove = 0x%0h ",pkt_str,this.io_writeback_21_bits_debugInfo_eliminatedMove);
    pkt_str = $sformatf("%sio_writeback_21_bits_debugInfo_renameTime = 0x%0h ",pkt_str,this.io_writeback_21_bits_debugInfo_renameTime);
    pkt_str = $sformatf("%sio_writeback_21_bits_debugInfo_dispatchTime = 0x%0h ",pkt_str,this.io_writeback_21_bits_debugInfo_dispatchTime);
    pkt_str = $sformatf("%sio_writeback_21_bits_debugInfo_enqRsTime = 0x%0h ",pkt_str,this.io_writeback_21_bits_debugInfo_enqRsTime);
    pkt_str = $sformatf("%sio_writeback_21_bits_debugInfo_selectTime = 0x%0h ",pkt_str,this.io_writeback_21_bits_debugInfo_selectTime);
    pkt_str = $sformatf("%sio_writeback_21_bits_debugInfo_issueTime = 0x%0h ",pkt_str,this.io_writeback_21_bits_debugInfo_issueTime);
    pkt_str = $sformatf("%sio_writeback_21_bits_debugInfo_writebackTime = 0x%0h ",pkt_str,this.io_writeback_21_bits_debugInfo_writebackTime);
    pkt_str = $sformatf("%sio_writeback_21_bits_debugInfo_runahead_checkpoint_id = 0x%0h ",pkt_str,this.io_writeback_21_bits_debugInfo_runahead_checkpoint_id);
    pkt_str = $sformatf("%sio_writeback_21_bits_debugInfo_tlbFirstReqTime = 0x%0h ",pkt_str,this.io_writeback_21_bits_debugInfo_tlbFirstReqTime);
    pkt_str = $sformatf("%sio_writeback_21_bits_debugInfo_tlbRespTime = 0x%0h ",pkt_str,this.io_writeback_21_bits_debugInfo_tlbRespTime);
    pkt_str = $sformatf("%sio_writeback_21_bits_debug_seqNum = 0x%0h ",pkt_str,this.io_writeback_21_bits_debug_seqNum);
    pkt_str = $sformatf("%sio_writeback_20_valid = 0x%0h ",pkt_str,this.io_writeback_20_valid);
    pkt_str = $sformatf("%sio_writeback_20_bits_data_0 = 0x%0h ",pkt_str,this.io_writeback_20_bits_data_0);
    pkt_str = $sformatf("%sio_writeback_20_bits_pdest = 0x%0h ",pkt_str,this.io_writeback_20_bits_pdest);
    pkt_str = $sformatf("%sio_writeback_20_bits_robIdx_flag = 0x%0h ",pkt_str,this.io_writeback_20_bits_robIdx_flag);
    pkt_str = $sformatf("%sio_writeback_20_bits_robIdx_value = 0x%0h ",pkt_str,this.io_writeback_20_bits_robIdx_value);
    pkt_str = $sformatf("%sio_writeback_20_bits_intWen = 0x%0h ",pkt_str,this.io_writeback_20_bits_intWen);
    pkt_str = $sformatf("%sio_writeback_20_bits_fpWen = 0x%0h ",pkt_str,this.io_writeback_20_bits_fpWen);
    pkt_str = $sformatf("%sio_writeback_20_bits_exceptionVec_0 = 0x%0h ",pkt_str,this.io_writeback_20_bits_exceptionVec_0);
    pkt_str = $sformatf("%sio_writeback_20_bits_exceptionVec_1 = 0x%0h ",pkt_str,this.io_writeback_20_bits_exceptionVec_1);
    pkt_str = $sformatf("%sio_writeback_20_bits_exceptionVec_2 = 0x%0h ",pkt_str,this.io_writeback_20_bits_exceptionVec_2);
    pkt_str = $sformatf("%sio_writeback_20_bits_exceptionVec_3 = 0x%0h ",pkt_str,this.io_writeback_20_bits_exceptionVec_3);
    pkt_str = $sformatf("%sio_writeback_20_bits_exceptionVec_4 = 0x%0h ",pkt_str,this.io_writeback_20_bits_exceptionVec_4);
    pkt_str = $sformatf("%sio_writeback_20_bits_exceptionVec_5 = 0x%0h ",pkt_str,this.io_writeback_20_bits_exceptionVec_5);
    pkt_str = $sformatf("%sio_writeback_20_bits_exceptionVec_6 = 0x%0h ",pkt_str,this.io_writeback_20_bits_exceptionVec_6);
    pkt_str = $sformatf("%sio_writeback_20_bits_exceptionVec_7 = 0x%0h ",pkt_str,this.io_writeback_20_bits_exceptionVec_7);
    pkt_str = $sformatf("%sio_writeback_20_bits_exceptionVec_8 = 0x%0h ",pkt_str,this.io_writeback_20_bits_exceptionVec_8);
    pkt_str = $sformatf("%sio_writeback_20_bits_exceptionVec_9 = 0x%0h ",pkt_str,this.io_writeback_20_bits_exceptionVec_9);
    pkt_str = $sformatf("%sio_writeback_20_bits_exceptionVec_10 = 0x%0h ",pkt_str,this.io_writeback_20_bits_exceptionVec_10);
    pkt_str = $sformatf("%sio_writeback_20_bits_exceptionVec_11 = 0x%0h ",pkt_str,this.io_writeback_20_bits_exceptionVec_11);
    pkt_str = $sformatf("%sio_writeback_20_bits_exceptionVec_12 = 0x%0h ",pkt_str,this.io_writeback_20_bits_exceptionVec_12);
    pkt_str = $sformatf("%sio_writeback_20_bits_exceptionVec_13 = 0x%0h ",pkt_str,this.io_writeback_20_bits_exceptionVec_13);
    pkt_str = $sformatf("%sio_writeback_20_bits_exceptionVec_14 = 0x%0h ",pkt_str,this.io_writeback_20_bits_exceptionVec_14);
    pkt_str = $sformatf("%sio_writeback_20_bits_exceptionVec_15 = 0x%0h ",pkt_str,this.io_writeback_20_bits_exceptionVec_15);
    pkt_str = $sformatf("%sio_writeback_20_bits_exceptionVec_16 = 0x%0h ",pkt_str,this.io_writeback_20_bits_exceptionVec_16);
    pkt_str = $sformatf("%sio_writeback_20_bits_exceptionVec_17 = 0x%0h ",pkt_str,this.io_writeback_20_bits_exceptionVec_17);
    pkt_str = $sformatf("%sio_writeback_20_bits_exceptionVec_18 = 0x%0h ",pkt_str,this.io_writeback_20_bits_exceptionVec_18);
    pkt_str = $sformatf("%sio_writeback_20_bits_exceptionVec_19 = 0x%0h ",pkt_str,this.io_writeback_20_bits_exceptionVec_19);
    pkt_str = $sformatf("%sio_writeback_20_bits_exceptionVec_20 = 0x%0h ",pkt_str,this.io_writeback_20_bits_exceptionVec_20);
    pkt_str = $sformatf("%sio_writeback_20_bits_exceptionVec_21 = 0x%0h ",pkt_str,this.io_writeback_20_bits_exceptionVec_21);
    pkt_str = $sformatf("%sio_writeback_20_bits_exceptionVec_22 = 0x%0h ",pkt_str,this.io_writeback_20_bits_exceptionVec_22);
    pkt_str = $sformatf("%sio_writeback_20_bits_exceptionVec_23 = 0x%0h ",pkt_str,this.io_writeback_20_bits_exceptionVec_23);
    pkt_str = $sformatf("%sio_writeback_20_bits_flushPipe = 0x%0h ",pkt_str,this.io_writeback_20_bits_flushPipe);
    pkt_str = $sformatf("%sio_writeback_20_bits_replay = 0x%0h ",pkt_str,this.io_writeback_20_bits_replay);
    pkt_str = $sformatf("%sio_writeback_20_bits_lqIdx_flag = 0x%0h ",pkt_str,this.io_writeback_20_bits_lqIdx_flag);
    pkt_str = $sformatf("%sio_writeback_20_bits_lqIdx_value = 0x%0h ",pkt_str,this.io_writeback_20_bits_lqIdx_value);
    pkt_str = $sformatf("%sio_writeback_20_bits_trigger = 0x%0h ",pkt_str,this.io_writeback_20_bits_trigger);
    pkt_str = $sformatf("%sio_writeback_20_bits_predecodeInfo_valid = 0x%0h ",pkt_str,this.io_writeback_20_bits_predecodeInfo_valid);
    pkt_str = $sformatf("%sio_writeback_20_bits_predecodeInfo_isRVC = 0x%0h ",pkt_str,this.io_writeback_20_bits_predecodeInfo_isRVC);
    pkt_str = $sformatf("%sio_writeback_20_bits_predecodeInfo_brType = 0x%0h ",pkt_str,this.io_writeback_20_bits_predecodeInfo_brType);
    pkt_str = $sformatf("%sio_writeback_20_bits_predecodeInfo_isCall = 0x%0h ",pkt_str,this.io_writeback_20_bits_predecodeInfo_isCall);
    pkt_str = $sformatf("%sio_writeback_20_bits_predecodeInfo_isRet = 0x%0h ",pkt_str,this.io_writeback_20_bits_predecodeInfo_isRet);
    pkt_str = $sformatf("%sio_writeback_20_bits_debug_isMMIO = 0x%0h ",pkt_str,this.io_writeback_20_bits_debug_isMMIO);
    pkt_str = $sformatf("%sio_writeback_20_bits_debug_isNCIO = 0x%0h ",pkt_str,this.io_writeback_20_bits_debug_isNCIO);
    pkt_str = $sformatf("%sio_writeback_20_bits_debug_isPerfCnt = 0x%0h ",pkt_str,this.io_writeback_20_bits_debug_isPerfCnt);
    pkt_str = $sformatf("%sio_writeback_20_bits_debug_paddr = 0x%0h ",pkt_str,this.io_writeback_20_bits_debug_paddr);
    pkt_str = $sformatf("%sio_writeback_20_bits_debug_vaddr = 0x%0h ",pkt_str,this.io_writeback_20_bits_debug_vaddr);
    pkt_str = $sformatf("%sio_writeback_20_bits_debugInfo_eliminatedMove = 0x%0h ",pkt_str,this.io_writeback_20_bits_debugInfo_eliminatedMove);
    pkt_str = $sformatf("%sio_writeback_20_bits_debugInfo_renameTime = 0x%0h ",pkt_str,this.io_writeback_20_bits_debugInfo_renameTime);
    pkt_str = $sformatf("%sio_writeback_20_bits_debugInfo_dispatchTime = 0x%0h ",pkt_str,this.io_writeback_20_bits_debugInfo_dispatchTime);
    pkt_str = $sformatf("%sio_writeback_20_bits_debugInfo_enqRsTime = 0x%0h ",pkt_str,this.io_writeback_20_bits_debugInfo_enqRsTime);
    pkt_str = $sformatf("%sio_writeback_20_bits_debugInfo_selectTime = 0x%0h ",pkt_str,this.io_writeback_20_bits_debugInfo_selectTime);
    pkt_str = $sformatf("%sio_writeback_20_bits_debugInfo_issueTime = 0x%0h ",pkt_str,this.io_writeback_20_bits_debugInfo_issueTime);
    pkt_str = $sformatf("%sio_writeback_20_bits_debugInfo_writebackTime = 0x%0h ",pkt_str,this.io_writeback_20_bits_debugInfo_writebackTime);
    pkt_str = $sformatf("%sio_writeback_20_bits_debugInfo_runahead_checkpoint_id = 0x%0h ",pkt_str,this.io_writeback_20_bits_debugInfo_runahead_checkpoint_id);
    pkt_str = $sformatf("%sio_writeback_20_bits_debugInfo_tlbFirstReqTime = 0x%0h ",pkt_str,this.io_writeback_20_bits_debugInfo_tlbFirstReqTime);
    pkt_str = $sformatf("%sio_writeback_20_bits_debugInfo_tlbRespTime = 0x%0h ",pkt_str,this.io_writeback_20_bits_debugInfo_tlbRespTime);
    pkt_str = $sformatf("%sio_writeback_20_bits_debug_seqNum = 0x%0h ",pkt_str,this.io_writeback_20_bits_debug_seqNum);
    pkt_str = $sformatf("%sio_writeback_19_valid = 0x%0h ",pkt_str,this.io_writeback_19_valid);
    pkt_str = $sformatf("%sio_writeback_19_bits_data_0 = 0x%0h ",pkt_str,this.io_writeback_19_bits_data_0);
    pkt_str = $sformatf("%sio_writeback_19_bits_pdest = 0x%0h ",pkt_str,this.io_writeback_19_bits_pdest);
    pkt_str = $sformatf("%sio_writeback_19_bits_robIdx_flag = 0x%0h ",pkt_str,this.io_writeback_19_bits_robIdx_flag);
    pkt_str = $sformatf("%sio_writeback_19_bits_robIdx_value = 0x%0h ",pkt_str,this.io_writeback_19_bits_robIdx_value);
    pkt_str = $sformatf("%sio_writeback_19_bits_intWen = 0x%0h ",pkt_str,this.io_writeback_19_bits_intWen);
    pkt_str = $sformatf("%sio_writeback_19_bits_exceptionVec_0 = 0x%0h ",pkt_str,this.io_writeback_19_bits_exceptionVec_0);
    pkt_str = $sformatf("%sio_writeback_19_bits_exceptionVec_1 = 0x%0h ",pkt_str,this.io_writeback_19_bits_exceptionVec_1);
    pkt_str = $sformatf("%sio_writeback_19_bits_exceptionVec_2 = 0x%0h ",pkt_str,this.io_writeback_19_bits_exceptionVec_2);
    pkt_str = $sformatf("%sio_writeback_19_bits_exceptionVec_3 = 0x%0h ",pkt_str,this.io_writeback_19_bits_exceptionVec_3);
    pkt_str = $sformatf("%sio_writeback_19_bits_exceptionVec_4 = 0x%0h ",pkt_str,this.io_writeback_19_bits_exceptionVec_4);
    pkt_str = $sformatf("%sio_writeback_19_bits_exceptionVec_5 = 0x%0h ",pkt_str,this.io_writeback_19_bits_exceptionVec_5);
    pkt_str = $sformatf("%sio_writeback_19_bits_exceptionVec_6 = 0x%0h ",pkt_str,this.io_writeback_19_bits_exceptionVec_6);
    pkt_str = $sformatf("%sio_writeback_19_bits_exceptionVec_7 = 0x%0h ",pkt_str,this.io_writeback_19_bits_exceptionVec_7);
    pkt_str = $sformatf("%sio_writeback_19_bits_exceptionVec_8 = 0x%0h ",pkt_str,this.io_writeback_19_bits_exceptionVec_8);
    pkt_str = $sformatf("%sio_writeback_19_bits_exceptionVec_9 = 0x%0h ",pkt_str,this.io_writeback_19_bits_exceptionVec_9);
    pkt_str = $sformatf("%sio_writeback_19_bits_exceptionVec_10 = 0x%0h ",pkt_str,this.io_writeback_19_bits_exceptionVec_10);
    pkt_str = $sformatf("%sio_writeback_19_bits_exceptionVec_11 = 0x%0h ",pkt_str,this.io_writeback_19_bits_exceptionVec_11);
    pkt_str = $sformatf("%sio_writeback_19_bits_exceptionVec_12 = 0x%0h ",pkt_str,this.io_writeback_19_bits_exceptionVec_12);
    pkt_str = $sformatf("%sio_writeback_19_bits_exceptionVec_13 = 0x%0h ",pkt_str,this.io_writeback_19_bits_exceptionVec_13);
    pkt_str = $sformatf("%sio_writeback_19_bits_exceptionVec_14 = 0x%0h ",pkt_str,this.io_writeback_19_bits_exceptionVec_14);
    pkt_str = $sformatf("%sio_writeback_19_bits_exceptionVec_15 = 0x%0h ",pkt_str,this.io_writeback_19_bits_exceptionVec_15);
    pkt_str = $sformatf("%sio_writeback_19_bits_exceptionVec_16 = 0x%0h ",pkt_str,this.io_writeback_19_bits_exceptionVec_16);
    pkt_str = $sformatf("%sio_writeback_19_bits_exceptionVec_17 = 0x%0h ",pkt_str,this.io_writeback_19_bits_exceptionVec_17);
    pkt_str = $sformatf("%sio_writeback_19_bits_exceptionVec_18 = 0x%0h ",pkt_str,this.io_writeback_19_bits_exceptionVec_18);
    pkt_str = $sformatf("%sio_writeback_19_bits_exceptionVec_19 = 0x%0h ",pkt_str,this.io_writeback_19_bits_exceptionVec_19);
    pkt_str = $sformatf("%sio_writeback_19_bits_exceptionVec_20 = 0x%0h ",pkt_str,this.io_writeback_19_bits_exceptionVec_20);
    pkt_str = $sformatf("%sio_writeback_19_bits_exceptionVec_21 = 0x%0h ",pkt_str,this.io_writeback_19_bits_exceptionVec_21);
    pkt_str = $sformatf("%sio_writeback_19_bits_exceptionVec_22 = 0x%0h ",pkt_str,this.io_writeback_19_bits_exceptionVec_22);
    pkt_str = $sformatf("%sio_writeback_19_bits_exceptionVec_23 = 0x%0h ",pkt_str,this.io_writeback_19_bits_exceptionVec_23);
    pkt_str = $sformatf("%sio_writeback_19_bits_flushPipe = 0x%0h ",pkt_str,this.io_writeback_19_bits_flushPipe);
    pkt_str = $sformatf("%sio_writeback_19_bits_sqIdx_flag = 0x%0h ",pkt_str,this.io_writeback_19_bits_sqIdx_flag);
    pkt_str = $sformatf("%sio_writeback_19_bits_sqIdx_value = 0x%0h ",pkt_str,this.io_writeback_19_bits_sqIdx_value);
    pkt_str = $sformatf("%sio_writeback_19_bits_trigger = 0x%0h ",pkt_str,this.io_writeback_19_bits_trigger);
    pkt_str = $sformatf("%sio_writeback_19_bits_debug_isMMIO = 0x%0h ",pkt_str,this.io_writeback_19_bits_debug_isMMIO);
    pkt_str = $sformatf("%sio_writeback_19_bits_debug_isNCIO = 0x%0h ",pkt_str,this.io_writeback_19_bits_debug_isNCIO);
    pkt_str = $sformatf("%sio_writeback_19_bits_debug_isPerfCnt = 0x%0h ",pkt_str,this.io_writeback_19_bits_debug_isPerfCnt);
    pkt_str = $sformatf("%sio_writeback_19_bits_debug_paddr = 0x%0h ",pkt_str,this.io_writeback_19_bits_debug_paddr);
    pkt_str = $sformatf("%sio_writeback_19_bits_debug_vaddr = 0x%0h ",pkt_str,this.io_writeback_19_bits_debug_vaddr);
    pkt_str = $sformatf("%sio_writeback_19_bits_debugInfo_eliminatedMove = 0x%0h ",pkt_str,this.io_writeback_19_bits_debugInfo_eliminatedMove);
    pkt_str = $sformatf("%sio_writeback_19_bits_debugInfo_renameTime = 0x%0h ",pkt_str,this.io_writeback_19_bits_debugInfo_renameTime);
    pkt_str = $sformatf("%sio_writeback_19_bits_debugInfo_dispatchTime = 0x%0h ",pkt_str,this.io_writeback_19_bits_debugInfo_dispatchTime);
    pkt_str = $sformatf("%sio_writeback_19_bits_debugInfo_enqRsTime = 0x%0h ",pkt_str,this.io_writeback_19_bits_debugInfo_enqRsTime);
    pkt_str = $sformatf("%sio_writeback_19_bits_debugInfo_selectTime = 0x%0h ",pkt_str,this.io_writeback_19_bits_debugInfo_selectTime);
    pkt_str = $sformatf("%sio_writeback_19_bits_debugInfo_issueTime = 0x%0h ",pkt_str,this.io_writeback_19_bits_debugInfo_issueTime);
    pkt_str = $sformatf("%sio_writeback_19_bits_debugInfo_writebackTime = 0x%0h ",pkt_str,this.io_writeback_19_bits_debugInfo_writebackTime);
    pkt_str = $sformatf("%sio_writeback_19_bits_debugInfo_runahead_checkpoint_id = 0x%0h ",pkt_str,this.io_writeback_19_bits_debugInfo_runahead_checkpoint_id);
    pkt_str = $sformatf("%sio_writeback_19_bits_debugInfo_tlbFirstReqTime = 0x%0h ",pkt_str,this.io_writeback_19_bits_debugInfo_tlbFirstReqTime);
    pkt_str = $sformatf("%sio_writeback_19_bits_debugInfo_tlbRespTime = 0x%0h ",pkt_str,this.io_writeback_19_bits_debugInfo_tlbRespTime);
    pkt_str = $sformatf("%sio_writeback_19_bits_debug_seqNum = 0x%0h ",pkt_str,this.io_writeback_19_bits_debug_seqNum);
    pkt_str = $sformatf("%sio_writeback_18_valid = 0x%0h ",pkt_str,this.io_writeback_18_valid);
    pkt_str = $sformatf("%sio_writeback_18_bits_data_0 = 0x%0h ",pkt_str,this.io_writeback_18_bits_data_0);
    pkt_str = $sformatf("%sio_writeback_18_bits_pdest = 0x%0h ",pkt_str,this.io_writeback_18_bits_pdest);
    pkt_str = $sformatf("%sio_writeback_18_bits_robIdx_flag = 0x%0h ",pkt_str,this.io_writeback_18_bits_robIdx_flag);
    pkt_str = $sformatf("%sio_writeback_18_bits_robIdx_value = 0x%0h ",pkt_str,this.io_writeback_18_bits_robIdx_value);
    pkt_str = $sformatf("%sio_writeback_18_bits_intWen = 0x%0h ",pkt_str,this.io_writeback_18_bits_intWen);
    pkt_str = $sformatf("%sio_writeback_18_bits_exceptionVec_0 = 0x%0h ",pkt_str,this.io_writeback_18_bits_exceptionVec_0);
    pkt_str = $sformatf("%sio_writeback_18_bits_exceptionVec_1 = 0x%0h ",pkt_str,this.io_writeback_18_bits_exceptionVec_1);
    pkt_str = $sformatf("%sio_writeback_18_bits_exceptionVec_2 = 0x%0h ",pkt_str,this.io_writeback_18_bits_exceptionVec_2);
    pkt_str = $sformatf("%sio_writeback_18_bits_exceptionVec_3 = 0x%0h ",pkt_str,this.io_writeback_18_bits_exceptionVec_3);
    pkt_str = $sformatf("%sio_writeback_18_bits_exceptionVec_4 = 0x%0h ",pkt_str,this.io_writeback_18_bits_exceptionVec_4);
    pkt_str = $sformatf("%sio_writeback_18_bits_exceptionVec_5 = 0x%0h ",pkt_str,this.io_writeback_18_bits_exceptionVec_5);
    pkt_str = $sformatf("%sio_writeback_18_bits_exceptionVec_6 = 0x%0h ",pkt_str,this.io_writeback_18_bits_exceptionVec_6);
    pkt_str = $sformatf("%sio_writeback_18_bits_exceptionVec_7 = 0x%0h ",pkt_str,this.io_writeback_18_bits_exceptionVec_7);
    pkt_str = $sformatf("%sio_writeback_18_bits_exceptionVec_8 = 0x%0h ",pkt_str,this.io_writeback_18_bits_exceptionVec_8);
    pkt_str = $sformatf("%sio_writeback_18_bits_exceptionVec_9 = 0x%0h ",pkt_str,this.io_writeback_18_bits_exceptionVec_9);
    pkt_str = $sformatf("%sio_writeback_18_bits_exceptionVec_10 = 0x%0h ",pkt_str,this.io_writeback_18_bits_exceptionVec_10);
    pkt_str = $sformatf("%sio_writeback_18_bits_exceptionVec_11 = 0x%0h ",pkt_str,this.io_writeback_18_bits_exceptionVec_11);
    pkt_str = $sformatf("%sio_writeback_18_bits_exceptionVec_12 = 0x%0h ",pkt_str,this.io_writeback_18_bits_exceptionVec_12);
    pkt_str = $sformatf("%sio_writeback_18_bits_exceptionVec_13 = 0x%0h ",pkt_str,this.io_writeback_18_bits_exceptionVec_13);
    pkt_str = $sformatf("%sio_writeback_18_bits_exceptionVec_14 = 0x%0h ",pkt_str,this.io_writeback_18_bits_exceptionVec_14);
    pkt_str = $sformatf("%sio_writeback_18_bits_exceptionVec_15 = 0x%0h ",pkt_str,this.io_writeback_18_bits_exceptionVec_15);
    pkt_str = $sformatf("%sio_writeback_18_bits_exceptionVec_16 = 0x%0h ",pkt_str,this.io_writeback_18_bits_exceptionVec_16);
    pkt_str = $sformatf("%sio_writeback_18_bits_exceptionVec_17 = 0x%0h ",pkt_str,this.io_writeback_18_bits_exceptionVec_17);
    pkt_str = $sformatf("%sio_writeback_18_bits_exceptionVec_18 = 0x%0h ",pkt_str,this.io_writeback_18_bits_exceptionVec_18);
    pkt_str = $sformatf("%sio_writeback_18_bits_exceptionVec_19 = 0x%0h ",pkt_str,this.io_writeback_18_bits_exceptionVec_19);
    pkt_str = $sformatf("%sio_writeback_18_bits_exceptionVec_20 = 0x%0h ",pkt_str,this.io_writeback_18_bits_exceptionVec_20);
    pkt_str = $sformatf("%sio_writeback_18_bits_exceptionVec_21 = 0x%0h ",pkt_str,this.io_writeback_18_bits_exceptionVec_21);
    pkt_str = $sformatf("%sio_writeback_18_bits_exceptionVec_22 = 0x%0h ",pkt_str,this.io_writeback_18_bits_exceptionVec_22);
    pkt_str = $sformatf("%sio_writeback_18_bits_exceptionVec_23 = 0x%0h ",pkt_str,this.io_writeback_18_bits_exceptionVec_23);
    pkt_str = $sformatf("%sio_writeback_18_bits_flushPipe = 0x%0h ",pkt_str,this.io_writeback_18_bits_flushPipe);
    pkt_str = $sformatf("%sio_writeback_18_bits_sqIdx_flag = 0x%0h ",pkt_str,this.io_writeback_18_bits_sqIdx_flag);
    pkt_str = $sformatf("%sio_writeback_18_bits_sqIdx_value = 0x%0h ",pkt_str,this.io_writeback_18_bits_sqIdx_value);
    pkt_str = $sformatf("%sio_writeback_18_bits_trigger = 0x%0h ",pkt_str,this.io_writeback_18_bits_trigger);
    pkt_str = $sformatf("%sio_writeback_18_bits_debug_isMMIO = 0x%0h ",pkt_str,this.io_writeback_18_bits_debug_isMMIO);
    pkt_str = $sformatf("%sio_writeback_18_bits_debug_isNCIO = 0x%0h ",pkt_str,this.io_writeback_18_bits_debug_isNCIO);
    pkt_str = $sformatf("%sio_writeback_18_bits_debug_isPerfCnt = 0x%0h ",pkt_str,this.io_writeback_18_bits_debug_isPerfCnt);
    pkt_str = $sformatf("%sio_writeback_18_bits_debug_paddr = 0x%0h ",pkt_str,this.io_writeback_18_bits_debug_paddr);
    pkt_str = $sformatf("%sio_writeback_18_bits_debug_vaddr = 0x%0h ",pkt_str,this.io_writeback_18_bits_debug_vaddr);
    pkt_str = $sformatf("%sio_writeback_18_bits_debugInfo_eliminatedMove = 0x%0h ",pkt_str,this.io_writeback_18_bits_debugInfo_eliminatedMove);
    pkt_str = $sformatf("%sio_writeback_18_bits_debugInfo_renameTime = 0x%0h ",pkt_str,this.io_writeback_18_bits_debugInfo_renameTime);
    pkt_str = $sformatf("%sio_writeback_18_bits_debugInfo_dispatchTime = 0x%0h ",pkt_str,this.io_writeback_18_bits_debugInfo_dispatchTime);
    pkt_str = $sformatf("%sio_writeback_18_bits_debugInfo_enqRsTime = 0x%0h ",pkt_str,this.io_writeback_18_bits_debugInfo_enqRsTime);
    pkt_str = $sformatf("%sio_writeback_18_bits_debugInfo_selectTime = 0x%0h ",pkt_str,this.io_writeback_18_bits_debugInfo_selectTime);
    pkt_str = $sformatf("%sio_writeback_18_bits_debugInfo_issueTime = 0x%0h ",pkt_str,this.io_writeback_18_bits_debugInfo_issueTime);
    pkt_str = $sformatf("%sio_writeback_18_bits_debugInfo_writebackTime = 0x%0h ",pkt_str,this.io_writeback_18_bits_debugInfo_writebackTime);
    pkt_str = $sformatf("%sio_writeback_18_bits_debugInfo_runahead_checkpoint_id = 0x%0h ",pkt_str,this.io_writeback_18_bits_debugInfo_runahead_checkpoint_id);
    pkt_str = $sformatf("%sio_writeback_18_bits_debugInfo_tlbFirstReqTime = 0x%0h ",pkt_str,this.io_writeback_18_bits_debugInfo_tlbFirstReqTime);
    pkt_str = $sformatf("%sio_writeback_18_bits_debugInfo_tlbRespTime = 0x%0h ",pkt_str,this.io_writeback_18_bits_debugInfo_tlbRespTime);
    pkt_str = $sformatf("%sio_writeback_18_bits_debug_seqNum = 0x%0h ",pkt_str,this.io_writeback_18_bits_debug_seqNum);
    pkt_str = $sformatf("%sio_writeback_17_valid = 0x%0h ",pkt_str,this.io_writeback_17_valid);
    pkt_str = $sformatf("%sio_writeback_17_bits_data_0 = 0x%0h ",pkt_str,this.io_writeback_17_bits_data_0);
    pkt_str = $sformatf("%sio_writeback_17_bits_data_1 = 0x%0h ",pkt_str,this.io_writeback_17_bits_data_1);
    pkt_str = $sformatf("%sio_writeback_17_bits_data_2 = 0x%0h ",pkt_str,this.io_writeback_17_bits_data_2);
    pkt_str = $sformatf("%sio_writeback_17_bits_pdest = 0x%0h ",pkt_str,this.io_writeback_17_bits_pdest);
    pkt_str = $sformatf("%sio_writeback_17_bits_robIdx_flag = 0x%0h ",pkt_str,this.io_writeback_17_bits_robIdx_flag);
    pkt_str = $sformatf("%sio_writeback_17_bits_robIdx_value = 0x%0h ",pkt_str,this.io_writeback_17_bits_robIdx_value);
    pkt_str = $sformatf("%sio_writeback_17_bits_vecWen = 0x%0h ",pkt_str,this.io_writeback_17_bits_vecWen);
    pkt_str = $sformatf("%sio_writeback_17_bits_v0Wen = 0x%0h ",pkt_str,this.io_writeback_17_bits_v0Wen);
    pkt_str = $sformatf("%sio_writeback_17_bits_fflags = 0x%0h ",pkt_str,this.io_writeback_17_bits_fflags);
    pkt_str = $sformatf("%sio_writeback_17_bits_wflags = 0x%0h ",pkt_str,this.io_writeback_17_bits_wflags);
    pkt_str = $sformatf("%sio_writeback_17_bits_debugInfo_eliminatedMove = 0x%0h ",pkt_str,this.io_writeback_17_bits_debugInfo_eliminatedMove);
    pkt_str = $sformatf("%sio_writeback_17_bits_debugInfo_renameTime = 0x%0h ",pkt_str,this.io_writeback_17_bits_debugInfo_renameTime);
    pkt_str = $sformatf("%sio_writeback_17_bits_debugInfo_dispatchTime = 0x%0h ",pkt_str,this.io_writeback_17_bits_debugInfo_dispatchTime);
    pkt_str = $sformatf("%sio_writeback_17_bits_debugInfo_enqRsTime = 0x%0h ",pkt_str,this.io_writeback_17_bits_debugInfo_enqRsTime);
    pkt_str = $sformatf("%sio_writeback_17_bits_debugInfo_selectTime = 0x%0h ",pkt_str,this.io_writeback_17_bits_debugInfo_selectTime);
    pkt_str = $sformatf("%sio_writeback_17_bits_debugInfo_issueTime = 0x%0h ",pkt_str,this.io_writeback_17_bits_debugInfo_issueTime);
    pkt_str = $sformatf("%sio_writeback_17_bits_debugInfo_writebackTime = 0x%0h ",pkt_str,this.io_writeback_17_bits_debugInfo_writebackTime);
    pkt_str = $sformatf("%sio_writeback_17_bits_debugInfo_runahead_checkpoint_id = 0x%0h ",pkt_str,this.io_writeback_17_bits_debugInfo_runahead_checkpoint_id);
    pkt_str = $sformatf("%sio_writeback_17_bits_debugInfo_tlbFirstReqTime = 0x%0h ",pkt_str,this.io_writeback_17_bits_debugInfo_tlbFirstReqTime);
    pkt_str = $sformatf("%sio_writeback_17_bits_debugInfo_tlbRespTime = 0x%0h ",pkt_str,this.io_writeback_17_bits_debugInfo_tlbRespTime);
    pkt_str = $sformatf("%sio_writeback_17_bits_debug_seqNum = 0x%0h ",pkt_str,this.io_writeback_17_bits_debug_seqNum);
    pkt_str = $sformatf("%sio_writeback_16_valid = 0x%0h ",pkt_str,this.io_writeback_16_valid);
    pkt_str = $sformatf("%sio_writeback_16_bits_data_0 = 0x%0h ",pkt_str,this.io_writeback_16_bits_data_0);
    pkt_str = $sformatf("%sio_writeback_16_bits_data_1 = 0x%0h ",pkt_str,this.io_writeback_16_bits_data_1);
    pkt_str = $sformatf("%sio_writeback_16_bits_data_2 = 0x%0h ",pkt_str,this.io_writeback_16_bits_data_2);
    pkt_str = $sformatf("%sio_writeback_16_bits_data_3 = 0x%0h ",pkt_str,this.io_writeback_16_bits_data_3);
    pkt_str = $sformatf("%sio_writeback_16_bits_pdest = 0x%0h ",pkt_str,this.io_writeback_16_bits_pdest);
    pkt_str = $sformatf("%sio_writeback_16_bits_robIdx_flag = 0x%0h ",pkt_str,this.io_writeback_16_bits_robIdx_flag);
    pkt_str = $sformatf("%sio_writeback_16_bits_robIdx_value = 0x%0h ",pkt_str,this.io_writeback_16_bits_robIdx_value);
    pkt_str = $sformatf("%sio_writeback_16_bits_fpWen = 0x%0h ",pkt_str,this.io_writeback_16_bits_fpWen);
    pkt_str = $sformatf("%sio_writeback_16_bits_vecWen = 0x%0h ",pkt_str,this.io_writeback_16_bits_vecWen);
    pkt_str = $sformatf("%sio_writeback_16_bits_v0Wen = 0x%0h ",pkt_str,this.io_writeback_16_bits_v0Wen);
    pkt_str = $sformatf("%sio_writeback_16_bits_fflags = 0x%0h ",pkt_str,this.io_writeback_16_bits_fflags);
    pkt_str = $sformatf("%sio_writeback_16_bits_wflags = 0x%0h ",pkt_str,this.io_writeback_16_bits_wflags);
    pkt_str = $sformatf("%sio_writeback_16_bits_debugInfo_eliminatedMove = 0x%0h ",pkt_str,this.io_writeback_16_bits_debugInfo_eliminatedMove);
    pkt_str = $sformatf("%sio_writeback_16_bits_debugInfo_renameTime = 0x%0h ",pkt_str,this.io_writeback_16_bits_debugInfo_renameTime);
    pkt_str = $sformatf("%sio_writeback_16_bits_debugInfo_dispatchTime = 0x%0h ",pkt_str,this.io_writeback_16_bits_debugInfo_dispatchTime);
    pkt_str = $sformatf("%sio_writeback_16_bits_debugInfo_enqRsTime = 0x%0h ",pkt_str,this.io_writeback_16_bits_debugInfo_enqRsTime);
    pkt_str = $sformatf("%sio_writeback_16_bits_debugInfo_selectTime = 0x%0h ",pkt_str,this.io_writeback_16_bits_debugInfo_selectTime);
    pkt_str = $sformatf("%sio_writeback_16_bits_debugInfo_issueTime = 0x%0h ",pkt_str,this.io_writeback_16_bits_debugInfo_issueTime);
    pkt_str = $sformatf("%sio_writeback_16_bits_debugInfo_writebackTime = 0x%0h ",pkt_str,this.io_writeback_16_bits_debugInfo_writebackTime);
    pkt_str = $sformatf("%sio_writeback_16_bits_debugInfo_runahead_checkpoint_id = 0x%0h ",pkt_str,this.io_writeback_16_bits_debugInfo_runahead_checkpoint_id);
    pkt_str = $sformatf("%sio_writeback_16_bits_debugInfo_tlbFirstReqTime = 0x%0h ",pkt_str,this.io_writeback_16_bits_debugInfo_tlbFirstReqTime);
    pkt_str = $sformatf("%sio_writeback_16_bits_debugInfo_tlbRespTime = 0x%0h ",pkt_str,this.io_writeback_16_bits_debugInfo_tlbRespTime);
    pkt_str = $sformatf("%sio_writeback_16_bits_debug_seqNum = 0x%0h ",pkt_str,this.io_writeback_16_bits_debug_seqNum);
    pkt_str = $sformatf("%sio_writeback_15_valid = 0x%0h ",pkt_str,this.io_writeback_15_valid);
    pkt_str = $sformatf("%sio_writeback_15_bits_data_0 = 0x%0h ",pkt_str,this.io_writeback_15_bits_data_0);
    pkt_str = $sformatf("%sio_writeback_15_bits_data_1 = 0x%0h ",pkt_str,this.io_writeback_15_bits_data_1);
    pkt_str = $sformatf("%sio_writeback_15_bits_data_2 = 0x%0h ",pkt_str,this.io_writeback_15_bits_data_2);
    pkt_str = $sformatf("%sio_writeback_15_bits_pdest = 0x%0h ",pkt_str,this.io_writeback_15_bits_pdest);
    pkt_str = $sformatf("%sio_writeback_15_bits_robIdx_flag = 0x%0h ",pkt_str,this.io_writeback_15_bits_robIdx_flag);
    pkt_str = $sformatf("%sio_writeback_15_bits_robIdx_value = 0x%0h ",pkt_str,this.io_writeback_15_bits_robIdx_value);
    pkt_str = $sformatf("%sio_writeback_15_bits_vecWen = 0x%0h ",pkt_str,this.io_writeback_15_bits_vecWen);
    pkt_str = $sformatf("%sio_writeback_15_bits_v0Wen = 0x%0h ",pkt_str,this.io_writeback_15_bits_v0Wen);
    pkt_str = $sformatf("%sio_writeback_15_bits_fflags = 0x%0h ",pkt_str,this.io_writeback_15_bits_fflags);
    pkt_str = $sformatf("%sio_writeback_15_bits_wflags = 0x%0h ",pkt_str,this.io_writeback_15_bits_wflags);
    pkt_str = $sformatf("%sio_writeback_15_bits_vxsat = 0x%0h ",pkt_str,this.io_writeback_15_bits_vxsat);
    pkt_str = $sformatf("%sio_writeback_15_bits_debugInfo_eliminatedMove = 0x%0h ",pkt_str,this.io_writeback_15_bits_debugInfo_eliminatedMove);
    pkt_str = $sformatf("%sio_writeback_15_bits_debugInfo_renameTime = 0x%0h ",pkt_str,this.io_writeback_15_bits_debugInfo_renameTime);
    pkt_str = $sformatf("%sio_writeback_15_bits_debugInfo_dispatchTime = 0x%0h ",pkt_str,this.io_writeback_15_bits_debugInfo_dispatchTime);
    pkt_str = $sformatf("%sio_writeback_15_bits_debugInfo_enqRsTime = 0x%0h ",pkt_str,this.io_writeback_15_bits_debugInfo_enqRsTime);
    pkt_str = $sformatf("%sio_writeback_15_bits_debugInfo_selectTime = 0x%0h ",pkt_str,this.io_writeback_15_bits_debugInfo_selectTime);
    pkt_str = $sformatf("%sio_writeback_15_bits_debugInfo_issueTime = 0x%0h ",pkt_str,this.io_writeback_15_bits_debugInfo_issueTime);
    pkt_str = $sformatf("%sio_writeback_15_bits_debugInfo_writebackTime = 0x%0h ",pkt_str,this.io_writeback_15_bits_debugInfo_writebackTime);
    pkt_str = $sformatf("%sio_writeback_15_bits_debugInfo_runahead_checkpoint_id = 0x%0h ",pkt_str,this.io_writeback_15_bits_debugInfo_runahead_checkpoint_id);
    pkt_str = $sformatf("%sio_writeback_15_bits_debugInfo_tlbFirstReqTime = 0x%0h ",pkt_str,this.io_writeback_15_bits_debugInfo_tlbFirstReqTime);
    pkt_str = $sformatf("%sio_writeback_15_bits_debugInfo_tlbRespTime = 0x%0h ",pkt_str,this.io_writeback_15_bits_debugInfo_tlbRespTime);
    pkt_str = $sformatf("%sio_writeback_15_bits_debug_seqNum = 0x%0h ",pkt_str,this.io_writeback_15_bits_debug_seqNum);
    pkt_str = $sformatf("%sio_writeback_14_valid = 0x%0h ",pkt_str,this.io_writeback_14_valid);
    pkt_str = $sformatf("%sio_writeback_14_bits_data_0 = 0x%0h ",pkt_str,this.io_writeback_14_bits_data_0);
    pkt_str = $sformatf("%sio_writeback_14_bits_data_1 = 0x%0h ",pkt_str,this.io_writeback_14_bits_data_1);
    pkt_str = $sformatf("%sio_writeback_14_bits_data_2 = 0x%0h ",pkt_str,this.io_writeback_14_bits_data_2);
    pkt_str = $sformatf("%sio_writeback_14_bits_data_3 = 0x%0h ",pkt_str,this.io_writeback_14_bits_data_3);
    pkt_str = $sformatf("%sio_writeback_14_bits_data_4 = 0x%0h ",pkt_str,this.io_writeback_14_bits_data_4);
    pkt_str = $sformatf("%sio_writeback_14_bits_data_5 = 0x%0h ",pkt_str,this.io_writeback_14_bits_data_5);
    pkt_str = $sformatf("%sio_writeback_14_bits_pdest = 0x%0h ",pkt_str,this.io_writeback_14_bits_pdest);
    pkt_str = $sformatf("%sio_writeback_14_bits_robIdx_flag = 0x%0h ",pkt_str,this.io_writeback_14_bits_robIdx_flag);
    pkt_str = $sformatf("%sio_writeback_14_bits_robIdx_value = 0x%0h ",pkt_str,this.io_writeback_14_bits_robIdx_value);
    pkt_str = $sformatf("%sio_writeback_14_bits_intWen = 0x%0h ",pkt_str,this.io_writeback_14_bits_intWen);
    pkt_str = $sformatf("%sio_writeback_14_bits_fpWen = 0x%0h ",pkt_str,this.io_writeback_14_bits_fpWen);
    pkt_str = $sformatf("%sio_writeback_14_bits_vecWen = 0x%0h ",pkt_str,this.io_writeback_14_bits_vecWen);
    pkt_str = $sformatf("%sio_writeback_14_bits_v0Wen = 0x%0h ",pkt_str,this.io_writeback_14_bits_v0Wen);
    pkt_str = $sformatf("%sio_writeback_14_bits_vlWen = 0x%0h ",pkt_str,this.io_writeback_14_bits_vlWen);
    pkt_str = $sformatf("%sio_writeback_14_bits_fflags = 0x%0h ",pkt_str,this.io_writeback_14_bits_fflags);
    pkt_str = $sformatf("%sio_writeback_14_bits_wflags = 0x%0h ",pkt_str,this.io_writeback_14_bits_wflags);
    pkt_str = $sformatf("%sio_writeback_14_bits_exceptionVec_2 = 0x%0h ",pkt_str,this.io_writeback_14_bits_exceptionVec_2);
    pkt_str = $sformatf("%sio_writeback_14_bits_debugInfo_eliminatedMove = 0x%0h ",pkt_str,this.io_writeback_14_bits_debugInfo_eliminatedMove);
    pkt_str = $sformatf("%sio_writeback_14_bits_debugInfo_renameTime = 0x%0h ",pkt_str,this.io_writeback_14_bits_debugInfo_renameTime);
    pkt_str = $sformatf("%sio_writeback_14_bits_debugInfo_dispatchTime = 0x%0h ",pkt_str,this.io_writeback_14_bits_debugInfo_dispatchTime);
    pkt_str = $sformatf("%sio_writeback_14_bits_debugInfo_enqRsTime = 0x%0h ",pkt_str,this.io_writeback_14_bits_debugInfo_enqRsTime);
    pkt_str = $sformatf("%sio_writeback_14_bits_debugInfo_selectTime = 0x%0h ",pkt_str,this.io_writeback_14_bits_debugInfo_selectTime);
    pkt_str = $sformatf("%sio_writeback_14_bits_debugInfo_issueTime = 0x%0h ",pkt_str,this.io_writeback_14_bits_debugInfo_issueTime);
    pkt_str = $sformatf("%sio_writeback_14_bits_debugInfo_writebackTime = 0x%0h ",pkt_str,this.io_writeback_14_bits_debugInfo_writebackTime);
    pkt_str = $sformatf("%sio_writeback_14_bits_debugInfo_runahead_checkpoint_id = 0x%0h ",pkt_str,this.io_writeback_14_bits_debugInfo_runahead_checkpoint_id);
    pkt_str = $sformatf("%sio_writeback_14_bits_debugInfo_tlbFirstReqTime = 0x%0h ",pkt_str,this.io_writeback_14_bits_debugInfo_tlbFirstReqTime);
    pkt_str = $sformatf("%sio_writeback_14_bits_debugInfo_tlbRespTime = 0x%0h ",pkt_str,this.io_writeback_14_bits_debugInfo_tlbRespTime);
    pkt_str = $sformatf("%sio_writeback_14_bits_debug_seqNum = 0x%0h ",pkt_str,this.io_writeback_14_bits_debug_seqNum);
    pkt_str = $sformatf("%sio_writeback_13_valid = 0x%0h ",pkt_str,this.io_writeback_13_valid);
    pkt_str = $sformatf("%sio_writeback_13_bits_data_0 = 0x%0h ",pkt_str,this.io_writeback_13_bits_data_0);
    pkt_str = $sformatf("%sio_writeback_13_bits_data_1 = 0x%0h ",pkt_str,this.io_writeback_13_bits_data_1);
    pkt_str = $sformatf("%sio_writeback_13_bits_data_2 = 0x%0h ",pkt_str,this.io_writeback_13_bits_data_2);
    pkt_str = $sformatf("%sio_writeback_13_bits_pdest = 0x%0h ",pkt_str,this.io_writeback_13_bits_pdest);
    pkt_str = $sformatf("%sio_writeback_13_bits_robIdx_flag = 0x%0h ",pkt_str,this.io_writeback_13_bits_robIdx_flag);
    pkt_str = $sformatf("%sio_writeback_13_bits_robIdx_value = 0x%0h ",pkt_str,this.io_writeback_13_bits_robIdx_value);
    pkt_str = $sformatf("%sio_writeback_13_bits_vecWen = 0x%0h ",pkt_str,this.io_writeback_13_bits_vecWen);
    pkt_str = $sformatf("%sio_writeback_13_bits_v0Wen = 0x%0h ",pkt_str,this.io_writeback_13_bits_v0Wen);
    pkt_str = $sformatf("%sio_writeback_13_bits_fflags = 0x%0h ",pkt_str,this.io_writeback_13_bits_fflags);
    pkt_str = $sformatf("%sio_writeback_13_bits_wflags = 0x%0h ",pkt_str,this.io_writeback_13_bits_wflags);
    pkt_str = $sformatf("%sio_writeback_13_bits_vxsat = 0x%0h ",pkt_str,this.io_writeback_13_bits_vxsat);
    pkt_str = $sformatf("%sio_writeback_13_bits_exceptionVec_2 = 0x%0h ",pkt_str,this.io_writeback_13_bits_exceptionVec_2);
    pkt_str = $sformatf("%sio_writeback_13_bits_debugInfo_eliminatedMove = 0x%0h ",pkt_str,this.io_writeback_13_bits_debugInfo_eliminatedMove);
    pkt_str = $sformatf("%sio_writeback_13_bits_debugInfo_renameTime = 0x%0h ",pkt_str,this.io_writeback_13_bits_debugInfo_renameTime);
    pkt_str = $sformatf("%sio_writeback_13_bits_debugInfo_dispatchTime = 0x%0h ",pkt_str,this.io_writeback_13_bits_debugInfo_dispatchTime);
    pkt_str = $sformatf("%sio_writeback_13_bits_debugInfo_enqRsTime = 0x%0h ",pkt_str,this.io_writeback_13_bits_debugInfo_enqRsTime);
    pkt_str = $sformatf("%sio_writeback_13_bits_debugInfo_selectTime = 0x%0h ",pkt_str,this.io_writeback_13_bits_debugInfo_selectTime);
    pkt_str = $sformatf("%sio_writeback_13_bits_debugInfo_issueTime = 0x%0h ",pkt_str,this.io_writeback_13_bits_debugInfo_issueTime);
    pkt_str = $sformatf("%sio_writeback_13_bits_debugInfo_writebackTime = 0x%0h ",pkt_str,this.io_writeback_13_bits_debugInfo_writebackTime);
    pkt_str = $sformatf("%sio_writeback_13_bits_debugInfo_runahead_checkpoint_id = 0x%0h ",pkt_str,this.io_writeback_13_bits_debugInfo_runahead_checkpoint_id);
    pkt_str = $sformatf("%sio_writeback_13_bits_debugInfo_tlbFirstReqTime = 0x%0h ",pkt_str,this.io_writeback_13_bits_debugInfo_tlbFirstReqTime);
    pkt_str = $sformatf("%sio_writeback_13_bits_debugInfo_tlbRespTime = 0x%0h ",pkt_str,this.io_writeback_13_bits_debugInfo_tlbRespTime);
    pkt_str = $sformatf("%sio_writeback_13_bits_debug_seqNum = 0x%0h ",pkt_str,this.io_writeback_13_bits_debug_seqNum);
    pkt_str = $sformatf("%sio_writeback_7_valid = 0x%0h ",pkt_str,this.io_writeback_7_valid);
    pkt_str = $sformatf("%sio_writeback_7_bits_data_0 = 0x%0h ",pkt_str,this.io_writeback_7_bits_data_0);
    pkt_str = $sformatf("%sio_writeback_7_bits_data_1 = 0x%0h ",pkt_str,this.io_writeback_7_bits_data_1);
    pkt_str = $sformatf("%sio_writeback_7_bits_pdest = 0x%0h ",pkt_str,this.io_writeback_7_bits_pdest);
    pkt_str = $sformatf("%sio_writeback_7_bits_robIdx_flag = 0x%0h ",pkt_str,this.io_writeback_7_bits_robIdx_flag);
    pkt_str = $sformatf("%sio_writeback_7_bits_robIdx_value = 0x%0h ",pkt_str,this.io_writeback_7_bits_robIdx_value);
    pkt_str = $sformatf("%sio_writeback_7_bits_intWen = 0x%0h ",pkt_str,this.io_writeback_7_bits_intWen);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_valid = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_valid);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_isRVC = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_isRVC);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_robIdx_flag = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_robIdx_flag);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_robIdx_value = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_robIdx_value);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_ftqIdx_flag = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_ftqIdx_flag);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_ftqIdx_value = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_ftqIdx_value);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_ftqOffset = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_ftqOffset);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_level = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_level);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_interrupt = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_interrupt);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_pc = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_pc);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_ssp = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_ssp);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_sctr = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_sctr);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_topAddr = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0 = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1 = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2 = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3 = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0 = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1 = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2 = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3 = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0 = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1 = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2 = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3 = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0 = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1 = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2 = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3 = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0 = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1 = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2 = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3 = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0 = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1 = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2 = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3 = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_ghr = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_ghr);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0 = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1 = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_br_hit = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_predTaken = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_target = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_target);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_taken = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_taken);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_shift = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_shift);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_fullTarget = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_fullTarget);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_stFtqIdx_flag = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_stFtqIdx_flag);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_stFtqIdx_value = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_stFtqIdx_value);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_stFtqOffset = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_stFtqOffset);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_debugIsCtrl = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_debugIsCtrl);
    pkt_str = $sformatf("%sio_writeback_7_bits_redirect_bits_debugIsMemVio = 0x%0h ",pkt_str,this.io_writeback_7_bits_redirect_bits_debugIsMemVio);
    pkt_str = $sformatf("%sio_writeback_7_bits_exceptionVec_2 = 0x%0h ",pkt_str,this.io_writeback_7_bits_exceptionVec_2);
    pkt_str = $sformatf("%sio_writeback_7_bits_exceptionVec_3 = 0x%0h ",pkt_str,this.io_writeback_7_bits_exceptionVec_3);
    pkt_str = $sformatf("%sio_writeback_7_bits_exceptionVec_8 = 0x%0h ",pkt_str,this.io_writeback_7_bits_exceptionVec_8);
    pkt_str = $sformatf("%sio_writeback_7_bits_exceptionVec_9 = 0x%0h ",pkt_str,this.io_writeback_7_bits_exceptionVec_9);
    pkt_str = $sformatf("%sio_writeback_7_bits_exceptionVec_10 = 0x%0h ",pkt_str,this.io_writeback_7_bits_exceptionVec_10);
    pkt_str = $sformatf("%sio_writeback_7_bits_exceptionVec_11 = 0x%0h ",pkt_str,this.io_writeback_7_bits_exceptionVec_11);
    pkt_str = $sformatf("%sio_writeback_7_bits_exceptionVec_22 = 0x%0h ",pkt_str,this.io_writeback_7_bits_exceptionVec_22);
    pkt_str = $sformatf("%sio_writeback_7_bits_flushPipe = 0x%0h ",pkt_str,this.io_writeback_7_bits_flushPipe);
    pkt_str = $sformatf("%sio_writeback_7_bits_predecodeInfo_valid = 0x%0h ",pkt_str,this.io_writeback_7_bits_predecodeInfo_valid);
    pkt_str = $sformatf("%sio_writeback_7_bits_predecodeInfo_isRVC = 0x%0h ",pkt_str,this.io_writeback_7_bits_predecodeInfo_isRVC);
    pkt_str = $sformatf("%sio_writeback_7_bits_predecodeInfo_brType = 0x%0h ",pkt_str,this.io_writeback_7_bits_predecodeInfo_brType);
    pkt_str = $sformatf("%sio_writeback_7_bits_predecodeInfo_isCall = 0x%0h ",pkt_str,this.io_writeback_7_bits_predecodeInfo_isCall);
    pkt_str = $sformatf("%sio_writeback_7_bits_predecodeInfo_isRet = 0x%0h ",pkt_str,this.io_writeback_7_bits_predecodeInfo_isRet);
    pkt_str = $sformatf("%sio_writeback_7_bits_debug_isPerfCnt = 0x%0h ",pkt_str,this.io_writeback_7_bits_debug_isPerfCnt);
    pkt_str = $sformatf("%sio_writeback_7_bits_debugInfo_eliminatedMove = 0x%0h ",pkt_str,this.io_writeback_7_bits_debugInfo_eliminatedMove);
    pkt_str = $sformatf("%sio_writeback_7_bits_debugInfo_renameTime = 0x%0h ",pkt_str,this.io_writeback_7_bits_debugInfo_renameTime);
    pkt_str = $sformatf("%sio_writeback_7_bits_debugInfo_dispatchTime = 0x%0h ",pkt_str,this.io_writeback_7_bits_debugInfo_dispatchTime);
    pkt_str = $sformatf("%sio_writeback_7_bits_debugInfo_enqRsTime = 0x%0h ",pkt_str,this.io_writeback_7_bits_debugInfo_enqRsTime);
    pkt_str = $sformatf("%sio_writeback_7_bits_debugInfo_selectTime = 0x%0h ",pkt_str,this.io_writeback_7_bits_debugInfo_selectTime);
    pkt_str = $sformatf("%sio_writeback_7_bits_debugInfo_issueTime = 0x%0h ",pkt_str,this.io_writeback_7_bits_debugInfo_issueTime);
    pkt_str = $sformatf("%sio_writeback_7_bits_debugInfo_writebackTime = 0x%0h ",pkt_str,this.io_writeback_7_bits_debugInfo_writebackTime);
    pkt_str = $sformatf("%sio_writeback_7_bits_debugInfo_runahead_checkpoint_id = 0x%0h ",pkt_str,this.io_writeback_7_bits_debugInfo_runahead_checkpoint_id);
    pkt_str = $sformatf("%sio_writeback_7_bits_debugInfo_tlbFirstReqTime = 0x%0h ",pkt_str,this.io_writeback_7_bits_debugInfo_tlbFirstReqTime);
    pkt_str = $sformatf("%sio_writeback_7_bits_debugInfo_tlbRespTime = 0x%0h ",pkt_str,this.io_writeback_7_bits_debugInfo_tlbRespTime);
    pkt_str = $sformatf("%sio_writeback_7_bits_debug_seqNum = 0x%0h ",pkt_str,this.io_writeback_7_bits_debug_seqNum);
    pkt_str = $sformatf("%sio_writeback_5_valid = 0x%0h ",pkt_str,this.io_writeback_5_valid);
    pkt_str = $sformatf("%sio_writeback_5_bits_redirect_valid = 0x%0h ",pkt_str,this.io_writeback_5_bits_redirect_valid);
    pkt_str = $sformatf("%sio_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred = 0x%0h ",pkt_str,this.io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred);
    pkt_str = $sformatf("%sio_writeback_3_valid = 0x%0h ",pkt_str,this.io_writeback_3_valid);
    pkt_str = $sformatf("%sio_writeback_3_bits_redirect_valid = 0x%0h ",pkt_str,this.io_writeback_3_bits_redirect_valid);
    pkt_str = $sformatf("%sio_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred = 0x%0h ",pkt_str,this.io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred);
    pkt_str = $sformatf("%sio_writeback_1_valid = 0x%0h ",pkt_str,this.io_writeback_1_valid);
    pkt_str = $sformatf("%sio_writeback_1_bits_redirect_valid = 0x%0h ",pkt_str,this.io_writeback_1_bits_redirect_valid);
    pkt_str = $sformatf("%sio_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred = 0x%0h ",pkt_str,this.io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred);
    pkt_str = $sformatf("%sio_exuWriteback_26_valid = 0x%0h ",pkt_str,this.io_exuWriteback_26_valid);
    pkt_str = $sformatf("%sio_exuWriteback_26_bits_robIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_26_bits_robIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_25_valid = 0x%0h ",pkt_str,this.io_exuWriteback_25_valid);
    pkt_str = $sformatf("%sio_exuWriteback_25_bits_robIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_25_bits_robIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_24_valid = 0x%0h ",pkt_str,this.io_exuWriteback_24_valid);
    pkt_str = $sformatf("%sio_exuWriteback_24_bits_data_0 = 0x%0h ",pkt_str,this.io_exuWriteback_24_bits_data_0);
    pkt_str = $sformatf("%sio_exuWriteback_24_bits_pdest = 0x%0h ",pkt_str,this.io_exuWriteback_24_bits_pdest);
    pkt_str = $sformatf("%sio_exuWriteback_24_bits_robIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_24_bits_robIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_24_bits_vecWen = 0x%0h ",pkt_str,this.io_exuWriteback_24_bits_vecWen);
    pkt_str = $sformatf("%sio_exuWriteback_24_bits_v0Wen = 0x%0h ",pkt_str,this.io_exuWriteback_24_bits_v0Wen);
    pkt_str = $sformatf("%sio_exuWriteback_24_bits_vls_vdIdx = 0x%0h ",pkt_str,this.io_exuWriteback_24_bits_vls_vdIdx);
    pkt_str = $sformatf("%sio_exuWriteback_24_bits_debug_isMMIO = 0x%0h ",pkt_str,this.io_exuWriteback_24_bits_debug_isMMIO);
    pkt_str = $sformatf("%sio_exuWriteback_24_bits_debug_isNCIO = 0x%0h ",pkt_str,this.io_exuWriteback_24_bits_debug_isNCIO);
    pkt_str = $sformatf("%sio_exuWriteback_24_bits_debug_isPerfCnt = 0x%0h ",pkt_str,this.io_exuWriteback_24_bits_debug_isPerfCnt);
    pkt_str = $sformatf("%sio_exuWriteback_24_bits_debug_paddr = 0x%0h ",pkt_str,this.io_exuWriteback_24_bits_debug_paddr);
    pkt_str = $sformatf("%sio_exuWriteback_23_valid = 0x%0h ",pkt_str,this.io_exuWriteback_23_valid);
    pkt_str = $sformatf("%sio_exuWriteback_23_bits_data_0 = 0x%0h ",pkt_str,this.io_exuWriteback_23_bits_data_0);
    pkt_str = $sformatf("%sio_exuWriteback_23_bits_pdest = 0x%0h ",pkt_str,this.io_exuWriteback_23_bits_pdest);
    pkt_str = $sformatf("%sio_exuWriteback_23_bits_robIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_23_bits_robIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_23_bits_vecWen = 0x%0h ",pkt_str,this.io_exuWriteback_23_bits_vecWen);
    pkt_str = $sformatf("%sio_exuWriteback_23_bits_v0Wen = 0x%0h ",pkt_str,this.io_exuWriteback_23_bits_v0Wen);
    pkt_str = $sformatf("%sio_exuWriteback_23_bits_vls_vdIdx = 0x%0h ",pkt_str,this.io_exuWriteback_23_bits_vls_vdIdx);
    pkt_str = $sformatf("%sio_exuWriteback_23_bits_debug_isMMIO = 0x%0h ",pkt_str,this.io_exuWriteback_23_bits_debug_isMMIO);
    pkt_str = $sformatf("%sio_exuWriteback_23_bits_debug_isNCIO = 0x%0h ",pkt_str,this.io_exuWriteback_23_bits_debug_isNCIO);
    pkt_str = $sformatf("%sio_exuWriteback_23_bits_debug_isPerfCnt = 0x%0h ",pkt_str,this.io_exuWriteback_23_bits_debug_isPerfCnt);
    pkt_str = $sformatf("%sio_exuWriteback_23_bits_debug_paddr = 0x%0h ",pkt_str,this.io_exuWriteback_23_bits_debug_paddr);
    pkt_str = $sformatf("%sio_exuWriteback_22_valid = 0x%0h ",pkt_str,this.io_exuWriteback_22_valid);
    pkt_str = $sformatf("%sio_exuWriteback_22_bits_data_0 = 0x%0h ",pkt_str,this.io_exuWriteback_22_bits_data_0);
    pkt_str = $sformatf("%sio_exuWriteback_22_bits_robIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_22_bits_robIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_22_bits_lqIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_22_bits_lqIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_22_bits_debug_isMMIO = 0x%0h ",pkt_str,this.io_exuWriteback_22_bits_debug_isMMIO);
    pkt_str = $sformatf("%sio_exuWriteback_22_bits_debug_isNCIO = 0x%0h ",pkt_str,this.io_exuWriteback_22_bits_debug_isNCIO);
    pkt_str = $sformatf("%sio_exuWriteback_22_bits_debug_isPerfCnt = 0x%0h ",pkt_str,this.io_exuWriteback_22_bits_debug_isPerfCnt);
    pkt_str = $sformatf("%sio_exuWriteback_22_bits_debug_paddr = 0x%0h ",pkt_str,this.io_exuWriteback_22_bits_debug_paddr);
    pkt_str = $sformatf("%sio_exuWriteback_21_valid = 0x%0h ",pkt_str,this.io_exuWriteback_21_valid);
    pkt_str = $sformatf("%sio_exuWriteback_21_bits_data_0 = 0x%0h ",pkt_str,this.io_exuWriteback_21_bits_data_0);
    pkt_str = $sformatf("%sio_exuWriteback_21_bits_robIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_21_bits_robIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_21_bits_lqIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_21_bits_lqIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_21_bits_debug_isMMIO = 0x%0h ",pkt_str,this.io_exuWriteback_21_bits_debug_isMMIO);
    pkt_str = $sformatf("%sio_exuWriteback_21_bits_debug_isNCIO = 0x%0h ",pkt_str,this.io_exuWriteback_21_bits_debug_isNCIO);
    pkt_str = $sformatf("%sio_exuWriteback_21_bits_debug_isPerfCnt = 0x%0h ",pkt_str,this.io_exuWriteback_21_bits_debug_isPerfCnt);
    pkt_str = $sformatf("%sio_exuWriteback_21_bits_debug_paddr = 0x%0h ",pkt_str,this.io_exuWriteback_21_bits_debug_paddr);
    pkt_str = $sformatf("%sio_exuWriteback_20_valid = 0x%0h ",pkt_str,this.io_exuWriteback_20_valid);
    pkt_str = $sformatf("%sio_exuWriteback_20_bits_data_0 = 0x%0h ",pkt_str,this.io_exuWriteback_20_bits_data_0);
    pkt_str = $sformatf("%sio_exuWriteback_20_bits_robIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_20_bits_robIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_20_bits_lqIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_20_bits_lqIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_20_bits_debug_isMMIO = 0x%0h ",pkt_str,this.io_exuWriteback_20_bits_debug_isMMIO);
    pkt_str = $sformatf("%sio_exuWriteback_20_bits_debug_isNCIO = 0x%0h ",pkt_str,this.io_exuWriteback_20_bits_debug_isNCIO);
    pkt_str = $sformatf("%sio_exuWriteback_20_bits_debug_isPerfCnt = 0x%0h ",pkt_str,this.io_exuWriteback_20_bits_debug_isPerfCnt);
    pkt_str = $sformatf("%sio_exuWriteback_20_bits_debug_paddr = 0x%0h ",pkt_str,this.io_exuWriteback_20_bits_debug_paddr);
    pkt_str = $sformatf("%sio_exuWriteback_19_valid = 0x%0h ",pkt_str,this.io_exuWriteback_19_valid);
    pkt_str = $sformatf("%sio_exuWriteback_19_bits_data_0 = 0x%0h ",pkt_str,this.io_exuWriteback_19_bits_data_0);
    pkt_str = $sformatf("%sio_exuWriteback_19_bits_robIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_19_bits_robIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_19_bits_sqIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_19_bits_sqIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_19_bits_debug_isMMIO = 0x%0h ",pkt_str,this.io_exuWriteback_19_bits_debug_isMMIO);
    pkt_str = $sformatf("%sio_exuWriteback_19_bits_debug_isNCIO = 0x%0h ",pkt_str,this.io_exuWriteback_19_bits_debug_isNCIO);
    pkt_str = $sformatf("%sio_exuWriteback_19_bits_debug_isPerfCnt = 0x%0h ",pkt_str,this.io_exuWriteback_19_bits_debug_isPerfCnt);
    pkt_str = $sformatf("%sio_exuWriteback_19_bits_debug_paddr = 0x%0h ",pkt_str,this.io_exuWriteback_19_bits_debug_paddr);
    pkt_str = $sformatf("%sio_exuWriteback_18_valid = 0x%0h ",pkt_str,this.io_exuWriteback_18_valid);
    pkt_str = $sformatf("%sio_exuWriteback_18_bits_data_0 = 0x%0h ",pkt_str,this.io_exuWriteback_18_bits_data_0);
    pkt_str = $sformatf("%sio_exuWriteback_18_bits_robIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_18_bits_robIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_18_bits_sqIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_18_bits_sqIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_18_bits_debug_isMMIO = 0x%0h ",pkt_str,this.io_exuWriteback_18_bits_debug_isMMIO);
    pkt_str = $sformatf("%sio_exuWriteback_18_bits_debug_isNCIO = 0x%0h ",pkt_str,this.io_exuWriteback_18_bits_debug_isNCIO);
    pkt_str = $sformatf("%sio_exuWriteback_18_bits_debug_isPerfCnt = 0x%0h ",pkt_str,this.io_exuWriteback_18_bits_debug_isPerfCnt);
    pkt_str = $sformatf("%sio_exuWriteback_18_bits_debug_paddr = 0x%0h ",pkt_str,this.io_exuWriteback_18_bits_debug_paddr);
    pkt_str = $sformatf("%sio_exuWriteback_17_valid = 0x%0h ",pkt_str,this.io_exuWriteback_17_valid);
    pkt_str = $sformatf("%sio_exuWriteback_17_bits_data_0 = 0x%0h ",pkt_str,this.io_exuWriteback_17_bits_data_0);
    pkt_str = $sformatf("%sio_exuWriteback_17_bits_robIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_17_bits_robIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_17_bits_fflags = 0x%0h ",pkt_str,this.io_exuWriteback_17_bits_fflags);
    pkt_str = $sformatf("%sio_exuWriteback_17_bits_wflags = 0x%0h ",pkt_str,this.io_exuWriteback_17_bits_wflags);
    pkt_str = $sformatf("%sio_exuWriteback_16_valid = 0x%0h ",pkt_str,this.io_exuWriteback_16_valid);
    pkt_str = $sformatf("%sio_exuWriteback_16_bits_data_0 = 0x%0h ",pkt_str,this.io_exuWriteback_16_bits_data_0);
    pkt_str = $sformatf("%sio_exuWriteback_16_bits_robIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_16_bits_robIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_16_bits_fflags = 0x%0h ",pkt_str,this.io_exuWriteback_16_bits_fflags);
    pkt_str = $sformatf("%sio_exuWriteback_16_bits_wflags = 0x%0h ",pkt_str,this.io_exuWriteback_16_bits_wflags);
    pkt_str = $sformatf("%sio_exuWriteback_15_valid = 0x%0h ",pkt_str,this.io_exuWriteback_15_valid);
    pkt_str = $sformatf("%sio_exuWriteback_15_bits_data_0 = 0x%0h ",pkt_str,this.io_exuWriteback_15_bits_data_0);
    pkt_str = $sformatf("%sio_exuWriteback_15_bits_robIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_15_bits_robIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_15_bits_fflags = 0x%0h ",pkt_str,this.io_exuWriteback_15_bits_fflags);
    pkt_str = $sformatf("%sio_exuWriteback_15_bits_wflags = 0x%0h ",pkt_str,this.io_exuWriteback_15_bits_wflags);
    pkt_str = $sformatf("%sio_exuWriteback_15_bits_vxsat = 0x%0h ",pkt_str,this.io_exuWriteback_15_bits_vxsat);
    pkt_str = $sformatf("%sio_exuWriteback_14_valid = 0x%0h ",pkt_str,this.io_exuWriteback_14_valid);
    pkt_str = $sformatf("%sio_exuWriteback_14_bits_data_0 = 0x%0h ",pkt_str,this.io_exuWriteback_14_bits_data_0);
    pkt_str = $sformatf("%sio_exuWriteback_14_bits_robIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_14_bits_robIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_14_bits_fflags = 0x%0h ",pkt_str,this.io_exuWriteback_14_bits_fflags);
    pkt_str = $sformatf("%sio_exuWriteback_14_bits_wflags = 0x%0h ",pkt_str,this.io_exuWriteback_14_bits_wflags);
    pkt_str = $sformatf("%sio_exuWriteback_13_valid = 0x%0h ",pkt_str,this.io_exuWriteback_13_valid);
    pkt_str = $sformatf("%sio_exuWriteback_13_bits_data_0 = 0x%0h ",pkt_str,this.io_exuWriteback_13_bits_data_0);
    pkt_str = $sformatf("%sio_exuWriteback_13_bits_robIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_13_bits_robIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_13_bits_fflags = 0x%0h ",pkt_str,this.io_exuWriteback_13_bits_fflags);
    pkt_str = $sformatf("%sio_exuWriteback_13_bits_wflags = 0x%0h ",pkt_str,this.io_exuWriteback_13_bits_wflags);
    pkt_str = $sformatf("%sio_exuWriteback_13_bits_vxsat = 0x%0h ",pkt_str,this.io_exuWriteback_13_bits_vxsat);
    pkt_str = $sformatf("%sio_exuWriteback_12_valid = 0x%0h ",pkt_str,this.io_exuWriteback_12_valid);
    pkt_str = $sformatf("%sio_exuWriteback_12_bits_data_0 = 0x%0h ",pkt_str,this.io_exuWriteback_12_bits_data_0);
    pkt_str = $sformatf("%sio_exuWriteback_12_bits_robIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_12_bits_robIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_12_bits_fflags = 0x%0h ",pkt_str,this.io_exuWriteback_12_bits_fflags);
    pkt_str = $sformatf("%sio_exuWriteback_12_bits_wflags = 0x%0h ",pkt_str,this.io_exuWriteback_12_bits_wflags);
    pkt_str = $sformatf("%sio_exuWriteback_11_valid = 0x%0h ",pkt_str,this.io_exuWriteback_11_valid);
    pkt_str = $sformatf("%sio_exuWriteback_11_bits_data_0 = 0x%0h ",pkt_str,this.io_exuWriteback_11_bits_data_0);
    pkt_str = $sformatf("%sio_exuWriteback_11_bits_robIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_11_bits_robIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_11_bits_fflags = 0x%0h ",pkt_str,this.io_exuWriteback_11_bits_fflags);
    pkt_str = $sformatf("%sio_exuWriteback_11_bits_wflags = 0x%0h ",pkt_str,this.io_exuWriteback_11_bits_wflags);
    pkt_str = $sformatf("%sio_exuWriteback_10_valid = 0x%0h ",pkt_str,this.io_exuWriteback_10_valid);
    pkt_str = $sformatf("%sio_exuWriteback_10_bits_data_0 = 0x%0h ",pkt_str,this.io_exuWriteback_10_bits_data_0);
    pkt_str = $sformatf("%sio_exuWriteback_10_bits_robIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_10_bits_robIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_10_bits_fflags = 0x%0h ",pkt_str,this.io_exuWriteback_10_bits_fflags);
    pkt_str = $sformatf("%sio_exuWriteback_10_bits_wflags = 0x%0h ",pkt_str,this.io_exuWriteback_10_bits_wflags);
    pkt_str = $sformatf("%sio_exuWriteback_9_valid = 0x%0h ",pkt_str,this.io_exuWriteback_9_valid);
    pkt_str = $sformatf("%sio_exuWriteback_9_bits_data_0 = 0x%0h ",pkt_str,this.io_exuWriteback_9_bits_data_0);
    pkt_str = $sformatf("%sio_exuWriteback_9_bits_robIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_9_bits_robIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_9_bits_fflags = 0x%0h ",pkt_str,this.io_exuWriteback_9_bits_fflags);
    pkt_str = $sformatf("%sio_exuWriteback_9_bits_wflags = 0x%0h ",pkt_str,this.io_exuWriteback_9_bits_wflags);
    pkt_str = $sformatf("%sio_exuWriteback_8_valid = 0x%0h ",pkt_str,this.io_exuWriteback_8_valid);
    pkt_str = $sformatf("%sio_exuWriteback_8_bits_data_0 = 0x%0h ",pkt_str,this.io_exuWriteback_8_bits_data_0);
    pkt_str = $sformatf("%sio_exuWriteback_8_bits_robIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_8_bits_robIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_8_bits_fflags = 0x%0h ",pkt_str,this.io_exuWriteback_8_bits_fflags);
    pkt_str = $sformatf("%sio_exuWriteback_8_bits_wflags = 0x%0h ",pkt_str,this.io_exuWriteback_8_bits_wflags);
    pkt_str = $sformatf("%sio_exuWriteback_7_valid = 0x%0h ",pkt_str,this.io_exuWriteback_7_valid);
    pkt_str = $sformatf("%sio_exuWriteback_7_bits_data_0 = 0x%0h ",pkt_str,this.io_exuWriteback_7_bits_data_0);
    pkt_str = $sformatf("%sio_exuWriteback_7_bits_robIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_7_bits_robIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_7_bits_debug_isPerfCnt = 0x%0h ",pkt_str,this.io_exuWriteback_7_bits_debug_isPerfCnt);
    pkt_str = $sformatf("%sio_exuWriteback_6_valid = 0x%0h ",pkt_str,this.io_exuWriteback_6_valid);
    pkt_str = $sformatf("%sio_exuWriteback_6_bits_data_0 = 0x%0h ",pkt_str,this.io_exuWriteback_6_bits_data_0);
    pkt_str = $sformatf("%sio_exuWriteback_6_bits_robIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_6_bits_robIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_5_valid = 0x%0h ",pkt_str,this.io_exuWriteback_5_valid);
    pkt_str = $sformatf("%sio_exuWriteback_5_bits_data_0 = 0x%0h ",pkt_str,this.io_exuWriteback_5_bits_data_0);
    pkt_str = $sformatf("%sio_exuWriteback_5_bits_robIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_5_bits_robIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_5_bits_redirect_valid = 0x%0h ",pkt_str,this.io_exuWriteback_5_bits_redirect_valid);
    pkt_str = $sformatf("%sio_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken = 0x%0h ",pkt_str,this.io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken);
    pkt_str = $sformatf("%sio_exuWriteback_5_bits_fflags = 0x%0h ",pkt_str,this.io_exuWriteback_5_bits_fflags);
    pkt_str = $sformatf("%sio_exuWriteback_5_bits_wflags = 0x%0h ",pkt_str,this.io_exuWriteback_5_bits_wflags);
    pkt_str = $sformatf("%sio_exuWriteback_4_valid = 0x%0h ",pkt_str,this.io_exuWriteback_4_valid);
    pkt_str = $sformatf("%sio_exuWriteback_4_bits_data_0 = 0x%0h ",pkt_str,this.io_exuWriteback_4_bits_data_0);
    pkt_str = $sformatf("%sio_exuWriteback_4_bits_robIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_4_bits_robIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_3_valid = 0x%0h ",pkt_str,this.io_exuWriteback_3_valid);
    pkt_str = $sformatf("%sio_exuWriteback_3_bits_data_0 = 0x%0h ",pkt_str,this.io_exuWriteback_3_bits_data_0);
    pkt_str = $sformatf("%sio_exuWriteback_3_bits_robIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_3_bits_robIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_3_bits_redirect_valid = 0x%0h ",pkt_str,this.io_exuWriteback_3_bits_redirect_valid);
    pkt_str = $sformatf("%sio_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken = 0x%0h ",pkt_str,this.io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken);
    pkt_str = $sformatf("%sio_exuWriteback_2_valid = 0x%0h ",pkt_str,this.io_exuWriteback_2_valid);
    pkt_str = $sformatf("%sio_exuWriteback_2_bits_data_0 = 0x%0h ",pkt_str,this.io_exuWriteback_2_bits_data_0);
    pkt_str = $sformatf("%sio_exuWriteback_2_bits_robIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_2_bits_robIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_1_valid = 0x%0h ",pkt_str,this.io_exuWriteback_1_valid);
    pkt_str = $sformatf("%sio_exuWriteback_1_bits_data_0 = 0x%0h ",pkt_str,this.io_exuWriteback_1_bits_data_0);
    pkt_str = $sformatf("%sio_exuWriteback_1_bits_robIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_1_bits_robIdx_value);
    pkt_str = $sformatf("%sio_exuWriteback_1_bits_redirect_valid = 0x%0h ",pkt_str,this.io_exuWriteback_1_bits_redirect_valid);
    pkt_str = $sformatf("%sio_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken = 0x%0h ",pkt_str,this.io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken);
    pkt_str = $sformatf("%sio_exuWriteback_0_valid = 0x%0h ",pkt_str,this.io_exuWriteback_0_valid);
    pkt_str = $sformatf("%sio_exuWriteback_0_bits_data_0 = 0x%0h ",pkt_str,this.io_exuWriteback_0_bits_data_0);
    pkt_str = $sformatf("%sio_exuWriteback_0_bits_robIdx_value = 0x%0h ",pkt_str,this.io_exuWriteback_0_bits_robIdx_value);
    pkt_str = $sformatf("%sio_writebackNums_0_bits = 0x%0h ",pkt_str,this.io_writebackNums_0_bits);
    pkt_str = $sformatf("%sio_writebackNums_1_bits = 0x%0h ",pkt_str,this.io_writebackNums_1_bits);
    pkt_str = $sformatf("%sio_writebackNums_2_bits = 0x%0h ",pkt_str,this.io_writebackNums_2_bits);
    pkt_str = $sformatf("%sio_writebackNums_3_bits = 0x%0h ",pkt_str,this.io_writebackNums_3_bits);
    pkt_str = $sformatf("%sio_writebackNums_4_bits = 0x%0h ",pkt_str,this.io_writebackNums_4_bits);
    pkt_str = $sformatf("%sio_writebackNums_5_bits = 0x%0h ",pkt_str,this.io_writebackNums_5_bits);
    pkt_str = $sformatf("%sio_writebackNums_6_bits = 0x%0h ",pkt_str,this.io_writebackNums_6_bits);
    pkt_str = $sformatf("%sio_writebackNums_7_bits = 0x%0h ",pkt_str,this.io_writebackNums_7_bits);
    pkt_str = $sformatf("%sio_writebackNums_8_bits = 0x%0h ",pkt_str,this.io_writebackNums_8_bits);
    pkt_str = $sformatf("%sio_writebackNums_9_bits = 0x%0h ",pkt_str,this.io_writebackNums_9_bits);
    pkt_str = $sformatf("%sio_writebackNums_10_bits = 0x%0h ",pkt_str,this.io_writebackNums_10_bits);
    pkt_str = $sformatf("%sio_writebackNums_11_bits = 0x%0h ",pkt_str,this.io_writebackNums_11_bits);
    pkt_str = $sformatf("%sio_writebackNums_12_bits = 0x%0h ",pkt_str,this.io_writebackNums_12_bits);
    pkt_str = $sformatf("%sio_writebackNums_13_bits = 0x%0h ",pkt_str,this.io_writebackNums_13_bits);
    pkt_str = $sformatf("%sio_writebackNums_14_bits = 0x%0h ",pkt_str,this.io_writebackNums_14_bits);
    pkt_str = $sformatf("%sio_writebackNums_15_bits = 0x%0h ",pkt_str,this.io_writebackNums_15_bits);
    pkt_str = $sformatf("%sio_writebackNums_16_bits = 0x%0h ",pkt_str,this.io_writebackNums_16_bits);
    pkt_str = $sformatf("%sio_writebackNums_17_bits = 0x%0h ",pkt_str,this.io_writebackNums_17_bits);
    pkt_str = $sformatf("%sio_writebackNums_18_bits = 0x%0h ",pkt_str,this.io_writebackNums_18_bits);
    pkt_str = $sformatf("%sio_writebackNums_19_bits = 0x%0h ",pkt_str,this.io_writebackNums_19_bits);
    pkt_str = $sformatf("%sio_writebackNums_20_bits = 0x%0h ",pkt_str,this.io_writebackNums_20_bits);
    pkt_str = $sformatf("%sio_writebackNums_21_bits = 0x%0h ",pkt_str,this.io_writebackNums_21_bits);
    pkt_str = $sformatf("%sio_writebackNums_22_bits = 0x%0h ",pkt_str,this.io_writebackNums_22_bits);
    pkt_str = $sformatf("%sio_writebackNums_23_bits = 0x%0h ",pkt_str,this.io_writebackNums_23_bits);
    pkt_str = $sformatf("%sio_writebackNums_24_bits = 0x%0h ",pkt_str,this.io_writebackNums_24_bits);
    pkt_str = $sformatf("%sio_writebackNeedFlush_0 = 0x%0h ",pkt_str,this.io_writebackNeedFlush_0);
    pkt_str = $sformatf("%sio_writebackNeedFlush_1 = 0x%0h ",pkt_str,this.io_writebackNeedFlush_1);
    pkt_str = $sformatf("%sio_writebackNeedFlush_2 = 0x%0h ",pkt_str,this.io_writebackNeedFlush_2);
    pkt_str = $sformatf("%sio_writebackNeedFlush_6 = 0x%0h ",pkt_str,this.io_writebackNeedFlush_6);
    pkt_str = $sformatf("%sio_writebackNeedFlush_7 = 0x%0h ",pkt_str,this.io_writebackNeedFlush_7);
    pkt_str = $sformatf("%sio_writebackNeedFlush_8 = 0x%0h ",pkt_str,this.io_writebackNeedFlush_8);
    pkt_str = $sformatf("%sio_writebackNeedFlush_9 = 0x%0h ",pkt_str,this.io_writebackNeedFlush_9);
    pkt_str = $sformatf("%sio_writebackNeedFlush_10 = 0x%0h ",pkt_str,this.io_writebackNeedFlush_10);
    pkt_str = $sformatf("%sio_writebackNeedFlush_11 = 0x%0h ",pkt_str,this.io_writebackNeedFlush_11);
    pkt_str = $sformatf("%sio_writebackNeedFlush_12 = 0x%0h ",pkt_str,this.io_writebackNeedFlush_12);

    return pkt_str;
endfunction:psdisplay

function bit WriteBack_in_agent_xaction::compare(uvm_object rhs, uvm_comparer comparer=null);
    bit super_result;
    WriteBack_in_agent_xaction  rhs_;
    if(!$cast(rhs_, rhs)) begin
        `uvm_fatal(get_type_name(),$sformatf("rhs is not a WriteBack_in_agent_xaction or its extend"))
    end
    super_result = super.compare(rhs_,comparer);
    if(super_result==0) begin
        super_result = 1;
        //foreach(this.pload_q[i]) begin
        //    if(this.pload_q[i]!=rhs_.pload_q[i]) begin
        //        super_result = 0;
        //        `uvm_info(get_type_name(),$sformatf("compare fail for this.pload[%0d]=0x%2h while the rhs_.pload[%0d]=0x%2h",i,this.pload_q[i],i,rhs_.pload_q[i]),UVM_NONE)
        //    end
        //end

        if(this.io_writeback_24_valid!=rhs_.io_writeback_24_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_valid=0x%0h while the rhs_.io_writeback_24_valid=0x%0h",this.io_writeback_24_valid,rhs_.io_writeback_24_valid),UVM_NONE)
        end

        if(this.io_writeback_24_bits_data_0!=rhs_.io_writeback_24_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_data_0=0x%0h while the rhs_.io_writeback_24_bits_data_0=0x%0h",this.io_writeback_24_bits_data_0,rhs_.io_writeback_24_bits_data_0),UVM_NONE)
        end

        if(this.io_writeback_24_bits_pdest!=rhs_.io_writeback_24_bits_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_pdest=0x%0h while the rhs_.io_writeback_24_bits_pdest=0x%0h",this.io_writeback_24_bits_pdest,rhs_.io_writeback_24_bits_pdest),UVM_NONE)
        end

        if(this.io_writeback_24_bits_robIdx_flag!=rhs_.io_writeback_24_bits_robIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_robIdx_flag=0x%0h while the rhs_.io_writeback_24_bits_robIdx_flag=0x%0h",this.io_writeback_24_bits_robIdx_flag,rhs_.io_writeback_24_bits_robIdx_flag),UVM_NONE)
        end

        if(this.io_writeback_24_bits_robIdx_value!=rhs_.io_writeback_24_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_robIdx_value=0x%0h while the rhs_.io_writeback_24_bits_robIdx_value=0x%0h",this.io_writeback_24_bits_robIdx_value,rhs_.io_writeback_24_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vecWen!=rhs_.io_writeback_24_bits_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vecWen=0x%0h while the rhs_.io_writeback_24_bits_vecWen=0x%0h",this.io_writeback_24_bits_vecWen,rhs_.io_writeback_24_bits_vecWen),UVM_NONE)
        end

        if(this.io_writeback_24_bits_v0Wen!=rhs_.io_writeback_24_bits_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_v0Wen=0x%0h while the rhs_.io_writeback_24_bits_v0Wen=0x%0h",this.io_writeback_24_bits_v0Wen,rhs_.io_writeback_24_bits_v0Wen),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vlWen!=rhs_.io_writeback_24_bits_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vlWen=0x%0h while the rhs_.io_writeback_24_bits_vlWen=0x%0h",this.io_writeback_24_bits_vlWen,rhs_.io_writeback_24_bits_vlWen),UVM_NONE)
        end

        if(this.io_writeback_24_bits_exceptionVec_0!=rhs_.io_writeback_24_bits_exceptionVec_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_exceptionVec_0=0x%0h while the rhs_.io_writeback_24_bits_exceptionVec_0=0x%0h",this.io_writeback_24_bits_exceptionVec_0,rhs_.io_writeback_24_bits_exceptionVec_0),UVM_NONE)
        end

        if(this.io_writeback_24_bits_exceptionVec_1!=rhs_.io_writeback_24_bits_exceptionVec_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_exceptionVec_1=0x%0h while the rhs_.io_writeback_24_bits_exceptionVec_1=0x%0h",this.io_writeback_24_bits_exceptionVec_1,rhs_.io_writeback_24_bits_exceptionVec_1),UVM_NONE)
        end

        if(this.io_writeback_24_bits_exceptionVec_2!=rhs_.io_writeback_24_bits_exceptionVec_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_exceptionVec_2=0x%0h while the rhs_.io_writeback_24_bits_exceptionVec_2=0x%0h",this.io_writeback_24_bits_exceptionVec_2,rhs_.io_writeback_24_bits_exceptionVec_2),UVM_NONE)
        end

        if(this.io_writeback_24_bits_exceptionVec_3!=rhs_.io_writeback_24_bits_exceptionVec_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_exceptionVec_3=0x%0h while the rhs_.io_writeback_24_bits_exceptionVec_3=0x%0h",this.io_writeback_24_bits_exceptionVec_3,rhs_.io_writeback_24_bits_exceptionVec_3),UVM_NONE)
        end

        if(this.io_writeback_24_bits_exceptionVec_4!=rhs_.io_writeback_24_bits_exceptionVec_4) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_exceptionVec_4=0x%0h while the rhs_.io_writeback_24_bits_exceptionVec_4=0x%0h",this.io_writeback_24_bits_exceptionVec_4,rhs_.io_writeback_24_bits_exceptionVec_4),UVM_NONE)
        end

        if(this.io_writeback_24_bits_exceptionVec_5!=rhs_.io_writeback_24_bits_exceptionVec_5) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_exceptionVec_5=0x%0h while the rhs_.io_writeback_24_bits_exceptionVec_5=0x%0h",this.io_writeback_24_bits_exceptionVec_5,rhs_.io_writeback_24_bits_exceptionVec_5),UVM_NONE)
        end

        if(this.io_writeback_24_bits_exceptionVec_6!=rhs_.io_writeback_24_bits_exceptionVec_6) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_exceptionVec_6=0x%0h while the rhs_.io_writeback_24_bits_exceptionVec_6=0x%0h",this.io_writeback_24_bits_exceptionVec_6,rhs_.io_writeback_24_bits_exceptionVec_6),UVM_NONE)
        end

        if(this.io_writeback_24_bits_exceptionVec_7!=rhs_.io_writeback_24_bits_exceptionVec_7) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_exceptionVec_7=0x%0h while the rhs_.io_writeback_24_bits_exceptionVec_7=0x%0h",this.io_writeback_24_bits_exceptionVec_7,rhs_.io_writeback_24_bits_exceptionVec_7),UVM_NONE)
        end

        if(this.io_writeback_24_bits_exceptionVec_8!=rhs_.io_writeback_24_bits_exceptionVec_8) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_exceptionVec_8=0x%0h while the rhs_.io_writeback_24_bits_exceptionVec_8=0x%0h",this.io_writeback_24_bits_exceptionVec_8,rhs_.io_writeback_24_bits_exceptionVec_8),UVM_NONE)
        end

        if(this.io_writeback_24_bits_exceptionVec_9!=rhs_.io_writeback_24_bits_exceptionVec_9) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_exceptionVec_9=0x%0h while the rhs_.io_writeback_24_bits_exceptionVec_9=0x%0h",this.io_writeback_24_bits_exceptionVec_9,rhs_.io_writeback_24_bits_exceptionVec_9),UVM_NONE)
        end

        if(this.io_writeback_24_bits_exceptionVec_10!=rhs_.io_writeback_24_bits_exceptionVec_10) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_exceptionVec_10=0x%0h while the rhs_.io_writeback_24_bits_exceptionVec_10=0x%0h",this.io_writeback_24_bits_exceptionVec_10,rhs_.io_writeback_24_bits_exceptionVec_10),UVM_NONE)
        end

        if(this.io_writeback_24_bits_exceptionVec_11!=rhs_.io_writeback_24_bits_exceptionVec_11) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_exceptionVec_11=0x%0h while the rhs_.io_writeback_24_bits_exceptionVec_11=0x%0h",this.io_writeback_24_bits_exceptionVec_11,rhs_.io_writeback_24_bits_exceptionVec_11),UVM_NONE)
        end

        if(this.io_writeback_24_bits_exceptionVec_12!=rhs_.io_writeback_24_bits_exceptionVec_12) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_exceptionVec_12=0x%0h while the rhs_.io_writeback_24_bits_exceptionVec_12=0x%0h",this.io_writeback_24_bits_exceptionVec_12,rhs_.io_writeback_24_bits_exceptionVec_12),UVM_NONE)
        end

        if(this.io_writeback_24_bits_exceptionVec_13!=rhs_.io_writeback_24_bits_exceptionVec_13) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_exceptionVec_13=0x%0h while the rhs_.io_writeback_24_bits_exceptionVec_13=0x%0h",this.io_writeback_24_bits_exceptionVec_13,rhs_.io_writeback_24_bits_exceptionVec_13),UVM_NONE)
        end

        if(this.io_writeback_24_bits_exceptionVec_14!=rhs_.io_writeback_24_bits_exceptionVec_14) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_exceptionVec_14=0x%0h while the rhs_.io_writeback_24_bits_exceptionVec_14=0x%0h",this.io_writeback_24_bits_exceptionVec_14,rhs_.io_writeback_24_bits_exceptionVec_14),UVM_NONE)
        end

        if(this.io_writeback_24_bits_exceptionVec_15!=rhs_.io_writeback_24_bits_exceptionVec_15) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_exceptionVec_15=0x%0h while the rhs_.io_writeback_24_bits_exceptionVec_15=0x%0h",this.io_writeback_24_bits_exceptionVec_15,rhs_.io_writeback_24_bits_exceptionVec_15),UVM_NONE)
        end

        if(this.io_writeback_24_bits_exceptionVec_16!=rhs_.io_writeback_24_bits_exceptionVec_16) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_exceptionVec_16=0x%0h while the rhs_.io_writeback_24_bits_exceptionVec_16=0x%0h",this.io_writeback_24_bits_exceptionVec_16,rhs_.io_writeback_24_bits_exceptionVec_16),UVM_NONE)
        end

        if(this.io_writeback_24_bits_exceptionVec_17!=rhs_.io_writeback_24_bits_exceptionVec_17) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_exceptionVec_17=0x%0h while the rhs_.io_writeback_24_bits_exceptionVec_17=0x%0h",this.io_writeback_24_bits_exceptionVec_17,rhs_.io_writeback_24_bits_exceptionVec_17),UVM_NONE)
        end

        if(this.io_writeback_24_bits_exceptionVec_18!=rhs_.io_writeback_24_bits_exceptionVec_18) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_exceptionVec_18=0x%0h while the rhs_.io_writeback_24_bits_exceptionVec_18=0x%0h",this.io_writeback_24_bits_exceptionVec_18,rhs_.io_writeback_24_bits_exceptionVec_18),UVM_NONE)
        end

        if(this.io_writeback_24_bits_exceptionVec_19!=rhs_.io_writeback_24_bits_exceptionVec_19) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_exceptionVec_19=0x%0h while the rhs_.io_writeback_24_bits_exceptionVec_19=0x%0h",this.io_writeback_24_bits_exceptionVec_19,rhs_.io_writeback_24_bits_exceptionVec_19),UVM_NONE)
        end

        if(this.io_writeback_24_bits_exceptionVec_20!=rhs_.io_writeback_24_bits_exceptionVec_20) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_exceptionVec_20=0x%0h while the rhs_.io_writeback_24_bits_exceptionVec_20=0x%0h",this.io_writeback_24_bits_exceptionVec_20,rhs_.io_writeback_24_bits_exceptionVec_20),UVM_NONE)
        end

        if(this.io_writeback_24_bits_exceptionVec_21!=rhs_.io_writeback_24_bits_exceptionVec_21) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_exceptionVec_21=0x%0h while the rhs_.io_writeback_24_bits_exceptionVec_21=0x%0h",this.io_writeback_24_bits_exceptionVec_21,rhs_.io_writeback_24_bits_exceptionVec_21),UVM_NONE)
        end

        if(this.io_writeback_24_bits_exceptionVec_22!=rhs_.io_writeback_24_bits_exceptionVec_22) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_exceptionVec_22=0x%0h while the rhs_.io_writeback_24_bits_exceptionVec_22=0x%0h",this.io_writeback_24_bits_exceptionVec_22,rhs_.io_writeback_24_bits_exceptionVec_22),UVM_NONE)
        end

        if(this.io_writeback_24_bits_exceptionVec_23!=rhs_.io_writeback_24_bits_exceptionVec_23) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_exceptionVec_23=0x%0h while the rhs_.io_writeback_24_bits_exceptionVec_23=0x%0h",this.io_writeback_24_bits_exceptionVec_23,rhs_.io_writeback_24_bits_exceptionVec_23),UVM_NONE)
        end

        if(this.io_writeback_24_bits_flushPipe!=rhs_.io_writeback_24_bits_flushPipe) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_flushPipe=0x%0h while the rhs_.io_writeback_24_bits_flushPipe=0x%0h",this.io_writeback_24_bits_flushPipe,rhs_.io_writeback_24_bits_flushPipe),UVM_NONE)
        end

        if(this.io_writeback_24_bits_replay!=rhs_.io_writeback_24_bits_replay) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_replay=0x%0h while the rhs_.io_writeback_24_bits_replay=0x%0h",this.io_writeback_24_bits_replay,rhs_.io_writeback_24_bits_replay),UVM_NONE)
        end

        if(this.io_writeback_24_bits_trigger!=rhs_.io_writeback_24_bits_trigger) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_trigger=0x%0h while the rhs_.io_writeback_24_bits_trigger=0x%0h",this.io_writeback_24_bits_trigger,rhs_.io_writeback_24_bits_trigger),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_vill!=rhs_.io_writeback_24_bits_vls_vpu_vill) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_vill=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_vill=0x%0h",this.io_writeback_24_bits_vls_vpu_vill,rhs_.io_writeback_24_bits_vls_vpu_vill),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_vma!=rhs_.io_writeback_24_bits_vls_vpu_vma) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_vma=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_vma=0x%0h",this.io_writeback_24_bits_vls_vpu_vma,rhs_.io_writeback_24_bits_vls_vpu_vma),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_vta!=rhs_.io_writeback_24_bits_vls_vpu_vta) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_vta=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_vta=0x%0h",this.io_writeback_24_bits_vls_vpu_vta,rhs_.io_writeback_24_bits_vls_vpu_vta),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_vsew!=rhs_.io_writeback_24_bits_vls_vpu_vsew) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_vsew=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_vsew=0x%0h",this.io_writeback_24_bits_vls_vpu_vsew,rhs_.io_writeback_24_bits_vls_vpu_vsew),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_vlmul!=rhs_.io_writeback_24_bits_vls_vpu_vlmul) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_vlmul=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_vlmul=0x%0h",this.io_writeback_24_bits_vls_vpu_vlmul,rhs_.io_writeback_24_bits_vls_vpu_vlmul),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_specVill!=rhs_.io_writeback_24_bits_vls_vpu_specVill) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_specVill=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_specVill=0x%0h",this.io_writeback_24_bits_vls_vpu_specVill,rhs_.io_writeback_24_bits_vls_vpu_specVill),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_specVma!=rhs_.io_writeback_24_bits_vls_vpu_specVma) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_specVma=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_specVma=0x%0h",this.io_writeback_24_bits_vls_vpu_specVma,rhs_.io_writeback_24_bits_vls_vpu_specVma),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_specVta!=rhs_.io_writeback_24_bits_vls_vpu_specVta) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_specVta=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_specVta=0x%0h",this.io_writeback_24_bits_vls_vpu_specVta,rhs_.io_writeback_24_bits_vls_vpu_specVta),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_specVsew!=rhs_.io_writeback_24_bits_vls_vpu_specVsew) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_specVsew=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_specVsew=0x%0h",this.io_writeback_24_bits_vls_vpu_specVsew,rhs_.io_writeback_24_bits_vls_vpu_specVsew),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_specVlmul!=rhs_.io_writeback_24_bits_vls_vpu_specVlmul) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_specVlmul=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_specVlmul=0x%0h",this.io_writeback_24_bits_vls_vpu_specVlmul,rhs_.io_writeback_24_bits_vls_vpu_specVlmul),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_vm!=rhs_.io_writeback_24_bits_vls_vpu_vm) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_vm=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_vm=0x%0h",this.io_writeback_24_bits_vls_vpu_vm,rhs_.io_writeback_24_bits_vls_vpu_vm),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_vstart!=rhs_.io_writeback_24_bits_vls_vpu_vstart) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_vstart=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_vstart=0x%0h",this.io_writeback_24_bits_vls_vpu_vstart,rhs_.io_writeback_24_bits_vls_vpu_vstart),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_frm!=rhs_.io_writeback_24_bits_vls_vpu_frm) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_frm=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_frm=0x%0h",this.io_writeback_24_bits_vls_vpu_frm,rhs_.io_writeback_24_bits_vls_vpu_frm),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst!=rhs_.io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst=0x%0h",this.io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst,rhs_.io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_fpu_isFP32Instr!=rhs_.io_writeback_24_bits_vls_vpu_fpu_isFP32Instr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_fpu_isFP32Instr=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_fpu_isFP32Instr=0x%0h",this.io_writeback_24_bits_vls_vpu_fpu_isFP32Instr,rhs_.io_writeback_24_bits_vls_vpu_fpu_isFP32Instr),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_fpu_isFP64Instr!=rhs_.io_writeback_24_bits_vls_vpu_fpu_isFP64Instr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_fpu_isFP64Instr=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_fpu_isFP64Instr=0x%0h",this.io_writeback_24_bits_vls_vpu_fpu_isFP64Instr,rhs_.io_writeback_24_bits_vls_vpu_fpu_isFP64Instr),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_fpu_isReduction!=rhs_.io_writeback_24_bits_vls_vpu_fpu_isReduction) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_fpu_isReduction=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_fpu_isReduction=0x%0h",this.io_writeback_24_bits_vls_vpu_fpu_isReduction,rhs_.io_writeback_24_bits_vls_vpu_fpu_isReduction),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2!=rhs_.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2=0x%0h",this.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2,rhs_.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4!=rhs_.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4=0x%0h",this.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4,rhs_.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8!=rhs_.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8=0x%0h",this.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8,rhs_.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_vxrm!=rhs_.io_writeback_24_bits_vls_vpu_vxrm) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_vxrm=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_vxrm=0x%0h",this.io_writeback_24_bits_vls_vpu_vxrm,rhs_.io_writeback_24_bits_vls_vpu_vxrm),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_vuopIdx!=rhs_.io_writeback_24_bits_vls_vpu_vuopIdx) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_vuopIdx=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_vuopIdx=0x%0h",this.io_writeback_24_bits_vls_vpu_vuopIdx,rhs_.io_writeback_24_bits_vls_vpu_vuopIdx),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_lastUop!=rhs_.io_writeback_24_bits_vls_vpu_lastUop) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_lastUop=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_lastUop=0x%0h",this.io_writeback_24_bits_vls_vpu_lastUop,rhs_.io_writeback_24_bits_vls_vpu_lastUop),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_vmask!=rhs_.io_writeback_24_bits_vls_vpu_vmask) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_vmask=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_vmask=0x%0h",this.io_writeback_24_bits_vls_vpu_vmask,rhs_.io_writeback_24_bits_vls_vpu_vmask),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_vl!=rhs_.io_writeback_24_bits_vls_vpu_vl) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_vl=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_vl=0x%0h",this.io_writeback_24_bits_vls_vpu_vl,rhs_.io_writeback_24_bits_vls_vpu_vl),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_nf!=rhs_.io_writeback_24_bits_vls_vpu_nf) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_nf=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_nf=0x%0h",this.io_writeback_24_bits_vls_vpu_nf,rhs_.io_writeback_24_bits_vls_vpu_nf),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_veew!=rhs_.io_writeback_24_bits_vls_vpu_veew) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_veew=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_veew=0x%0h",this.io_writeback_24_bits_vls_vpu_veew,rhs_.io_writeback_24_bits_vls_vpu_veew),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_isReverse!=rhs_.io_writeback_24_bits_vls_vpu_isReverse) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_isReverse=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_isReverse=0x%0h",this.io_writeback_24_bits_vls_vpu_isReverse,rhs_.io_writeback_24_bits_vls_vpu_isReverse),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_isExt!=rhs_.io_writeback_24_bits_vls_vpu_isExt) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_isExt=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_isExt=0x%0h",this.io_writeback_24_bits_vls_vpu_isExt,rhs_.io_writeback_24_bits_vls_vpu_isExt),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_isNarrow!=rhs_.io_writeback_24_bits_vls_vpu_isNarrow) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_isNarrow=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_isNarrow=0x%0h",this.io_writeback_24_bits_vls_vpu_isNarrow,rhs_.io_writeback_24_bits_vls_vpu_isNarrow),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_isDstMask!=rhs_.io_writeback_24_bits_vls_vpu_isDstMask) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_isDstMask=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_isDstMask=0x%0h",this.io_writeback_24_bits_vls_vpu_isDstMask,rhs_.io_writeback_24_bits_vls_vpu_isDstMask),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_isOpMask!=rhs_.io_writeback_24_bits_vls_vpu_isOpMask) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_isOpMask=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_isOpMask=0x%0h",this.io_writeback_24_bits_vls_vpu_isOpMask,rhs_.io_writeback_24_bits_vls_vpu_isOpMask),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_isMove!=rhs_.io_writeback_24_bits_vls_vpu_isMove) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_isMove=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_isMove=0x%0h",this.io_writeback_24_bits_vls_vpu_isMove,rhs_.io_writeback_24_bits_vls_vpu_isMove),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_isDependOldVd!=rhs_.io_writeback_24_bits_vls_vpu_isDependOldVd) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_isDependOldVd=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_isDependOldVd=0x%0h",this.io_writeback_24_bits_vls_vpu_isDependOldVd,rhs_.io_writeback_24_bits_vls_vpu_isDependOldVd),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_isWritePartVd!=rhs_.io_writeback_24_bits_vls_vpu_isWritePartVd) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_isWritePartVd=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_isWritePartVd=0x%0h",this.io_writeback_24_bits_vls_vpu_isWritePartVd,rhs_.io_writeback_24_bits_vls_vpu_isWritePartVd),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vpu_isVleff!=rhs_.io_writeback_24_bits_vls_vpu_isVleff) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vpu_isVleff=0x%0h while the rhs_.io_writeback_24_bits_vls_vpu_isVleff=0x%0h",this.io_writeback_24_bits_vls_vpu_isVleff,rhs_.io_writeback_24_bits_vls_vpu_isVleff),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_oldVdPsrc!=rhs_.io_writeback_24_bits_vls_oldVdPsrc) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_oldVdPsrc=0x%0h while the rhs_.io_writeback_24_bits_vls_oldVdPsrc=0x%0h",this.io_writeback_24_bits_vls_oldVdPsrc,rhs_.io_writeback_24_bits_vls_oldVdPsrc),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vdIdx!=rhs_.io_writeback_24_bits_vls_vdIdx) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vdIdx=0x%0h while the rhs_.io_writeback_24_bits_vls_vdIdx=0x%0h",this.io_writeback_24_bits_vls_vdIdx,rhs_.io_writeback_24_bits_vls_vdIdx),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_vdIdxInField!=rhs_.io_writeback_24_bits_vls_vdIdxInField) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_vdIdxInField=0x%0h while the rhs_.io_writeback_24_bits_vls_vdIdxInField=0x%0h",this.io_writeback_24_bits_vls_vdIdxInField,rhs_.io_writeback_24_bits_vls_vdIdxInField),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_isIndexed!=rhs_.io_writeback_24_bits_vls_isIndexed) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_isIndexed=0x%0h while the rhs_.io_writeback_24_bits_vls_isIndexed=0x%0h",this.io_writeback_24_bits_vls_isIndexed,rhs_.io_writeback_24_bits_vls_isIndexed),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_isMasked!=rhs_.io_writeback_24_bits_vls_isMasked) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_isMasked=0x%0h while the rhs_.io_writeback_24_bits_vls_isMasked=0x%0h",this.io_writeback_24_bits_vls_isMasked,rhs_.io_writeback_24_bits_vls_isMasked),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_isStrided!=rhs_.io_writeback_24_bits_vls_isStrided) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_isStrided=0x%0h while the rhs_.io_writeback_24_bits_vls_isStrided=0x%0h",this.io_writeback_24_bits_vls_isStrided,rhs_.io_writeback_24_bits_vls_isStrided),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_isWhole!=rhs_.io_writeback_24_bits_vls_isWhole) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_isWhole=0x%0h while the rhs_.io_writeback_24_bits_vls_isWhole=0x%0h",this.io_writeback_24_bits_vls_isWhole,rhs_.io_writeback_24_bits_vls_isWhole),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_isVecLoad!=rhs_.io_writeback_24_bits_vls_isVecLoad) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_isVecLoad=0x%0h while the rhs_.io_writeback_24_bits_vls_isVecLoad=0x%0h",this.io_writeback_24_bits_vls_isVecLoad,rhs_.io_writeback_24_bits_vls_isVecLoad),UVM_NONE)
        end

        if(this.io_writeback_24_bits_vls_isVlm!=rhs_.io_writeback_24_bits_vls_isVlm) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_vls_isVlm=0x%0h while the rhs_.io_writeback_24_bits_vls_isVlm=0x%0h",this.io_writeback_24_bits_vls_isVlm,rhs_.io_writeback_24_bits_vls_isVlm),UVM_NONE)
        end

        if(this.io_writeback_24_bits_debug_isMMIO!=rhs_.io_writeback_24_bits_debug_isMMIO) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_debug_isMMIO=0x%0h while the rhs_.io_writeback_24_bits_debug_isMMIO=0x%0h",this.io_writeback_24_bits_debug_isMMIO,rhs_.io_writeback_24_bits_debug_isMMIO),UVM_NONE)
        end

        if(this.io_writeback_24_bits_debug_isNCIO!=rhs_.io_writeback_24_bits_debug_isNCIO) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_debug_isNCIO=0x%0h while the rhs_.io_writeback_24_bits_debug_isNCIO=0x%0h",this.io_writeback_24_bits_debug_isNCIO,rhs_.io_writeback_24_bits_debug_isNCIO),UVM_NONE)
        end

        if(this.io_writeback_24_bits_debug_isPerfCnt!=rhs_.io_writeback_24_bits_debug_isPerfCnt) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_debug_isPerfCnt=0x%0h while the rhs_.io_writeback_24_bits_debug_isPerfCnt=0x%0h",this.io_writeback_24_bits_debug_isPerfCnt,rhs_.io_writeback_24_bits_debug_isPerfCnt),UVM_NONE)
        end

        if(this.io_writeback_24_bits_debug_paddr!=rhs_.io_writeback_24_bits_debug_paddr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_debug_paddr=0x%0h while the rhs_.io_writeback_24_bits_debug_paddr=0x%0h",this.io_writeback_24_bits_debug_paddr,rhs_.io_writeback_24_bits_debug_paddr),UVM_NONE)
        end

        if(this.io_writeback_24_bits_debug_vaddr!=rhs_.io_writeback_24_bits_debug_vaddr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_debug_vaddr=0x%0h while the rhs_.io_writeback_24_bits_debug_vaddr=0x%0h",this.io_writeback_24_bits_debug_vaddr,rhs_.io_writeback_24_bits_debug_vaddr),UVM_NONE)
        end

        if(this.io_writeback_24_bits_debugInfo_eliminatedMove!=rhs_.io_writeback_24_bits_debugInfo_eliminatedMove) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_debugInfo_eliminatedMove=0x%0h while the rhs_.io_writeback_24_bits_debugInfo_eliminatedMove=0x%0h",this.io_writeback_24_bits_debugInfo_eliminatedMove,rhs_.io_writeback_24_bits_debugInfo_eliminatedMove),UVM_NONE)
        end

        if(this.io_writeback_24_bits_debugInfo_renameTime!=rhs_.io_writeback_24_bits_debugInfo_renameTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_debugInfo_renameTime=0x%0h while the rhs_.io_writeback_24_bits_debugInfo_renameTime=0x%0h",this.io_writeback_24_bits_debugInfo_renameTime,rhs_.io_writeback_24_bits_debugInfo_renameTime),UVM_NONE)
        end

        if(this.io_writeback_24_bits_debugInfo_dispatchTime!=rhs_.io_writeback_24_bits_debugInfo_dispatchTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_debugInfo_dispatchTime=0x%0h while the rhs_.io_writeback_24_bits_debugInfo_dispatchTime=0x%0h",this.io_writeback_24_bits_debugInfo_dispatchTime,rhs_.io_writeback_24_bits_debugInfo_dispatchTime),UVM_NONE)
        end

        if(this.io_writeback_24_bits_debugInfo_enqRsTime!=rhs_.io_writeback_24_bits_debugInfo_enqRsTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_debugInfo_enqRsTime=0x%0h while the rhs_.io_writeback_24_bits_debugInfo_enqRsTime=0x%0h",this.io_writeback_24_bits_debugInfo_enqRsTime,rhs_.io_writeback_24_bits_debugInfo_enqRsTime),UVM_NONE)
        end

        if(this.io_writeback_24_bits_debugInfo_selectTime!=rhs_.io_writeback_24_bits_debugInfo_selectTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_debugInfo_selectTime=0x%0h while the rhs_.io_writeback_24_bits_debugInfo_selectTime=0x%0h",this.io_writeback_24_bits_debugInfo_selectTime,rhs_.io_writeback_24_bits_debugInfo_selectTime),UVM_NONE)
        end

        if(this.io_writeback_24_bits_debugInfo_issueTime!=rhs_.io_writeback_24_bits_debugInfo_issueTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_debugInfo_issueTime=0x%0h while the rhs_.io_writeback_24_bits_debugInfo_issueTime=0x%0h",this.io_writeback_24_bits_debugInfo_issueTime,rhs_.io_writeback_24_bits_debugInfo_issueTime),UVM_NONE)
        end

        if(this.io_writeback_24_bits_debugInfo_writebackTime!=rhs_.io_writeback_24_bits_debugInfo_writebackTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_debugInfo_writebackTime=0x%0h while the rhs_.io_writeback_24_bits_debugInfo_writebackTime=0x%0h",this.io_writeback_24_bits_debugInfo_writebackTime,rhs_.io_writeback_24_bits_debugInfo_writebackTime),UVM_NONE)
        end

        if(this.io_writeback_24_bits_debugInfo_runahead_checkpoint_id!=rhs_.io_writeback_24_bits_debugInfo_runahead_checkpoint_id) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_debugInfo_runahead_checkpoint_id=0x%0h while the rhs_.io_writeback_24_bits_debugInfo_runahead_checkpoint_id=0x%0h",this.io_writeback_24_bits_debugInfo_runahead_checkpoint_id,rhs_.io_writeback_24_bits_debugInfo_runahead_checkpoint_id),UVM_NONE)
        end

        if(this.io_writeback_24_bits_debugInfo_tlbFirstReqTime!=rhs_.io_writeback_24_bits_debugInfo_tlbFirstReqTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_debugInfo_tlbFirstReqTime=0x%0h while the rhs_.io_writeback_24_bits_debugInfo_tlbFirstReqTime=0x%0h",this.io_writeback_24_bits_debugInfo_tlbFirstReqTime,rhs_.io_writeback_24_bits_debugInfo_tlbFirstReqTime),UVM_NONE)
        end

        if(this.io_writeback_24_bits_debugInfo_tlbRespTime!=rhs_.io_writeback_24_bits_debugInfo_tlbRespTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_debugInfo_tlbRespTime=0x%0h while the rhs_.io_writeback_24_bits_debugInfo_tlbRespTime=0x%0h",this.io_writeback_24_bits_debugInfo_tlbRespTime,rhs_.io_writeback_24_bits_debugInfo_tlbRespTime),UVM_NONE)
        end

        if(this.io_writeback_24_bits_debug_seqNum!=rhs_.io_writeback_24_bits_debug_seqNum) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_24_bits_debug_seqNum=0x%0h while the rhs_.io_writeback_24_bits_debug_seqNum=0x%0h",this.io_writeback_24_bits_debug_seqNum,rhs_.io_writeback_24_bits_debug_seqNum),UVM_NONE)
        end

        if(this.io_writeback_23_valid!=rhs_.io_writeback_23_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_valid=0x%0h while the rhs_.io_writeback_23_valid=0x%0h",this.io_writeback_23_valid,rhs_.io_writeback_23_valid),UVM_NONE)
        end

        if(this.io_writeback_23_bits_data_0!=rhs_.io_writeback_23_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_data_0=0x%0h while the rhs_.io_writeback_23_bits_data_0=0x%0h",this.io_writeback_23_bits_data_0,rhs_.io_writeback_23_bits_data_0),UVM_NONE)
        end

        if(this.io_writeback_23_bits_pdest!=rhs_.io_writeback_23_bits_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_pdest=0x%0h while the rhs_.io_writeback_23_bits_pdest=0x%0h",this.io_writeback_23_bits_pdest,rhs_.io_writeback_23_bits_pdest),UVM_NONE)
        end

        if(this.io_writeback_23_bits_robIdx_flag!=rhs_.io_writeback_23_bits_robIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_robIdx_flag=0x%0h while the rhs_.io_writeback_23_bits_robIdx_flag=0x%0h",this.io_writeback_23_bits_robIdx_flag,rhs_.io_writeback_23_bits_robIdx_flag),UVM_NONE)
        end

        if(this.io_writeback_23_bits_robIdx_value!=rhs_.io_writeback_23_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_robIdx_value=0x%0h while the rhs_.io_writeback_23_bits_robIdx_value=0x%0h",this.io_writeback_23_bits_robIdx_value,rhs_.io_writeback_23_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vecWen!=rhs_.io_writeback_23_bits_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vecWen=0x%0h while the rhs_.io_writeback_23_bits_vecWen=0x%0h",this.io_writeback_23_bits_vecWen,rhs_.io_writeback_23_bits_vecWen),UVM_NONE)
        end

        if(this.io_writeback_23_bits_v0Wen!=rhs_.io_writeback_23_bits_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_v0Wen=0x%0h while the rhs_.io_writeback_23_bits_v0Wen=0x%0h",this.io_writeback_23_bits_v0Wen,rhs_.io_writeback_23_bits_v0Wen),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vlWen!=rhs_.io_writeback_23_bits_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vlWen=0x%0h while the rhs_.io_writeback_23_bits_vlWen=0x%0h",this.io_writeback_23_bits_vlWen,rhs_.io_writeback_23_bits_vlWen),UVM_NONE)
        end

        if(this.io_writeback_23_bits_exceptionVec_0!=rhs_.io_writeback_23_bits_exceptionVec_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_exceptionVec_0=0x%0h while the rhs_.io_writeback_23_bits_exceptionVec_0=0x%0h",this.io_writeback_23_bits_exceptionVec_0,rhs_.io_writeback_23_bits_exceptionVec_0),UVM_NONE)
        end

        if(this.io_writeback_23_bits_exceptionVec_1!=rhs_.io_writeback_23_bits_exceptionVec_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_exceptionVec_1=0x%0h while the rhs_.io_writeback_23_bits_exceptionVec_1=0x%0h",this.io_writeback_23_bits_exceptionVec_1,rhs_.io_writeback_23_bits_exceptionVec_1),UVM_NONE)
        end

        if(this.io_writeback_23_bits_exceptionVec_2!=rhs_.io_writeback_23_bits_exceptionVec_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_exceptionVec_2=0x%0h while the rhs_.io_writeback_23_bits_exceptionVec_2=0x%0h",this.io_writeback_23_bits_exceptionVec_2,rhs_.io_writeback_23_bits_exceptionVec_2),UVM_NONE)
        end

        if(this.io_writeback_23_bits_exceptionVec_3!=rhs_.io_writeback_23_bits_exceptionVec_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_exceptionVec_3=0x%0h while the rhs_.io_writeback_23_bits_exceptionVec_3=0x%0h",this.io_writeback_23_bits_exceptionVec_3,rhs_.io_writeback_23_bits_exceptionVec_3),UVM_NONE)
        end

        if(this.io_writeback_23_bits_exceptionVec_4!=rhs_.io_writeback_23_bits_exceptionVec_4) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_exceptionVec_4=0x%0h while the rhs_.io_writeback_23_bits_exceptionVec_4=0x%0h",this.io_writeback_23_bits_exceptionVec_4,rhs_.io_writeback_23_bits_exceptionVec_4),UVM_NONE)
        end

        if(this.io_writeback_23_bits_exceptionVec_5!=rhs_.io_writeback_23_bits_exceptionVec_5) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_exceptionVec_5=0x%0h while the rhs_.io_writeback_23_bits_exceptionVec_5=0x%0h",this.io_writeback_23_bits_exceptionVec_5,rhs_.io_writeback_23_bits_exceptionVec_5),UVM_NONE)
        end

        if(this.io_writeback_23_bits_exceptionVec_6!=rhs_.io_writeback_23_bits_exceptionVec_6) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_exceptionVec_6=0x%0h while the rhs_.io_writeback_23_bits_exceptionVec_6=0x%0h",this.io_writeback_23_bits_exceptionVec_6,rhs_.io_writeback_23_bits_exceptionVec_6),UVM_NONE)
        end

        if(this.io_writeback_23_bits_exceptionVec_7!=rhs_.io_writeback_23_bits_exceptionVec_7) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_exceptionVec_7=0x%0h while the rhs_.io_writeback_23_bits_exceptionVec_7=0x%0h",this.io_writeback_23_bits_exceptionVec_7,rhs_.io_writeback_23_bits_exceptionVec_7),UVM_NONE)
        end

        if(this.io_writeback_23_bits_exceptionVec_8!=rhs_.io_writeback_23_bits_exceptionVec_8) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_exceptionVec_8=0x%0h while the rhs_.io_writeback_23_bits_exceptionVec_8=0x%0h",this.io_writeback_23_bits_exceptionVec_8,rhs_.io_writeback_23_bits_exceptionVec_8),UVM_NONE)
        end

        if(this.io_writeback_23_bits_exceptionVec_9!=rhs_.io_writeback_23_bits_exceptionVec_9) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_exceptionVec_9=0x%0h while the rhs_.io_writeback_23_bits_exceptionVec_9=0x%0h",this.io_writeback_23_bits_exceptionVec_9,rhs_.io_writeback_23_bits_exceptionVec_9),UVM_NONE)
        end

        if(this.io_writeback_23_bits_exceptionVec_10!=rhs_.io_writeback_23_bits_exceptionVec_10) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_exceptionVec_10=0x%0h while the rhs_.io_writeback_23_bits_exceptionVec_10=0x%0h",this.io_writeback_23_bits_exceptionVec_10,rhs_.io_writeback_23_bits_exceptionVec_10),UVM_NONE)
        end

        if(this.io_writeback_23_bits_exceptionVec_11!=rhs_.io_writeback_23_bits_exceptionVec_11) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_exceptionVec_11=0x%0h while the rhs_.io_writeback_23_bits_exceptionVec_11=0x%0h",this.io_writeback_23_bits_exceptionVec_11,rhs_.io_writeback_23_bits_exceptionVec_11),UVM_NONE)
        end

        if(this.io_writeback_23_bits_exceptionVec_12!=rhs_.io_writeback_23_bits_exceptionVec_12) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_exceptionVec_12=0x%0h while the rhs_.io_writeback_23_bits_exceptionVec_12=0x%0h",this.io_writeback_23_bits_exceptionVec_12,rhs_.io_writeback_23_bits_exceptionVec_12),UVM_NONE)
        end

        if(this.io_writeback_23_bits_exceptionVec_13!=rhs_.io_writeback_23_bits_exceptionVec_13) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_exceptionVec_13=0x%0h while the rhs_.io_writeback_23_bits_exceptionVec_13=0x%0h",this.io_writeback_23_bits_exceptionVec_13,rhs_.io_writeback_23_bits_exceptionVec_13),UVM_NONE)
        end

        if(this.io_writeback_23_bits_exceptionVec_14!=rhs_.io_writeback_23_bits_exceptionVec_14) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_exceptionVec_14=0x%0h while the rhs_.io_writeback_23_bits_exceptionVec_14=0x%0h",this.io_writeback_23_bits_exceptionVec_14,rhs_.io_writeback_23_bits_exceptionVec_14),UVM_NONE)
        end

        if(this.io_writeback_23_bits_exceptionVec_15!=rhs_.io_writeback_23_bits_exceptionVec_15) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_exceptionVec_15=0x%0h while the rhs_.io_writeback_23_bits_exceptionVec_15=0x%0h",this.io_writeback_23_bits_exceptionVec_15,rhs_.io_writeback_23_bits_exceptionVec_15),UVM_NONE)
        end

        if(this.io_writeback_23_bits_exceptionVec_16!=rhs_.io_writeback_23_bits_exceptionVec_16) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_exceptionVec_16=0x%0h while the rhs_.io_writeback_23_bits_exceptionVec_16=0x%0h",this.io_writeback_23_bits_exceptionVec_16,rhs_.io_writeback_23_bits_exceptionVec_16),UVM_NONE)
        end

        if(this.io_writeback_23_bits_exceptionVec_17!=rhs_.io_writeback_23_bits_exceptionVec_17) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_exceptionVec_17=0x%0h while the rhs_.io_writeback_23_bits_exceptionVec_17=0x%0h",this.io_writeback_23_bits_exceptionVec_17,rhs_.io_writeback_23_bits_exceptionVec_17),UVM_NONE)
        end

        if(this.io_writeback_23_bits_exceptionVec_18!=rhs_.io_writeback_23_bits_exceptionVec_18) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_exceptionVec_18=0x%0h while the rhs_.io_writeback_23_bits_exceptionVec_18=0x%0h",this.io_writeback_23_bits_exceptionVec_18,rhs_.io_writeback_23_bits_exceptionVec_18),UVM_NONE)
        end

        if(this.io_writeback_23_bits_exceptionVec_19!=rhs_.io_writeback_23_bits_exceptionVec_19) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_exceptionVec_19=0x%0h while the rhs_.io_writeback_23_bits_exceptionVec_19=0x%0h",this.io_writeback_23_bits_exceptionVec_19,rhs_.io_writeback_23_bits_exceptionVec_19),UVM_NONE)
        end

        if(this.io_writeback_23_bits_exceptionVec_20!=rhs_.io_writeback_23_bits_exceptionVec_20) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_exceptionVec_20=0x%0h while the rhs_.io_writeback_23_bits_exceptionVec_20=0x%0h",this.io_writeback_23_bits_exceptionVec_20,rhs_.io_writeback_23_bits_exceptionVec_20),UVM_NONE)
        end

        if(this.io_writeback_23_bits_exceptionVec_21!=rhs_.io_writeback_23_bits_exceptionVec_21) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_exceptionVec_21=0x%0h while the rhs_.io_writeback_23_bits_exceptionVec_21=0x%0h",this.io_writeback_23_bits_exceptionVec_21,rhs_.io_writeback_23_bits_exceptionVec_21),UVM_NONE)
        end

        if(this.io_writeback_23_bits_exceptionVec_22!=rhs_.io_writeback_23_bits_exceptionVec_22) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_exceptionVec_22=0x%0h while the rhs_.io_writeback_23_bits_exceptionVec_22=0x%0h",this.io_writeback_23_bits_exceptionVec_22,rhs_.io_writeback_23_bits_exceptionVec_22),UVM_NONE)
        end

        if(this.io_writeback_23_bits_exceptionVec_23!=rhs_.io_writeback_23_bits_exceptionVec_23) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_exceptionVec_23=0x%0h while the rhs_.io_writeback_23_bits_exceptionVec_23=0x%0h",this.io_writeback_23_bits_exceptionVec_23,rhs_.io_writeback_23_bits_exceptionVec_23),UVM_NONE)
        end

        if(this.io_writeback_23_bits_flushPipe!=rhs_.io_writeback_23_bits_flushPipe) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_flushPipe=0x%0h while the rhs_.io_writeback_23_bits_flushPipe=0x%0h",this.io_writeback_23_bits_flushPipe,rhs_.io_writeback_23_bits_flushPipe),UVM_NONE)
        end

        if(this.io_writeback_23_bits_replay!=rhs_.io_writeback_23_bits_replay) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_replay=0x%0h while the rhs_.io_writeback_23_bits_replay=0x%0h",this.io_writeback_23_bits_replay,rhs_.io_writeback_23_bits_replay),UVM_NONE)
        end

        if(this.io_writeback_23_bits_trigger!=rhs_.io_writeback_23_bits_trigger) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_trigger=0x%0h while the rhs_.io_writeback_23_bits_trigger=0x%0h",this.io_writeback_23_bits_trigger,rhs_.io_writeback_23_bits_trigger),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_vill!=rhs_.io_writeback_23_bits_vls_vpu_vill) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_vill=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_vill=0x%0h",this.io_writeback_23_bits_vls_vpu_vill,rhs_.io_writeback_23_bits_vls_vpu_vill),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_vma!=rhs_.io_writeback_23_bits_vls_vpu_vma) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_vma=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_vma=0x%0h",this.io_writeback_23_bits_vls_vpu_vma,rhs_.io_writeback_23_bits_vls_vpu_vma),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_vta!=rhs_.io_writeback_23_bits_vls_vpu_vta) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_vta=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_vta=0x%0h",this.io_writeback_23_bits_vls_vpu_vta,rhs_.io_writeback_23_bits_vls_vpu_vta),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_vsew!=rhs_.io_writeback_23_bits_vls_vpu_vsew) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_vsew=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_vsew=0x%0h",this.io_writeback_23_bits_vls_vpu_vsew,rhs_.io_writeback_23_bits_vls_vpu_vsew),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_vlmul!=rhs_.io_writeback_23_bits_vls_vpu_vlmul) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_vlmul=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_vlmul=0x%0h",this.io_writeback_23_bits_vls_vpu_vlmul,rhs_.io_writeback_23_bits_vls_vpu_vlmul),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_specVill!=rhs_.io_writeback_23_bits_vls_vpu_specVill) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_specVill=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_specVill=0x%0h",this.io_writeback_23_bits_vls_vpu_specVill,rhs_.io_writeback_23_bits_vls_vpu_specVill),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_specVma!=rhs_.io_writeback_23_bits_vls_vpu_specVma) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_specVma=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_specVma=0x%0h",this.io_writeback_23_bits_vls_vpu_specVma,rhs_.io_writeback_23_bits_vls_vpu_specVma),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_specVta!=rhs_.io_writeback_23_bits_vls_vpu_specVta) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_specVta=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_specVta=0x%0h",this.io_writeback_23_bits_vls_vpu_specVta,rhs_.io_writeback_23_bits_vls_vpu_specVta),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_specVsew!=rhs_.io_writeback_23_bits_vls_vpu_specVsew) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_specVsew=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_specVsew=0x%0h",this.io_writeback_23_bits_vls_vpu_specVsew,rhs_.io_writeback_23_bits_vls_vpu_specVsew),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_specVlmul!=rhs_.io_writeback_23_bits_vls_vpu_specVlmul) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_specVlmul=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_specVlmul=0x%0h",this.io_writeback_23_bits_vls_vpu_specVlmul,rhs_.io_writeback_23_bits_vls_vpu_specVlmul),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_vm!=rhs_.io_writeback_23_bits_vls_vpu_vm) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_vm=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_vm=0x%0h",this.io_writeback_23_bits_vls_vpu_vm,rhs_.io_writeback_23_bits_vls_vpu_vm),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_vstart!=rhs_.io_writeback_23_bits_vls_vpu_vstart) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_vstart=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_vstart=0x%0h",this.io_writeback_23_bits_vls_vpu_vstart,rhs_.io_writeback_23_bits_vls_vpu_vstart),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_frm!=rhs_.io_writeback_23_bits_vls_vpu_frm) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_frm=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_frm=0x%0h",this.io_writeback_23_bits_vls_vpu_frm,rhs_.io_writeback_23_bits_vls_vpu_frm),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst!=rhs_.io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst=0x%0h",this.io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst,rhs_.io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_fpu_isFP32Instr!=rhs_.io_writeback_23_bits_vls_vpu_fpu_isFP32Instr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_fpu_isFP32Instr=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_fpu_isFP32Instr=0x%0h",this.io_writeback_23_bits_vls_vpu_fpu_isFP32Instr,rhs_.io_writeback_23_bits_vls_vpu_fpu_isFP32Instr),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_fpu_isFP64Instr!=rhs_.io_writeback_23_bits_vls_vpu_fpu_isFP64Instr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_fpu_isFP64Instr=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_fpu_isFP64Instr=0x%0h",this.io_writeback_23_bits_vls_vpu_fpu_isFP64Instr,rhs_.io_writeback_23_bits_vls_vpu_fpu_isFP64Instr),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_fpu_isReduction!=rhs_.io_writeback_23_bits_vls_vpu_fpu_isReduction) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_fpu_isReduction=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_fpu_isReduction=0x%0h",this.io_writeback_23_bits_vls_vpu_fpu_isReduction,rhs_.io_writeback_23_bits_vls_vpu_fpu_isReduction),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2!=rhs_.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2=0x%0h",this.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2,rhs_.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4!=rhs_.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4=0x%0h",this.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4,rhs_.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8!=rhs_.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8=0x%0h",this.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8,rhs_.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_vxrm!=rhs_.io_writeback_23_bits_vls_vpu_vxrm) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_vxrm=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_vxrm=0x%0h",this.io_writeback_23_bits_vls_vpu_vxrm,rhs_.io_writeback_23_bits_vls_vpu_vxrm),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_vuopIdx!=rhs_.io_writeback_23_bits_vls_vpu_vuopIdx) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_vuopIdx=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_vuopIdx=0x%0h",this.io_writeback_23_bits_vls_vpu_vuopIdx,rhs_.io_writeback_23_bits_vls_vpu_vuopIdx),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_lastUop!=rhs_.io_writeback_23_bits_vls_vpu_lastUop) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_lastUop=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_lastUop=0x%0h",this.io_writeback_23_bits_vls_vpu_lastUop,rhs_.io_writeback_23_bits_vls_vpu_lastUop),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_vmask!=rhs_.io_writeback_23_bits_vls_vpu_vmask) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_vmask=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_vmask=0x%0h",this.io_writeback_23_bits_vls_vpu_vmask,rhs_.io_writeback_23_bits_vls_vpu_vmask),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_vl!=rhs_.io_writeback_23_bits_vls_vpu_vl) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_vl=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_vl=0x%0h",this.io_writeback_23_bits_vls_vpu_vl,rhs_.io_writeback_23_bits_vls_vpu_vl),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_nf!=rhs_.io_writeback_23_bits_vls_vpu_nf) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_nf=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_nf=0x%0h",this.io_writeback_23_bits_vls_vpu_nf,rhs_.io_writeback_23_bits_vls_vpu_nf),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_veew!=rhs_.io_writeback_23_bits_vls_vpu_veew) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_veew=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_veew=0x%0h",this.io_writeback_23_bits_vls_vpu_veew,rhs_.io_writeback_23_bits_vls_vpu_veew),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_isReverse!=rhs_.io_writeback_23_bits_vls_vpu_isReverse) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_isReverse=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_isReverse=0x%0h",this.io_writeback_23_bits_vls_vpu_isReverse,rhs_.io_writeback_23_bits_vls_vpu_isReverse),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_isExt!=rhs_.io_writeback_23_bits_vls_vpu_isExt) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_isExt=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_isExt=0x%0h",this.io_writeback_23_bits_vls_vpu_isExt,rhs_.io_writeback_23_bits_vls_vpu_isExt),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_isNarrow!=rhs_.io_writeback_23_bits_vls_vpu_isNarrow) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_isNarrow=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_isNarrow=0x%0h",this.io_writeback_23_bits_vls_vpu_isNarrow,rhs_.io_writeback_23_bits_vls_vpu_isNarrow),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_isDstMask!=rhs_.io_writeback_23_bits_vls_vpu_isDstMask) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_isDstMask=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_isDstMask=0x%0h",this.io_writeback_23_bits_vls_vpu_isDstMask,rhs_.io_writeback_23_bits_vls_vpu_isDstMask),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_isOpMask!=rhs_.io_writeback_23_bits_vls_vpu_isOpMask) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_isOpMask=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_isOpMask=0x%0h",this.io_writeback_23_bits_vls_vpu_isOpMask,rhs_.io_writeback_23_bits_vls_vpu_isOpMask),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_isMove!=rhs_.io_writeback_23_bits_vls_vpu_isMove) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_isMove=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_isMove=0x%0h",this.io_writeback_23_bits_vls_vpu_isMove,rhs_.io_writeback_23_bits_vls_vpu_isMove),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_isDependOldVd!=rhs_.io_writeback_23_bits_vls_vpu_isDependOldVd) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_isDependOldVd=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_isDependOldVd=0x%0h",this.io_writeback_23_bits_vls_vpu_isDependOldVd,rhs_.io_writeback_23_bits_vls_vpu_isDependOldVd),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_isWritePartVd!=rhs_.io_writeback_23_bits_vls_vpu_isWritePartVd) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_isWritePartVd=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_isWritePartVd=0x%0h",this.io_writeback_23_bits_vls_vpu_isWritePartVd,rhs_.io_writeback_23_bits_vls_vpu_isWritePartVd),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vpu_isVleff!=rhs_.io_writeback_23_bits_vls_vpu_isVleff) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vpu_isVleff=0x%0h while the rhs_.io_writeback_23_bits_vls_vpu_isVleff=0x%0h",this.io_writeback_23_bits_vls_vpu_isVleff,rhs_.io_writeback_23_bits_vls_vpu_isVleff),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_oldVdPsrc!=rhs_.io_writeback_23_bits_vls_oldVdPsrc) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_oldVdPsrc=0x%0h while the rhs_.io_writeback_23_bits_vls_oldVdPsrc=0x%0h",this.io_writeback_23_bits_vls_oldVdPsrc,rhs_.io_writeback_23_bits_vls_oldVdPsrc),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vdIdx!=rhs_.io_writeback_23_bits_vls_vdIdx) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vdIdx=0x%0h while the rhs_.io_writeback_23_bits_vls_vdIdx=0x%0h",this.io_writeback_23_bits_vls_vdIdx,rhs_.io_writeback_23_bits_vls_vdIdx),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_vdIdxInField!=rhs_.io_writeback_23_bits_vls_vdIdxInField) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_vdIdxInField=0x%0h while the rhs_.io_writeback_23_bits_vls_vdIdxInField=0x%0h",this.io_writeback_23_bits_vls_vdIdxInField,rhs_.io_writeback_23_bits_vls_vdIdxInField),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_isIndexed!=rhs_.io_writeback_23_bits_vls_isIndexed) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_isIndexed=0x%0h while the rhs_.io_writeback_23_bits_vls_isIndexed=0x%0h",this.io_writeback_23_bits_vls_isIndexed,rhs_.io_writeback_23_bits_vls_isIndexed),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_isMasked!=rhs_.io_writeback_23_bits_vls_isMasked) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_isMasked=0x%0h while the rhs_.io_writeback_23_bits_vls_isMasked=0x%0h",this.io_writeback_23_bits_vls_isMasked,rhs_.io_writeback_23_bits_vls_isMasked),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_isStrided!=rhs_.io_writeback_23_bits_vls_isStrided) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_isStrided=0x%0h while the rhs_.io_writeback_23_bits_vls_isStrided=0x%0h",this.io_writeback_23_bits_vls_isStrided,rhs_.io_writeback_23_bits_vls_isStrided),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_isWhole!=rhs_.io_writeback_23_bits_vls_isWhole) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_isWhole=0x%0h while the rhs_.io_writeback_23_bits_vls_isWhole=0x%0h",this.io_writeback_23_bits_vls_isWhole,rhs_.io_writeback_23_bits_vls_isWhole),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_isVecLoad!=rhs_.io_writeback_23_bits_vls_isVecLoad) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_isVecLoad=0x%0h while the rhs_.io_writeback_23_bits_vls_isVecLoad=0x%0h",this.io_writeback_23_bits_vls_isVecLoad,rhs_.io_writeback_23_bits_vls_isVecLoad),UVM_NONE)
        end

        if(this.io_writeback_23_bits_vls_isVlm!=rhs_.io_writeback_23_bits_vls_isVlm) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_vls_isVlm=0x%0h while the rhs_.io_writeback_23_bits_vls_isVlm=0x%0h",this.io_writeback_23_bits_vls_isVlm,rhs_.io_writeback_23_bits_vls_isVlm),UVM_NONE)
        end

        if(this.io_writeback_23_bits_debug_isMMIO!=rhs_.io_writeback_23_bits_debug_isMMIO) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_debug_isMMIO=0x%0h while the rhs_.io_writeback_23_bits_debug_isMMIO=0x%0h",this.io_writeback_23_bits_debug_isMMIO,rhs_.io_writeback_23_bits_debug_isMMIO),UVM_NONE)
        end

        if(this.io_writeback_23_bits_debug_isNCIO!=rhs_.io_writeback_23_bits_debug_isNCIO) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_debug_isNCIO=0x%0h while the rhs_.io_writeback_23_bits_debug_isNCIO=0x%0h",this.io_writeback_23_bits_debug_isNCIO,rhs_.io_writeback_23_bits_debug_isNCIO),UVM_NONE)
        end

        if(this.io_writeback_23_bits_debug_isPerfCnt!=rhs_.io_writeback_23_bits_debug_isPerfCnt) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_debug_isPerfCnt=0x%0h while the rhs_.io_writeback_23_bits_debug_isPerfCnt=0x%0h",this.io_writeback_23_bits_debug_isPerfCnt,rhs_.io_writeback_23_bits_debug_isPerfCnt),UVM_NONE)
        end

        if(this.io_writeback_23_bits_debug_paddr!=rhs_.io_writeback_23_bits_debug_paddr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_debug_paddr=0x%0h while the rhs_.io_writeback_23_bits_debug_paddr=0x%0h",this.io_writeback_23_bits_debug_paddr,rhs_.io_writeback_23_bits_debug_paddr),UVM_NONE)
        end

        if(this.io_writeback_23_bits_debug_vaddr!=rhs_.io_writeback_23_bits_debug_vaddr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_debug_vaddr=0x%0h while the rhs_.io_writeback_23_bits_debug_vaddr=0x%0h",this.io_writeback_23_bits_debug_vaddr,rhs_.io_writeback_23_bits_debug_vaddr),UVM_NONE)
        end

        if(this.io_writeback_23_bits_debugInfo_eliminatedMove!=rhs_.io_writeback_23_bits_debugInfo_eliminatedMove) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_debugInfo_eliminatedMove=0x%0h while the rhs_.io_writeback_23_bits_debugInfo_eliminatedMove=0x%0h",this.io_writeback_23_bits_debugInfo_eliminatedMove,rhs_.io_writeback_23_bits_debugInfo_eliminatedMove),UVM_NONE)
        end

        if(this.io_writeback_23_bits_debugInfo_renameTime!=rhs_.io_writeback_23_bits_debugInfo_renameTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_debugInfo_renameTime=0x%0h while the rhs_.io_writeback_23_bits_debugInfo_renameTime=0x%0h",this.io_writeback_23_bits_debugInfo_renameTime,rhs_.io_writeback_23_bits_debugInfo_renameTime),UVM_NONE)
        end

        if(this.io_writeback_23_bits_debugInfo_dispatchTime!=rhs_.io_writeback_23_bits_debugInfo_dispatchTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_debugInfo_dispatchTime=0x%0h while the rhs_.io_writeback_23_bits_debugInfo_dispatchTime=0x%0h",this.io_writeback_23_bits_debugInfo_dispatchTime,rhs_.io_writeback_23_bits_debugInfo_dispatchTime),UVM_NONE)
        end

        if(this.io_writeback_23_bits_debugInfo_enqRsTime!=rhs_.io_writeback_23_bits_debugInfo_enqRsTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_debugInfo_enqRsTime=0x%0h while the rhs_.io_writeback_23_bits_debugInfo_enqRsTime=0x%0h",this.io_writeback_23_bits_debugInfo_enqRsTime,rhs_.io_writeback_23_bits_debugInfo_enqRsTime),UVM_NONE)
        end

        if(this.io_writeback_23_bits_debugInfo_selectTime!=rhs_.io_writeback_23_bits_debugInfo_selectTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_debugInfo_selectTime=0x%0h while the rhs_.io_writeback_23_bits_debugInfo_selectTime=0x%0h",this.io_writeback_23_bits_debugInfo_selectTime,rhs_.io_writeback_23_bits_debugInfo_selectTime),UVM_NONE)
        end

        if(this.io_writeback_23_bits_debugInfo_issueTime!=rhs_.io_writeback_23_bits_debugInfo_issueTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_debugInfo_issueTime=0x%0h while the rhs_.io_writeback_23_bits_debugInfo_issueTime=0x%0h",this.io_writeback_23_bits_debugInfo_issueTime,rhs_.io_writeback_23_bits_debugInfo_issueTime),UVM_NONE)
        end

        if(this.io_writeback_23_bits_debugInfo_writebackTime!=rhs_.io_writeback_23_bits_debugInfo_writebackTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_debugInfo_writebackTime=0x%0h while the rhs_.io_writeback_23_bits_debugInfo_writebackTime=0x%0h",this.io_writeback_23_bits_debugInfo_writebackTime,rhs_.io_writeback_23_bits_debugInfo_writebackTime),UVM_NONE)
        end

        if(this.io_writeback_23_bits_debugInfo_runahead_checkpoint_id!=rhs_.io_writeback_23_bits_debugInfo_runahead_checkpoint_id) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_debugInfo_runahead_checkpoint_id=0x%0h while the rhs_.io_writeback_23_bits_debugInfo_runahead_checkpoint_id=0x%0h",this.io_writeback_23_bits_debugInfo_runahead_checkpoint_id,rhs_.io_writeback_23_bits_debugInfo_runahead_checkpoint_id),UVM_NONE)
        end

        if(this.io_writeback_23_bits_debugInfo_tlbFirstReqTime!=rhs_.io_writeback_23_bits_debugInfo_tlbFirstReqTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_debugInfo_tlbFirstReqTime=0x%0h while the rhs_.io_writeback_23_bits_debugInfo_tlbFirstReqTime=0x%0h",this.io_writeback_23_bits_debugInfo_tlbFirstReqTime,rhs_.io_writeback_23_bits_debugInfo_tlbFirstReqTime),UVM_NONE)
        end

        if(this.io_writeback_23_bits_debugInfo_tlbRespTime!=rhs_.io_writeback_23_bits_debugInfo_tlbRespTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_debugInfo_tlbRespTime=0x%0h while the rhs_.io_writeback_23_bits_debugInfo_tlbRespTime=0x%0h",this.io_writeback_23_bits_debugInfo_tlbRespTime,rhs_.io_writeback_23_bits_debugInfo_tlbRespTime),UVM_NONE)
        end

        if(this.io_writeback_23_bits_debug_seqNum!=rhs_.io_writeback_23_bits_debug_seqNum) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_23_bits_debug_seqNum=0x%0h while the rhs_.io_writeback_23_bits_debug_seqNum=0x%0h",this.io_writeback_23_bits_debug_seqNum,rhs_.io_writeback_23_bits_debug_seqNum),UVM_NONE)
        end

        if(this.io_writeback_22_valid!=rhs_.io_writeback_22_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_valid=0x%0h while the rhs_.io_writeback_22_valid=0x%0h",this.io_writeback_22_valid,rhs_.io_writeback_22_valid),UVM_NONE)
        end

        if(this.io_writeback_22_bits_data_0!=rhs_.io_writeback_22_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_data_0=0x%0h while the rhs_.io_writeback_22_bits_data_0=0x%0h",this.io_writeback_22_bits_data_0,rhs_.io_writeback_22_bits_data_0),UVM_NONE)
        end

        if(this.io_writeback_22_bits_pdest!=rhs_.io_writeback_22_bits_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_pdest=0x%0h while the rhs_.io_writeback_22_bits_pdest=0x%0h",this.io_writeback_22_bits_pdest,rhs_.io_writeback_22_bits_pdest),UVM_NONE)
        end

        if(this.io_writeback_22_bits_robIdx_flag!=rhs_.io_writeback_22_bits_robIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_robIdx_flag=0x%0h while the rhs_.io_writeback_22_bits_robIdx_flag=0x%0h",this.io_writeback_22_bits_robIdx_flag,rhs_.io_writeback_22_bits_robIdx_flag),UVM_NONE)
        end

        if(this.io_writeback_22_bits_robIdx_value!=rhs_.io_writeback_22_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_robIdx_value=0x%0h while the rhs_.io_writeback_22_bits_robIdx_value=0x%0h",this.io_writeback_22_bits_robIdx_value,rhs_.io_writeback_22_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_writeback_22_bits_intWen!=rhs_.io_writeback_22_bits_intWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_intWen=0x%0h while the rhs_.io_writeback_22_bits_intWen=0x%0h",this.io_writeback_22_bits_intWen,rhs_.io_writeback_22_bits_intWen),UVM_NONE)
        end

        if(this.io_writeback_22_bits_fpWen!=rhs_.io_writeback_22_bits_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_fpWen=0x%0h while the rhs_.io_writeback_22_bits_fpWen=0x%0h",this.io_writeback_22_bits_fpWen,rhs_.io_writeback_22_bits_fpWen),UVM_NONE)
        end

        if(this.io_writeback_22_bits_exceptionVec_0!=rhs_.io_writeback_22_bits_exceptionVec_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_exceptionVec_0=0x%0h while the rhs_.io_writeback_22_bits_exceptionVec_0=0x%0h",this.io_writeback_22_bits_exceptionVec_0,rhs_.io_writeback_22_bits_exceptionVec_0),UVM_NONE)
        end

        if(this.io_writeback_22_bits_exceptionVec_1!=rhs_.io_writeback_22_bits_exceptionVec_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_exceptionVec_1=0x%0h while the rhs_.io_writeback_22_bits_exceptionVec_1=0x%0h",this.io_writeback_22_bits_exceptionVec_1,rhs_.io_writeback_22_bits_exceptionVec_1),UVM_NONE)
        end

        if(this.io_writeback_22_bits_exceptionVec_2!=rhs_.io_writeback_22_bits_exceptionVec_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_exceptionVec_2=0x%0h while the rhs_.io_writeback_22_bits_exceptionVec_2=0x%0h",this.io_writeback_22_bits_exceptionVec_2,rhs_.io_writeback_22_bits_exceptionVec_2),UVM_NONE)
        end

        if(this.io_writeback_22_bits_exceptionVec_3!=rhs_.io_writeback_22_bits_exceptionVec_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_exceptionVec_3=0x%0h while the rhs_.io_writeback_22_bits_exceptionVec_3=0x%0h",this.io_writeback_22_bits_exceptionVec_3,rhs_.io_writeback_22_bits_exceptionVec_3),UVM_NONE)
        end

        if(this.io_writeback_22_bits_exceptionVec_4!=rhs_.io_writeback_22_bits_exceptionVec_4) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_exceptionVec_4=0x%0h while the rhs_.io_writeback_22_bits_exceptionVec_4=0x%0h",this.io_writeback_22_bits_exceptionVec_4,rhs_.io_writeback_22_bits_exceptionVec_4),UVM_NONE)
        end

        if(this.io_writeback_22_bits_exceptionVec_5!=rhs_.io_writeback_22_bits_exceptionVec_5) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_exceptionVec_5=0x%0h while the rhs_.io_writeback_22_bits_exceptionVec_5=0x%0h",this.io_writeback_22_bits_exceptionVec_5,rhs_.io_writeback_22_bits_exceptionVec_5),UVM_NONE)
        end

        if(this.io_writeback_22_bits_exceptionVec_6!=rhs_.io_writeback_22_bits_exceptionVec_6) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_exceptionVec_6=0x%0h while the rhs_.io_writeback_22_bits_exceptionVec_6=0x%0h",this.io_writeback_22_bits_exceptionVec_6,rhs_.io_writeback_22_bits_exceptionVec_6),UVM_NONE)
        end

        if(this.io_writeback_22_bits_exceptionVec_7!=rhs_.io_writeback_22_bits_exceptionVec_7) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_exceptionVec_7=0x%0h while the rhs_.io_writeback_22_bits_exceptionVec_7=0x%0h",this.io_writeback_22_bits_exceptionVec_7,rhs_.io_writeback_22_bits_exceptionVec_7),UVM_NONE)
        end

        if(this.io_writeback_22_bits_exceptionVec_8!=rhs_.io_writeback_22_bits_exceptionVec_8) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_exceptionVec_8=0x%0h while the rhs_.io_writeback_22_bits_exceptionVec_8=0x%0h",this.io_writeback_22_bits_exceptionVec_8,rhs_.io_writeback_22_bits_exceptionVec_8),UVM_NONE)
        end

        if(this.io_writeback_22_bits_exceptionVec_9!=rhs_.io_writeback_22_bits_exceptionVec_9) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_exceptionVec_9=0x%0h while the rhs_.io_writeback_22_bits_exceptionVec_9=0x%0h",this.io_writeback_22_bits_exceptionVec_9,rhs_.io_writeback_22_bits_exceptionVec_9),UVM_NONE)
        end

        if(this.io_writeback_22_bits_exceptionVec_10!=rhs_.io_writeback_22_bits_exceptionVec_10) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_exceptionVec_10=0x%0h while the rhs_.io_writeback_22_bits_exceptionVec_10=0x%0h",this.io_writeback_22_bits_exceptionVec_10,rhs_.io_writeback_22_bits_exceptionVec_10),UVM_NONE)
        end

        if(this.io_writeback_22_bits_exceptionVec_11!=rhs_.io_writeback_22_bits_exceptionVec_11) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_exceptionVec_11=0x%0h while the rhs_.io_writeback_22_bits_exceptionVec_11=0x%0h",this.io_writeback_22_bits_exceptionVec_11,rhs_.io_writeback_22_bits_exceptionVec_11),UVM_NONE)
        end

        if(this.io_writeback_22_bits_exceptionVec_12!=rhs_.io_writeback_22_bits_exceptionVec_12) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_exceptionVec_12=0x%0h while the rhs_.io_writeback_22_bits_exceptionVec_12=0x%0h",this.io_writeback_22_bits_exceptionVec_12,rhs_.io_writeback_22_bits_exceptionVec_12),UVM_NONE)
        end

        if(this.io_writeback_22_bits_exceptionVec_13!=rhs_.io_writeback_22_bits_exceptionVec_13) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_exceptionVec_13=0x%0h while the rhs_.io_writeback_22_bits_exceptionVec_13=0x%0h",this.io_writeback_22_bits_exceptionVec_13,rhs_.io_writeback_22_bits_exceptionVec_13),UVM_NONE)
        end

        if(this.io_writeback_22_bits_exceptionVec_14!=rhs_.io_writeback_22_bits_exceptionVec_14) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_exceptionVec_14=0x%0h while the rhs_.io_writeback_22_bits_exceptionVec_14=0x%0h",this.io_writeback_22_bits_exceptionVec_14,rhs_.io_writeback_22_bits_exceptionVec_14),UVM_NONE)
        end

        if(this.io_writeback_22_bits_exceptionVec_15!=rhs_.io_writeback_22_bits_exceptionVec_15) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_exceptionVec_15=0x%0h while the rhs_.io_writeback_22_bits_exceptionVec_15=0x%0h",this.io_writeback_22_bits_exceptionVec_15,rhs_.io_writeback_22_bits_exceptionVec_15),UVM_NONE)
        end

        if(this.io_writeback_22_bits_exceptionVec_16!=rhs_.io_writeback_22_bits_exceptionVec_16) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_exceptionVec_16=0x%0h while the rhs_.io_writeback_22_bits_exceptionVec_16=0x%0h",this.io_writeback_22_bits_exceptionVec_16,rhs_.io_writeback_22_bits_exceptionVec_16),UVM_NONE)
        end

        if(this.io_writeback_22_bits_exceptionVec_17!=rhs_.io_writeback_22_bits_exceptionVec_17) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_exceptionVec_17=0x%0h while the rhs_.io_writeback_22_bits_exceptionVec_17=0x%0h",this.io_writeback_22_bits_exceptionVec_17,rhs_.io_writeback_22_bits_exceptionVec_17),UVM_NONE)
        end

        if(this.io_writeback_22_bits_exceptionVec_18!=rhs_.io_writeback_22_bits_exceptionVec_18) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_exceptionVec_18=0x%0h while the rhs_.io_writeback_22_bits_exceptionVec_18=0x%0h",this.io_writeback_22_bits_exceptionVec_18,rhs_.io_writeback_22_bits_exceptionVec_18),UVM_NONE)
        end

        if(this.io_writeback_22_bits_exceptionVec_19!=rhs_.io_writeback_22_bits_exceptionVec_19) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_exceptionVec_19=0x%0h while the rhs_.io_writeback_22_bits_exceptionVec_19=0x%0h",this.io_writeback_22_bits_exceptionVec_19,rhs_.io_writeback_22_bits_exceptionVec_19),UVM_NONE)
        end

        if(this.io_writeback_22_bits_exceptionVec_20!=rhs_.io_writeback_22_bits_exceptionVec_20) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_exceptionVec_20=0x%0h while the rhs_.io_writeback_22_bits_exceptionVec_20=0x%0h",this.io_writeback_22_bits_exceptionVec_20,rhs_.io_writeback_22_bits_exceptionVec_20),UVM_NONE)
        end

        if(this.io_writeback_22_bits_exceptionVec_21!=rhs_.io_writeback_22_bits_exceptionVec_21) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_exceptionVec_21=0x%0h while the rhs_.io_writeback_22_bits_exceptionVec_21=0x%0h",this.io_writeback_22_bits_exceptionVec_21,rhs_.io_writeback_22_bits_exceptionVec_21),UVM_NONE)
        end

        if(this.io_writeback_22_bits_exceptionVec_22!=rhs_.io_writeback_22_bits_exceptionVec_22) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_exceptionVec_22=0x%0h while the rhs_.io_writeback_22_bits_exceptionVec_22=0x%0h",this.io_writeback_22_bits_exceptionVec_22,rhs_.io_writeback_22_bits_exceptionVec_22),UVM_NONE)
        end

        if(this.io_writeback_22_bits_exceptionVec_23!=rhs_.io_writeback_22_bits_exceptionVec_23) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_exceptionVec_23=0x%0h while the rhs_.io_writeback_22_bits_exceptionVec_23=0x%0h",this.io_writeback_22_bits_exceptionVec_23,rhs_.io_writeback_22_bits_exceptionVec_23),UVM_NONE)
        end

        if(this.io_writeback_22_bits_flushPipe!=rhs_.io_writeback_22_bits_flushPipe) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_flushPipe=0x%0h while the rhs_.io_writeback_22_bits_flushPipe=0x%0h",this.io_writeback_22_bits_flushPipe,rhs_.io_writeback_22_bits_flushPipe),UVM_NONE)
        end

        if(this.io_writeback_22_bits_replay!=rhs_.io_writeback_22_bits_replay) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_replay=0x%0h while the rhs_.io_writeback_22_bits_replay=0x%0h",this.io_writeback_22_bits_replay,rhs_.io_writeback_22_bits_replay),UVM_NONE)
        end

        if(this.io_writeback_22_bits_lqIdx_flag!=rhs_.io_writeback_22_bits_lqIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_lqIdx_flag=0x%0h while the rhs_.io_writeback_22_bits_lqIdx_flag=0x%0h",this.io_writeback_22_bits_lqIdx_flag,rhs_.io_writeback_22_bits_lqIdx_flag),UVM_NONE)
        end

        if(this.io_writeback_22_bits_lqIdx_value!=rhs_.io_writeback_22_bits_lqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_lqIdx_value=0x%0h while the rhs_.io_writeback_22_bits_lqIdx_value=0x%0h",this.io_writeback_22_bits_lqIdx_value,rhs_.io_writeback_22_bits_lqIdx_value),UVM_NONE)
        end

        if(this.io_writeback_22_bits_trigger!=rhs_.io_writeback_22_bits_trigger) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_trigger=0x%0h while the rhs_.io_writeback_22_bits_trigger=0x%0h",this.io_writeback_22_bits_trigger,rhs_.io_writeback_22_bits_trigger),UVM_NONE)
        end

        if(this.io_writeback_22_bits_predecodeInfo_valid!=rhs_.io_writeback_22_bits_predecodeInfo_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_predecodeInfo_valid=0x%0h while the rhs_.io_writeback_22_bits_predecodeInfo_valid=0x%0h",this.io_writeback_22_bits_predecodeInfo_valid,rhs_.io_writeback_22_bits_predecodeInfo_valid),UVM_NONE)
        end

        if(this.io_writeback_22_bits_predecodeInfo_isRVC!=rhs_.io_writeback_22_bits_predecodeInfo_isRVC) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_predecodeInfo_isRVC=0x%0h while the rhs_.io_writeback_22_bits_predecodeInfo_isRVC=0x%0h",this.io_writeback_22_bits_predecodeInfo_isRVC,rhs_.io_writeback_22_bits_predecodeInfo_isRVC),UVM_NONE)
        end

        if(this.io_writeback_22_bits_predecodeInfo_brType!=rhs_.io_writeback_22_bits_predecodeInfo_brType) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_predecodeInfo_brType=0x%0h while the rhs_.io_writeback_22_bits_predecodeInfo_brType=0x%0h",this.io_writeback_22_bits_predecodeInfo_brType,rhs_.io_writeback_22_bits_predecodeInfo_brType),UVM_NONE)
        end

        if(this.io_writeback_22_bits_predecodeInfo_isCall!=rhs_.io_writeback_22_bits_predecodeInfo_isCall) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_predecodeInfo_isCall=0x%0h while the rhs_.io_writeback_22_bits_predecodeInfo_isCall=0x%0h",this.io_writeback_22_bits_predecodeInfo_isCall,rhs_.io_writeback_22_bits_predecodeInfo_isCall),UVM_NONE)
        end

        if(this.io_writeback_22_bits_predecodeInfo_isRet!=rhs_.io_writeback_22_bits_predecodeInfo_isRet) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_predecodeInfo_isRet=0x%0h while the rhs_.io_writeback_22_bits_predecodeInfo_isRet=0x%0h",this.io_writeback_22_bits_predecodeInfo_isRet,rhs_.io_writeback_22_bits_predecodeInfo_isRet),UVM_NONE)
        end

        if(this.io_writeback_22_bits_debug_isMMIO!=rhs_.io_writeback_22_bits_debug_isMMIO) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_debug_isMMIO=0x%0h while the rhs_.io_writeback_22_bits_debug_isMMIO=0x%0h",this.io_writeback_22_bits_debug_isMMIO,rhs_.io_writeback_22_bits_debug_isMMIO),UVM_NONE)
        end

        if(this.io_writeback_22_bits_debug_isNCIO!=rhs_.io_writeback_22_bits_debug_isNCIO) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_debug_isNCIO=0x%0h while the rhs_.io_writeback_22_bits_debug_isNCIO=0x%0h",this.io_writeback_22_bits_debug_isNCIO,rhs_.io_writeback_22_bits_debug_isNCIO),UVM_NONE)
        end

        if(this.io_writeback_22_bits_debug_isPerfCnt!=rhs_.io_writeback_22_bits_debug_isPerfCnt) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_debug_isPerfCnt=0x%0h while the rhs_.io_writeback_22_bits_debug_isPerfCnt=0x%0h",this.io_writeback_22_bits_debug_isPerfCnt,rhs_.io_writeback_22_bits_debug_isPerfCnt),UVM_NONE)
        end

        if(this.io_writeback_22_bits_debug_paddr!=rhs_.io_writeback_22_bits_debug_paddr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_debug_paddr=0x%0h while the rhs_.io_writeback_22_bits_debug_paddr=0x%0h",this.io_writeback_22_bits_debug_paddr,rhs_.io_writeback_22_bits_debug_paddr),UVM_NONE)
        end

        if(this.io_writeback_22_bits_debug_vaddr!=rhs_.io_writeback_22_bits_debug_vaddr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_debug_vaddr=0x%0h while the rhs_.io_writeback_22_bits_debug_vaddr=0x%0h",this.io_writeback_22_bits_debug_vaddr,rhs_.io_writeback_22_bits_debug_vaddr),UVM_NONE)
        end

        if(this.io_writeback_22_bits_debugInfo_eliminatedMove!=rhs_.io_writeback_22_bits_debugInfo_eliminatedMove) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_debugInfo_eliminatedMove=0x%0h while the rhs_.io_writeback_22_bits_debugInfo_eliminatedMove=0x%0h",this.io_writeback_22_bits_debugInfo_eliminatedMove,rhs_.io_writeback_22_bits_debugInfo_eliminatedMove),UVM_NONE)
        end

        if(this.io_writeback_22_bits_debugInfo_renameTime!=rhs_.io_writeback_22_bits_debugInfo_renameTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_debugInfo_renameTime=0x%0h while the rhs_.io_writeback_22_bits_debugInfo_renameTime=0x%0h",this.io_writeback_22_bits_debugInfo_renameTime,rhs_.io_writeback_22_bits_debugInfo_renameTime),UVM_NONE)
        end

        if(this.io_writeback_22_bits_debugInfo_dispatchTime!=rhs_.io_writeback_22_bits_debugInfo_dispatchTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_debugInfo_dispatchTime=0x%0h while the rhs_.io_writeback_22_bits_debugInfo_dispatchTime=0x%0h",this.io_writeback_22_bits_debugInfo_dispatchTime,rhs_.io_writeback_22_bits_debugInfo_dispatchTime),UVM_NONE)
        end

        if(this.io_writeback_22_bits_debugInfo_enqRsTime!=rhs_.io_writeback_22_bits_debugInfo_enqRsTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_debugInfo_enqRsTime=0x%0h while the rhs_.io_writeback_22_bits_debugInfo_enqRsTime=0x%0h",this.io_writeback_22_bits_debugInfo_enqRsTime,rhs_.io_writeback_22_bits_debugInfo_enqRsTime),UVM_NONE)
        end

        if(this.io_writeback_22_bits_debugInfo_selectTime!=rhs_.io_writeback_22_bits_debugInfo_selectTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_debugInfo_selectTime=0x%0h while the rhs_.io_writeback_22_bits_debugInfo_selectTime=0x%0h",this.io_writeback_22_bits_debugInfo_selectTime,rhs_.io_writeback_22_bits_debugInfo_selectTime),UVM_NONE)
        end

        if(this.io_writeback_22_bits_debugInfo_issueTime!=rhs_.io_writeback_22_bits_debugInfo_issueTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_debugInfo_issueTime=0x%0h while the rhs_.io_writeback_22_bits_debugInfo_issueTime=0x%0h",this.io_writeback_22_bits_debugInfo_issueTime,rhs_.io_writeback_22_bits_debugInfo_issueTime),UVM_NONE)
        end

        if(this.io_writeback_22_bits_debugInfo_writebackTime!=rhs_.io_writeback_22_bits_debugInfo_writebackTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_debugInfo_writebackTime=0x%0h while the rhs_.io_writeback_22_bits_debugInfo_writebackTime=0x%0h",this.io_writeback_22_bits_debugInfo_writebackTime,rhs_.io_writeback_22_bits_debugInfo_writebackTime),UVM_NONE)
        end

        if(this.io_writeback_22_bits_debugInfo_runahead_checkpoint_id!=rhs_.io_writeback_22_bits_debugInfo_runahead_checkpoint_id) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_debugInfo_runahead_checkpoint_id=0x%0h while the rhs_.io_writeback_22_bits_debugInfo_runahead_checkpoint_id=0x%0h",this.io_writeback_22_bits_debugInfo_runahead_checkpoint_id,rhs_.io_writeback_22_bits_debugInfo_runahead_checkpoint_id),UVM_NONE)
        end

        if(this.io_writeback_22_bits_debugInfo_tlbFirstReqTime!=rhs_.io_writeback_22_bits_debugInfo_tlbFirstReqTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_debugInfo_tlbFirstReqTime=0x%0h while the rhs_.io_writeback_22_bits_debugInfo_tlbFirstReqTime=0x%0h",this.io_writeback_22_bits_debugInfo_tlbFirstReqTime,rhs_.io_writeback_22_bits_debugInfo_tlbFirstReqTime),UVM_NONE)
        end

        if(this.io_writeback_22_bits_debugInfo_tlbRespTime!=rhs_.io_writeback_22_bits_debugInfo_tlbRespTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_debugInfo_tlbRespTime=0x%0h while the rhs_.io_writeback_22_bits_debugInfo_tlbRespTime=0x%0h",this.io_writeback_22_bits_debugInfo_tlbRespTime,rhs_.io_writeback_22_bits_debugInfo_tlbRespTime),UVM_NONE)
        end

        if(this.io_writeback_22_bits_debug_seqNum!=rhs_.io_writeback_22_bits_debug_seqNum) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_22_bits_debug_seqNum=0x%0h while the rhs_.io_writeback_22_bits_debug_seqNum=0x%0h",this.io_writeback_22_bits_debug_seqNum,rhs_.io_writeback_22_bits_debug_seqNum),UVM_NONE)
        end

        if(this.io_writeback_21_valid!=rhs_.io_writeback_21_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_valid=0x%0h while the rhs_.io_writeback_21_valid=0x%0h",this.io_writeback_21_valid,rhs_.io_writeback_21_valid),UVM_NONE)
        end

        if(this.io_writeback_21_bits_data_0!=rhs_.io_writeback_21_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_data_0=0x%0h while the rhs_.io_writeback_21_bits_data_0=0x%0h",this.io_writeback_21_bits_data_0,rhs_.io_writeback_21_bits_data_0),UVM_NONE)
        end

        if(this.io_writeback_21_bits_pdest!=rhs_.io_writeback_21_bits_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_pdest=0x%0h while the rhs_.io_writeback_21_bits_pdest=0x%0h",this.io_writeback_21_bits_pdest,rhs_.io_writeback_21_bits_pdest),UVM_NONE)
        end

        if(this.io_writeback_21_bits_robIdx_flag!=rhs_.io_writeback_21_bits_robIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_robIdx_flag=0x%0h while the rhs_.io_writeback_21_bits_robIdx_flag=0x%0h",this.io_writeback_21_bits_robIdx_flag,rhs_.io_writeback_21_bits_robIdx_flag),UVM_NONE)
        end

        if(this.io_writeback_21_bits_robIdx_value!=rhs_.io_writeback_21_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_robIdx_value=0x%0h while the rhs_.io_writeback_21_bits_robIdx_value=0x%0h",this.io_writeback_21_bits_robIdx_value,rhs_.io_writeback_21_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_writeback_21_bits_intWen!=rhs_.io_writeback_21_bits_intWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_intWen=0x%0h while the rhs_.io_writeback_21_bits_intWen=0x%0h",this.io_writeback_21_bits_intWen,rhs_.io_writeback_21_bits_intWen),UVM_NONE)
        end

        if(this.io_writeback_21_bits_fpWen!=rhs_.io_writeback_21_bits_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_fpWen=0x%0h while the rhs_.io_writeback_21_bits_fpWen=0x%0h",this.io_writeback_21_bits_fpWen,rhs_.io_writeback_21_bits_fpWen),UVM_NONE)
        end

        if(this.io_writeback_21_bits_exceptionVec_0!=rhs_.io_writeback_21_bits_exceptionVec_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_exceptionVec_0=0x%0h while the rhs_.io_writeback_21_bits_exceptionVec_0=0x%0h",this.io_writeback_21_bits_exceptionVec_0,rhs_.io_writeback_21_bits_exceptionVec_0),UVM_NONE)
        end

        if(this.io_writeback_21_bits_exceptionVec_1!=rhs_.io_writeback_21_bits_exceptionVec_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_exceptionVec_1=0x%0h while the rhs_.io_writeback_21_bits_exceptionVec_1=0x%0h",this.io_writeback_21_bits_exceptionVec_1,rhs_.io_writeback_21_bits_exceptionVec_1),UVM_NONE)
        end

        if(this.io_writeback_21_bits_exceptionVec_2!=rhs_.io_writeback_21_bits_exceptionVec_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_exceptionVec_2=0x%0h while the rhs_.io_writeback_21_bits_exceptionVec_2=0x%0h",this.io_writeback_21_bits_exceptionVec_2,rhs_.io_writeback_21_bits_exceptionVec_2),UVM_NONE)
        end

        if(this.io_writeback_21_bits_exceptionVec_3!=rhs_.io_writeback_21_bits_exceptionVec_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_exceptionVec_3=0x%0h while the rhs_.io_writeback_21_bits_exceptionVec_3=0x%0h",this.io_writeback_21_bits_exceptionVec_3,rhs_.io_writeback_21_bits_exceptionVec_3),UVM_NONE)
        end

        if(this.io_writeback_21_bits_exceptionVec_4!=rhs_.io_writeback_21_bits_exceptionVec_4) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_exceptionVec_4=0x%0h while the rhs_.io_writeback_21_bits_exceptionVec_4=0x%0h",this.io_writeback_21_bits_exceptionVec_4,rhs_.io_writeback_21_bits_exceptionVec_4),UVM_NONE)
        end

        if(this.io_writeback_21_bits_exceptionVec_5!=rhs_.io_writeback_21_bits_exceptionVec_5) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_exceptionVec_5=0x%0h while the rhs_.io_writeback_21_bits_exceptionVec_5=0x%0h",this.io_writeback_21_bits_exceptionVec_5,rhs_.io_writeback_21_bits_exceptionVec_5),UVM_NONE)
        end

        if(this.io_writeback_21_bits_exceptionVec_6!=rhs_.io_writeback_21_bits_exceptionVec_6) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_exceptionVec_6=0x%0h while the rhs_.io_writeback_21_bits_exceptionVec_6=0x%0h",this.io_writeback_21_bits_exceptionVec_6,rhs_.io_writeback_21_bits_exceptionVec_6),UVM_NONE)
        end

        if(this.io_writeback_21_bits_exceptionVec_7!=rhs_.io_writeback_21_bits_exceptionVec_7) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_exceptionVec_7=0x%0h while the rhs_.io_writeback_21_bits_exceptionVec_7=0x%0h",this.io_writeback_21_bits_exceptionVec_7,rhs_.io_writeback_21_bits_exceptionVec_7),UVM_NONE)
        end

        if(this.io_writeback_21_bits_exceptionVec_8!=rhs_.io_writeback_21_bits_exceptionVec_8) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_exceptionVec_8=0x%0h while the rhs_.io_writeback_21_bits_exceptionVec_8=0x%0h",this.io_writeback_21_bits_exceptionVec_8,rhs_.io_writeback_21_bits_exceptionVec_8),UVM_NONE)
        end

        if(this.io_writeback_21_bits_exceptionVec_9!=rhs_.io_writeback_21_bits_exceptionVec_9) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_exceptionVec_9=0x%0h while the rhs_.io_writeback_21_bits_exceptionVec_9=0x%0h",this.io_writeback_21_bits_exceptionVec_9,rhs_.io_writeback_21_bits_exceptionVec_9),UVM_NONE)
        end

        if(this.io_writeback_21_bits_exceptionVec_10!=rhs_.io_writeback_21_bits_exceptionVec_10) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_exceptionVec_10=0x%0h while the rhs_.io_writeback_21_bits_exceptionVec_10=0x%0h",this.io_writeback_21_bits_exceptionVec_10,rhs_.io_writeback_21_bits_exceptionVec_10),UVM_NONE)
        end

        if(this.io_writeback_21_bits_exceptionVec_11!=rhs_.io_writeback_21_bits_exceptionVec_11) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_exceptionVec_11=0x%0h while the rhs_.io_writeback_21_bits_exceptionVec_11=0x%0h",this.io_writeback_21_bits_exceptionVec_11,rhs_.io_writeback_21_bits_exceptionVec_11),UVM_NONE)
        end

        if(this.io_writeback_21_bits_exceptionVec_12!=rhs_.io_writeback_21_bits_exceptionVec_12) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_exceptionVec_12=0x%0h while the rhs_.io_writeback_21_bits_exceptionVec_12=0x%0h",this.io_writeback_21_bits_exceptionVec_12,rhs_.io_writeback_21_bits_exceptionVec_12),UVM_NONE)
        end

        if(this.io_writeback_21_bits_exceptionVec_13!=rhs_.io_writeback_21_bits_exceptionVec_13) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_exceptionVec_13=0x%0h while the rhs_.io_writeback_21_bits_exceptionVec_13=0x%0h",this.io_writeback_21_bits_exceptionVec_13,rhs_.io_writeback_21_bits_exceptionVec_13),UVM_NONE)
        end

        if(this.io_writeback_21_bits_exceptionVec_14!=rhs_.io_writeback_21_bits_exceptionVec_14) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_exceptionVec_14=0x%0h while the rhs_.io_writeback_21_bits_exceptionVec_14=0x%0h",this.io_writeback_21_bits_exceptionVec_14,rhs_.io_writeback_21_bits_exceptionVec_14),UVM_NONE)
        end

        if(this.io_writeback_21_bits_exceptionVec_15!=rhs_.io_writeback_21_bits_exceptionVec_15) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_exceptionVec_15=0x%0h while the rhs_.io_writeback_21_bits_exceptionVec_15=0x%0h",this.io_writeback_21_bits_exceptionVec_15,rhs_.io_writeback_21_bits_exceptionVec_15),UVM_NONE)
        end

        if(this.io_writeback_21_bits_exceptionVec_16!=rhs_.io_writeback_21_bits_exceptionVec_16) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_exceptionVec_16=0x%0h while the rhs_.io_writeback_21_bits_exceptionVec_16=0x%0h",this.io_writeback_21_bits_exceptionVec_16,rhs_.io_writeback_21_bits_exceptionVec_16),UVM_NONE)
        end

        if(this.io_writeback_21_bits_exceptionVec_17!=rhs_.io_writeback_21_bits_exceptionVec_17) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_exceptionVec_17=0x%0h while the rhs_.io_writeback_21_bits_exceptionVec_17=0x%0h",this.io_writeback_21_bits_exceptionVec_17,rhs_.io_writeback_21_bits_exceptionVec_17),UVM_NONE)
        end

        if(this.io_writeback_21_bits_exceptionVec_18!=rhs_.io_writeback_21_bits_exceptionVec_18) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_exceptionVec_18=0x%0h while the rhs_.io_writeback_21_bits_exceptionVec_18=0x%0h",this.io_writeback_21_bits_exceptionVec_18,rhs_.io_writeback_21_bits_exceptionVec_18),UVM_NONE)
        end

        if(this.io_writeback_21_bits_exceptionVec_19!=rhs_.io_writeback_21_bits_exceptionVec_19) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_exceptionVec_19=0x%0h while the rhs_.io_writeback_21_bits_exceptionVec_19=0x%0h",this.io_writeback_21_bits_exceptionVec_19,rhs_.io_writeback_21_bits_exceptionVec_19),UVM_NONE)
        end

        if(this.io_writeback_21_bits_exceptionVec_20!=rhs_.io_writeback_21_bits_exceptionVec_20) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_exceptionVec_20=0x%0h while the rhs_.io_writeback_21_bits_exceptionVec_20=0x%0h",this.io_writeback_21_bits_exceptionVec_20,rhs_.io_writeback_21_bits_exceptionVec_20),UVM_NONE)
        end

        if(this.io_writeback_21_bits_exceptionVec_21!=rhs_.io_writeback_21_bits_exceptionVec_21) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_exceptionVec_21=0x%0h while the rhs_.io_writeback_21_bits_exceptionVec_21=0x%0h",this.io_writeback_21_bits_exceptionVec_21,rhs_.io_writeback_21_bits_exceptionVec_21),UVM_NONE)
        end

        if(this.io_writeback_21_bits_exceptionVec_22!=rhs_.io_writeback_21_bits_exceptionVec_22) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_exceptionVec_22=0x%0h while the rhs_.io_writeback_21_bits_exceptionVec_22=0x%0h",this.io_writeback_21_bits_exceptionVec_22,rhs_.io_writeback_21_bits_exceptionVec_22),UVM_NONE)
        end

        if(this.io_writeback_21_bits_exceptionVec_23!=rhs_.io_writeback_21_bits_exceptionVec_23) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_exceptionVec_23=0x%0h while the rhs_.io_writeback_21_bits_exceptionVec_23=0x%0h",this.io_writeback_21_bits_exceptionVec_23,rhs_.io_writeback_21_bits_exceptionVec_23),UVM_NONE)
        end

        if(this.io_writeback_21_bits_flushPipe!=rhs_.io_writeback_21_bits_flushPipe) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_flushPipe=0x%0h while the rhs_.io_writeback_21_bits_flushPipe=0x%0h",this.io_writeback_21_bits_flushPipe,rhs_.io_writeback_21_bits_flushPipe),UVM_NONE)
        end

        if(this.io_writeback_21_bits_replay!=rhs_.io_writeback_21_bits_replay) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_replay=0x%0h while the rhs_.io_writeback_21_bits_replay=0x%0h",this.io_writeback_21_bits_replay,rhs_.io_writeback_21_bits_replay),UVM_NONE)
        end

        if(this.io_writeback_21_bits_lqIdx_flag!=rhs_.io_writeback_21_bits_lqIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_lqIdx_flag=0x%0h while the rhs_.io_writeback_21_bits_lqIdx_flag=0x%0h",this.io_writeback_21_bits_lqIdx_flag,rhs_.io_writeback_21_bits_lqIdx_flag),UVM_NONE)
        end

        if(this.io_writeback_21_bits_lqIdx_value!=rhs_.io_writeback_21_bits_lqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_lqIdx_value=0x%0h while the rhs_.io_writeback_21_bits_lqIdx_value=0x%0h",this.io_writeback_21_bits_lqIdx_value,rhs_.io_writeback_21_bits_lqIdx_value),UVM_NONE)
        end

        if(this.io_writeback_21_bits_trigger!=rhs_.io_writeback_21_bits_trigger) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_trigger=0x%0h while the rhs_.io_writeback_21_bits_trigger=0x%0h",this.io_writeback_21_bits_trigger,rhs_.io_writeback_21_bits_trigger),UVM_NONE)
        end

        if(this.io_writeback_21_bits_predecodeInfo_valid!=rhs_.io_writeback_21_bits_predecodeInfo_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_predecodeInfo_valid=0x%0h while the rhs_.io_writeback_21_bits_predecodeInfo_valid=0x%0h",this.io_writeback_21_bits_predecodeInfo_valid,rhs_.io_writeback_21_bits_predecodeInfo_valid),UVM_NONE)
        end

        if(this.io_writeback_21_bits_predecodeInfo_isRVC!=rhs_.io_writeback_21_bits_predecodeInfo_isRVC) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_predecodeInfo_isRVC=0x%0h while the rhs_.io_writeback_21_bits_predecodeInfo_isRVC=0x%0h",this.io_writeback_21_bits_predecodeInfo_isRVC,rhs_.io_writeback_21_bits_predecodeInfo_isRVC),UVM_NONE)
        end

        if(this.io_writeback_21_bits_predecodeInfo_brType!=rhs_.io_writeback_21_bits_predecodeInfo_brType) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_predecodeInfo_brType=0x%0h while the rhs_.io_writeback_21_bits_predecodeInfo_brType=0x%0h",this.io_writeback_21_bits_predecodeInfo_brType,rhs_.io_writeback_21_bits_predecodeInfo_brType),UVM_NONE)
        end

        if(this.io_writeback_21_bits_predecodeInfo_isCall!=rhs_.io_writeback_21_bits_predecodeInfo_isCall) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_predecodeInfo_isCall=0x%0h while the rhs_.io_writeback_21_bits_predecodeInfo_isCall=0x%0h",this.io_writeback_21_bits_predecodeInfo_isCall,rhs_.io_writeback_21_bits_predecodeInfo_isCall),UVM_NONE)
        end

        if(this.io_writeback_21_bits_predecodeInfo_isRet!=rhs_.io_writeback_21_bits_predecodeInfo_isRet) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_predecodeInfo_isRet=0x%0h while the rhs_.io_writeback_21_bits_predecodeInfo_isRet=0x%0h",this.io_writeback_21_bits_predecodeInfo_isRet,rhs_.io_writeback_21_bits_predecodeInfo_isRet),UVM_NONE)
        end

        if(this.io_writeback_21_bits_debug_isMMIO!=rhs_.io_writeback_21_bits_debug_isMMIO) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_debug_isMMIO=0x%0h while the rhs_.io_writeback_21_bits_debug_isMMIO=0x%0h",this.io_writeback_21_bits_debug_isMMIO,rhs_.io_writeback_21_bits_debug_isMMIO),UVM_NONE)
        end

        if(this.io_writeback_21_bits_debug_isNCIO!=rhs_.io_writeback_21_bits_debug_isNCIO) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_debug_isNCIO=0x%0h while the rhs_.io_writeback_21_bits_debug_isNCIO=0x%0h",this.io_writeback_21_bits_debug_isNCIO,rhs_.io_writeback_21_bits_debug_isNCIO),UVM_NONE)
        end

        if(this.io_writeback_21_bits_debug_isPerfCnt!=rhs_.io_writeback_21_bits_debug_isPerfCnt) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_debug_isPerfCnt=0x%0h while the rhs_.io_writeback_21_bits_debug_isPerfCnt=0x%0h",this.io_writeback_21_bits_debug_isPerfCnt,rhs_.io_writeback_21_bits_debug_isPerfCnt),UVM_NONE)
        end

        if(this.io_writeback_21_bits_debug_paddr!=rhs_.io_writeback_21_bits_debug_paddr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_debug_paddr=0x%0h while the rhs_.io_writeback_21_bits_debug_paddr=0x%0h",this.io_writeback_21_bits_debug_paddr,rhs_.io_writeback_21_bits_debug_paddr),UVM_NONE)
        end

        if(this.io_writeback_21_bits_debug_vaddr!=rhs_.io_writeback_21_bits_debug_vaddr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_debug_vaddr=0x%0h while the rhs_.io_writeback_21_bits_debug_vaddr=0x%0h",this.io_writeback_21_bits_debug_vaddr,rhs_.io_writeback_21_bits_debug_vaddr),UVM_NONE)
        end

        if(this.io_writeback_21_bits_debugInfo_eliminatedMove!=rhs_.io_writeback_21_bits_debugInfo_eliminatedMove) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_debugInfo_eliminatedMove=0x%0h while the rhs_.io_writeback_21_bits_debugInfo_eliminatedMove=0x%0h",this.io_writeback_21_bits_debugInfo_eliminatedMove,rhs_.io_writeback_21_bits_debugInfo_eliminatedMove),UVM_NONE)
        end

        if(this.io_writeback_21_bits_debugInfo_renameTime!=rhs_.io_writeback_21_bits_debugInfo_renameTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_debugInfo_renameTime=0x%0h while the rhs_.io_writeback_21_bits_debugInfo_renameTime=0x%0h",this.io_writeback_21_bits_debugInfo_renameTime,rhs_.io_writeback_21_bits_debugInfo_renameTime),UVM_NONE)
        end

        if(this.io_writeback_21_bits_debugInfo_dispatchTime!=rhs_.io_writeback_21_bits_debugInfo_dispatchTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_debugInfo_dispatchTime=0x%0h while the rhs_.io_writeback_21_bits_debugInfo_dispatchTime=0x%0h",this.io_writeback_21_bits_debugInfo_dispatchTime,rhs_.io_writeback_21_bits_debugInfo_dispatchTime),UVM_NONE)
        end

        if(this.io_writeback_21_bits_debugInfo_enqRsTime!=rhs_.io_writeback_21_bits_debugInfo_enqRsTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_debugInfo_enqRsTime=0x%0h while the rhs_.io_writeback_21_bits_debugInfo_enqRsTime=0x%0h",this.io_writeback_21_bits_debugInfo_enqRsTime,rhs_.io_writeback_21_bits_debugInfo_enqRsTime),UVM_NONE)
        end

        if(this.io_writeback_21_bits_debugInfo_selectTime!=rhs_.io_writeback_21_bits_debugInfo_selectTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_debugInfo_selectTime=0x%0h while the rhs_.io_writeback_21_bits_debugInfo_selectTime=0x%0h",this.io_writeback_21_bits_debugInfo_selectTime,rhs_.io_writeback_21_bits_debugInfo_selectTime),UVM_NONE)
        end

        if(this.io_writeback_21_bits_debugInfo_issueTime!=rhs_.io_writeback_21_bits_debugInfo_issueTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_debugInfo_issueTime=0x%0h while the rhs_.io_writeback_21_bits_debugInfo_issueTime=0x%0h",this.io_writeback_21_bits_debugInfo_issueTime,rhs_.io_writeback_21_bits_debugInfo_issueTime),UVM_NONE)
        end

        if(this.io_writeback_21_bits_debugInfo_writebackTime!=rhs_.io_writeback_21_bits_debugInfo_writebackTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_debugInfo_writebackTime=0x%0h while the rhs_.io_writeback_21_bits_debugInfo_writebackTime=0x%0h",this.io_writeback_21_bits_debugInfo_writebackTime,rhs_.io_writeback_21_bits_debugInfo_writebackTime),UVM_NONE)
        end

        if(this.io_writeback_21_bits_debugInfo_runahead_checkpoint_id!=rhs_.io_writeback_21_bits_debugInfo_runahead_checkpoint_id) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_debugInfo_runahead_checkpoint_id=0x%0h while the rhs_.io_writeback_21_bits_debugInfo_runahead_checkpoint_id=0x%0h",this.io_writeback_21_bits_debugInfo_runahead_checkpoint_id,rhs_.io_writeback_21_bits_debugInfo_runahead_checkpoint_id),UVM_NONE)
        end

        if(this.io_writeback_21_bits_debugInfo_tlbFirstReqTime!=rhs_.io_writeback_21_bits_debugInfo_tlbFirstReqTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_debugInfo_tlbFirstReqTime=0x%0h while the rhs_.io_writeback_21_bits_debugInfo_tlbFirstReqTime=0x%0h",this.io_writeback_21_bits_debugInfo_tlbFirstReqTime,rhs_.io_writeback_21_bits_debugInfo_tlbFirstReqTime),UVM_NONE)
        end

        if(this.io_writeback_21_bits_debugInfo_tlbRespTime!=rhs_.io_writeback_21_bits_debugInfo_tlbRespTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_debugInfo_tlbRespTime=0x%0h while the rhs_.io_writeback_21_bits_debugInfo_tlbRespTime=0x%0h",this.io_writeback_21_bits_debugInfo_tlbRespTime,rhs_.io_writeback_21_bits_debugInfo_tlbRespTime),UVM_NONE)
        end

        if(this.io_writeback_21_bits_debug_seqNum!=rhs_.io_writeback_21_bits_debug_seqNum) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_21_bits_debug_seqNum=0x%0h while the rhs_.io_writeback_21_bits_debug_seqNum=0x%0h",this.io_writeback_21_bits_debug_seqNum,rhs_.io_writeback_21_bits_debug_seqNum),UVM_NONE)
        end

        if(this.io_writeback_20_valid!=rhs_.io_writeback_20_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_valid=0x%0h while the rhs_.io_writeback_20_valid=0x%0h",this.io_writeback_20_valid,rhs_.io_writeback_20_valid),UVM_NONE)
        end

        if(this.io_writeback_20_bits_data_0!=rhs_.io_writeback_20_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_data_0=0x%0h while the rhs_.io_writeback_20_bits_data_0=0x%0h",this.io_writeback_20_bits_data_0,rhs_.io_writeback_20_bits_data_0),UVM_NONE)
        end

        if(this.io_writeback_20_bits_pdest!=rhs_.io_writeback_20_bits_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_pdest=0x%0h while the rhs_.io_writeback_20_bits_pdest=0x%0h",this.io_writeback_20_bits_pdest,rhs_.io_writeback_20_bits_pdest),UVM_NONE)
        end

        if(this.io_writeback_20_bits_robIdx_flag!=rhs_.io_writeback_20_bits_robIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_robIdx_flag=0x%0h while the rhs_.io_writeback_20_bits_robIdx_flag=0x%0h",this.io_writeback_20_bits_robIdx_flag,rhs_.io_writeback_20_bits_robIdx_flag),UVM_NONE)
        end

        if(this.io_writeback_20_bits_robIdx_value!=rhs_.io_writeback_20_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_robIdx_value=0x%0h while the rhs_.io_writeback_20_bits_robIdx_value=0x%0h",this.io_writeback_20_bits_robIdx_value,rhs_.io_writeback_20_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_writeback_20_bits_intWen!=rhs_.io_writeback_20_bits_intWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_intWen=0x%0h while the rhs_.io_writeback_20_bits_intWen=0x%0h",this.io_writeback_20_bits_intWen,rhs_.io_writeback_20_bits_intWen),UVM_NONE)
        end

        if(this.io_writeback_20_bits_fpWen!=rhs_.io_writeback_20_bits_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_fpWen=0x%0h while the rhs_.io_writeback_20_bits_fpWen=0x%0h",this.io_writeback_20_bits_fpWen,rhs_.io_writeback_20_bits_fpWen),UVM_NONE)
        end

        if(this.io_writeback_20_bits_exceptionVec_0!=rhs_.io_writeback_20_bits_exceptionVec_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_exceptionVec_0=0x%0h while the rhs_.io_writeback_20_bits_exceptionVec_0=0x%0h",this.io_writeback_20_bits_exceptionVec_0,rhs_.io_writeback_20_bits_exceptionVec_0),UVM_NONE)
        end

        if(this.io_writeback_20_bits_exceptionVec_1!=rhs_.io_writeback_20_bits_exceptionVec_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_exceptionVec_1=0x%0h while the rhs_.io_writeback_20_bits_exceptionVec_1=0x%0h",this.io_writeback_20_bits_exceptionVec_1,rhs_.io_writeback_20_bits_exceptionVec_1),UVM_NONE)
        end

        if(this.io_writeback_20_bits_exceptionVec_2!=rhs_.io_writeback_20_bits_exceptionVec_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_exceptionVec_2=0x%0h while the rhs_.io_writeback_20_bits_exceptionVec_2=0x%0h",this.io_writeback_20_bits_exceptionVec_2,rhs_.io_writeback_20_bits_exceptionVec_2),UVM_NONE)
        end

        if(this.io_writeback_20_bits_exceptionVec_3!=rhs_.io_writeback_20_bits_exceptionVec_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_exceptionVec_3=0x%0h while the rhs_.io_writeback_20_bits_exceptionVec_3=0x%0h",this.io_writeback_20_bits_exceptionVec_3,rhs_.io_writeback_20_bits_exceptionVec_3),UVM_NONE)
        end

        if(this.io_writeback_20_bits_exceptionVec_4!=rhs_.io_writeback_20_bits_exceptionVec_4) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_exceptionVec_4=0x%0h while the rhs_.io_writeback_20_bits_exceptionVec_4=0x%0h",this.io_writeback_20_bits_exceptionVec_4,rhs_.io_writeback_20_bits_exceptionVec_4),UVM_NONE)
        end

        if(this.io_writeback_20_bits_exceptionVec_5!=rhs_.io_writeback_20_bits_exceptionVec_5) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_exceptionVec_5=0x%0h while the rhs_.io_writeback_20_bits_exceptionVec_5=0x%0h",this.io_writeback_20_bits_exceptionVec_5,rhs_.io_writeback_20_bits_exceptionVec_5),UVM_NONE)
        end

        if(this.io_writeback_20_bits_exceptionVec_6!=rhs_.io_writeback_20_bits_exceptionVec_6) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_exceptionVec_6=0x%0h while the rhs_.io_writeback_20_bits_exceptionVec_6=0x%0h",this.io_writeback_20_bits_exceptionVec_6,rhs_.io_writeback_20_bits_exceptionVec_6),UVM_NONE)
        end

        if(this.io_writeback_20_bits_exceptionVec_7!=rhs_.io_writeback_20_bits_exceptionVec_7) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_exceptionVec_7=0x%0h while the rhs_.io_writeback_20_bits_exceptionVec_7=0x%0h",this.io_writeback_20_bits_exceptionVec_7,rhs_.io_writeback_20_bits_exceptionVec_7),UVM_NONE)
        end

        if(this.io_writeback_20_bits_exceptionVec_8!=rhs_.io_writeback_20_bits_exceptionVec_8) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_exceptionVec_8=0x%0h while the rhs_.io_writeback_20_bits_exceptionVec_8=0x%0h",this.io_writeback_20_bits_exceptionVec_8,rhs_.io_writeback_20_bits_exceptionVec_8),UVM_NONE)
        end

        if(this.io_writeback_20_bits_exceptionVec_9!=rhs_.io_writeback_20_bits_exceptionVec_9) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_exceptionVec_9=0x%0h while the rhs_.io_writeback_20_bits_exceptionVec_9=0x%0h",this.io_writeback_20_bits_exceptionVec_9,rhs_.io_writeback_20_bits_exceptionVec_9),UVM_NONE)
        end

        if(this.io_writeback_20_bits_exceptionVec_10!=rhs_.io_writeback_20_bits_exceptionVec_10) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_exceptionVec_10=0x%0h while the rhs_.io_writeback_20_bits_exceptionVec_10=0x%0h",this.io_writeback_20_bits_exceptionVec_10,rhs_.io_writeback_20_bits_exceptionVec_10),UVM_NONE)
        end

        if(this.io_writeback_20_bits_exceptionVec_11!=rhs_.io_writeback_20_bits_exceptionVec_11) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_exceptionVec_11=0x%0h while the rhs_.io_writeback_20_bits_exceptionVec_11=0x%0h",this.io_writeback_20_bits_exceptionVec_11,rhs_.io_writeback_20_bits_exceptionVec_11),UVM_NONE)
        end

        if(this.io_writeback_20_bits_exceptionVec_12!=rhs_.io_writeback_20_bits_exceptionVec_12) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_exceptionVec_12=0x%0h while the rhs_.io_writeback_20_bits_exceptionVec_12=0x%0h",this.io_writeback_20_bits_exceptionVec_12,rhs_.io_writeback_20_bits_exceptionVec_12),UVM_NONE)
        end

        if(this.io_writeback_20_bits_exceptionVec_13!=rhs_.io_writeback_20_bits_exceptionVec_13) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_exceptionVec_13=0x%0h while the rhs_.io_writeback_20_bits_exceptionVec_13=0x%0h",this.io_writeback_20_bits_exceptionVec_13,rhs_.io_writeback_20_bits_exceptionVec_13),UVM_NONE)
        end

        if(this.io_writeback_20_bits_exceptionVec_14!=rhs_.io_writeback_20_bits_exceptionVec_14) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_exceptionVec_14=0x%0h while the rhs_.io_writeback_20_bits_exceptionVec_14=0x%0h",this.io_writeback_20_bits_exceptionVec_14,rhs_.io_writeback_20_bits_exceptionVec_14),UVM_NONE)
        end

        if(this.io_writeback_20_bits_exceptionVec_15!=rhs_.io_writeback_20_bits_exceptionVec_15) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_exceptionVec_15=0x%0h while the rhs_.io_writeback_20_bits_exceptionVec_15=0x%0h",this.io_writeback_20_bits_exceptionVec_15,rhs_.io_writeback_20_bits_exceptionVec_15),UVM_NONE)
        end

        if(this.io_writeback_20_bits_exceptionVec_16!=rhs_.io_writeback_20_bits_exceptionVec_16) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_exceptionVec_16=0x%0h while the rhs_.io_writeback_20_bits_exceptionVec_16=0x%0h",this.io_writeback_20_bits_exceptionVec_16,rhs_.io_writeback_20_bits_exceptionVec_16),UVM_NONE)
        end

        if(this.io_writeback_20_bits_exceptionVec_17!=rhs_.io_writeback_20_bits_exceptionVec_17) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_exceptionVec_17=0x%0h while the rhs_.io_writeback_20_bits_exceptionVec_17=0x%0h",this.io_writeback_20_bits_exceptionVec_17,rhs_.io_writeback_20_bits_exceptionVec_17),UVM_NONE)
        end

        if(this.io_writeback_20_bits_exceptionVec_18!=rhs_.io_writeback_20_bits_exceptionVec_18) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_exceptionVec_18=0x%0h while the rhs_.io_writeback_20_bits_exceptionVec_18=0x%0h",this.io_writeback_20_bits_exceptionVec_18,rhs_.io_writeback_20_bits_exceptionVec_18),UVM_NONE)
        end

        if(this.io_writeback_20_bits_exceptionVec_19!=rhs_.io_writeback_20_bits_exceptionVec_19) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_exceptionVec_19=0x%0h while the rhs_.io_writeback_20_bits_exceptionVec_19=0x%0h",this.io_writeback_20_bits_exceptionVec_19,rhs_.io_writeback_20_bits_exceptionVec_19),UVM_NONE)
        end

        if(this.io_writeback_20_bits_exceptionVec_20!=rhs_.io_writeback_20_bits_exceptionVec_20) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_exceptionVec_20=0x%0h while the rhs_.io_writeback_20_bits_exceptionVec_20=0x%0h",this.io_writeback_20_bits_exceptionVec_20,rhs_.io_writeback_20_bits_exceptionVec_20),UVM_NONE)
        end

        if(this.io_writeback_20_bits_exceptionVec_21!=rhs_.io_writeback_20_bits_exceptionVec_21) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_exceptionVec_21=0x%0h while the rhs_.io_writeback_20_bits_exceptionVec_21=0x%0h",this.io_writeback_20_bits_exceptionVec_21,rhs_.io_writeback_20_bits_exceptionVec_21),UVM_NONE)
        end

        if(this.io_writeback_20_bits_exceptionVec_22!=rhs_.io_writeback_20_bits_exceptionVec_22) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_exceptionVec_22=0x%0h while the rhs_.io_writeback_20_bits_exceptionVec_22=0x%0h",this.io_writeback_20_bits_exceptionVec_22,rhs_.io_writeback_20_bits_exceptionVec_22),UVM_NONE)
        end

        if(this.io_writeback_20_bits_exceptionVec_23!=rhs_.io_writeback_20_bits_exceptionVec_23) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_exceptionVec_23=0x%0h while the rhs_.io_writeback_20_bits_exceptionVec_23=0x%0h",this.io_writeback_20_bits_exceptionVec_23,rhs_.io_writeback_20_bits_exceptionVec_23),UVM_NONE)
        end

        if(this.io_writeback_20_bits_flushPipe!=rhs_.io_writeback_20_bits_flushPipe) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_flushPipe=0x%0h while the rhs_.io_writeback_20_bits_flushPipe=0x%0h",this.io_writeback_20_bits_flushPipe,rhs_.io_writeback_20_bits_flushPipe),UVM_NONE)
        end

        if(this.io_writeback_20_bits_replay!=rhs_.io_writeback_20_bits_replay) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_replay=0x%0h while the rhs_.io_writeback_20_bits_replay=0x%0h",this.io_writeback_20_bits_replay,rhs_.io_writeback_20_bits_replay),UVM_NONE)
        end

        if(this.io_writeback_20_bits_lqIdx_flag!=rhs_.io_writeback_20_bits_lqIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_lqIdx_flag=0x%0h while the rhs_.io_writeback_20_bits_lqIdx_flag=0x%0h",this.io_writeback_20_bits_lqIdx_flag,rhs_.io_writeback_20_bits_lqIdx_flag),UVM_NONE)
        end

        if(this.io_writeback_20_bits_lqIdx_value!=rhs_.io_writeback_20_bits_lqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_lqIdx_value=0x%0h while the rhs_.io_writeback_20_bits_lqIdx_value=0x%0h",this.io_writeback_20_bits_lqIdx_value,rhs_.io_writeback_20_bits_lqIdx_value),UVM_NONE)
        end

        if(this.io_writeback_20_bits_trigger!=rhs_.io_writeback_20_bits_trigger) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_trigger=0x%0h while the rhs_.io_writeback_20_bits_trigger=0x%0h",this.io_writeback_20_bits_trigger,rhs_.io_writeback_20_bits_trigger),UVM_NONE)
        end

        if(this.io_writeback_20_bits_predecodeInfo_valid!=rhs_.io_writeback_20_bits_predecodeInfo_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_predecodeInfo_valid=0x%0h while the rhs_.io_writeback_20_bits_predecodeInfo_valid=0x%0h",this.io_writeback_20_bits_predecodeInfo_valid,rhs_.io_writeback_20_bits_predecodeInfo_valid),UVM_NONE)
        end

        if(this.io_writeback_20_bits_predecodeInfo_isRVC!=rhs_.io_writeback_20_bits_predecodeInfo_isRVC) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_predecodeInfo_isRVC=0x%0h while the rhs_.io_writeback_20_bits_predecodeInfo_isRVC=0x%0h",this.io_writeback_20_bits_predecodeInfo_isRVC,rhs_.io_writeback_20_bits_predecodeInfo_isRVC),UVM_NONE)
        end

        if(this.io_writeback_20_bits_predecodeInfo_brType!=rhs_.io_writeback_20_bits_predecodeInfo_brType) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_predecodeInfo_brType=0x%0h while the rhs_.io_writeback_20_bits_predecodeInfo_brType=0x%0h",this.io_writeback_20_bits_predecodeInfo_brType,rhs_.io_writeback_20_bits_predecodeInfo_brType),UVM_NONE)
        end

        if(this.io_writeback_20_bits_predecodeInfo_isCall!=rhs_.io_writeback_20_bits_predecodeInfo_isCall) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_predecodeInfo_isCall=0x%0h while the rhs_.io_writeback_20_bits_predecodeInfo_isCall=0x%0h",this.io_writeback_20_bits_predecodeInfo_isCall,rhs_.io_writeback_20_bits_predecodeInfo_isCall),UVM_NONE)
        end

        if(this.io_writeback_20_bits_predecodeInfo_isRet!=rhs_.io_writeback_20_bits_predecodeInfo_isRet) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_predecodeInfo_isRet=0x%0h while the rhs_.io_writeback_20_bits_predecodeInfo_isRet=0x%0h",this.io_writeback_20_bits_predecodeInfo_isRet,rhs_.io_writeback_20_bits_predecodeInfo_isRet),UVM_NONE)
        end

        if(this.io_writeback_20_bits_debug_isMMIO!=rhs_.io_writeback_20_bits_debug_isMMIO) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_debug_isMMIO=0x%0h while the rhs_.io_writeback_20_bits_debug_isMMIO=0x%0h",this.io_writeback_20_bits_debug_isMMIO,rhs_.io_writeback_20_bits_debug_isMMIO),UVM_NONE)
        end

        if(this.io_writeback_20_bits_debug_isNCIO!=rhs_.io_writeback_20_bits_debug_isNCIO) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_debug_isNCIO=0x%0h while the rhs_.io_writeback_20_bits_debug_isNCIO=0x%0h",this.io_writeback_20_bits_debug_isNCIO,rhs_.io_writeback_20_bits_debug_isNCIO),UVM_NONE)
        end

        if(this.io_writeback_20_bits_debug_isPerfCnt!=rhs_.io_writeback_20_bits_debug_isPerfCnt) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_debug_isPerfCnt=0x%0h while the rhs_.io_writeback_20_bits_debug_isPerfCnt=0x%0h",this.io_writeback_20_bits_debug_isPerfCnt,rhs_.io_writeback_20_bits_debug_isPerfCnt),UVM_NONE)
        end

        if(this.io_writeback_20_bits_debug_paddr!=rhs_.io_writeback_20_bits_debug_paddr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_debug_paddr=0x%0h while the rhs_.io_writeback_20_bits_debug_paddr=0x%0h",this.io_writeback_20_bits_debug_paddr,rhs_.io_writeback_20_bits_debug_paddr),UVM_NONE)
        end

        if(this.io_writeback_20_bits_debug_vaddr!=rhs_.io_writeback_20_bits_debug_vaddr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_debug_vaddr=0x%0h while the rhs_.io_writeback_20_bits_debug_vaddr=0x%0h",this.io_writeback_20_bits_debug_vaddr,rhs_.io_writeback_20_bits_debug_vaddr),UVM_NONE)
        end

        if(this.io_writeback_20_bits_debugInfo_eliminatedMove!=rhs_.io_writeback_20_bits_debugInfo_eliminatedMove) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_debugInfo_eliminatedMove=0x%0h while the rhs_.io_writeback_20_bits_debugInfo_eliminatedMove=0x%0h",this.io_writeback_20_bits_debugInfo_eliminatedMove,rhs_.io_writeback_20_bits_debugInfo_eliminatedMove),UVM_NONE)
        end

        if(this.io_writeback_20_bits_debugInfo_renameTime!=rhs_.io_writeback_20_bits_debugInfo_renameTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_debugInfo_renameTime=0x%0h while the rhs_.io_writeback_20_bits_debugInfo_renameTime=0x%0h",this.io_writeback_20_bits_debugInfo_renameTime,rhs_.io_writeback_20_bits_debugInfo_renameTime),UVM_NONE)
        end

        if(this.io_writeback_20_bits_debugInfo_dispatchTime!=rhs_.io_writeback_20_bits_debugInfo_dispatchTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_debugInfo_dispatchTime=0x%0h while the rhs_.io_writeback_20_bits_debugInfo_dispatchTime=0x%0h",this.io_writeback_20_bits_debugInfo_dispatchTime,rhs_.io_writeback_20_bits_debugInfo_dispatchTime),UVM_NONE)
        end

        if(this.io_writeback_20_bits_debugInfo_enqRsTime!=rhs_.io_writeback_20_bits_debugInfo_enqRsTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_debugInfo_enqRsTime=0x%0h while the rhs_.io_writeback_20_bits_debugInfo_enqRsTime=0x%0h",this.io_writeback_20_bits_debugInfo_enqRsTime,rhs_.io_writeback_20_bits_debugInfo_enqRsTime),UVM_NONE)
        end

        if(this.io_writeback_20_bits_debugInfo_selectTime!=rhs_.io_writeback_20_bits_debugInfo_selectTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_debugInfo_selectTime=0x%0h while the rhs_.io_writeback_20_bits_debugInfo_selectTime=0x%0h",this.io_writeback_20_bits_debugInfo_selectTime,rhs_.io_writeback_20_bits_debugInfo_selectTime),UVM_NONE)
        end

        if(this.io_writeback_20_bits_debugInfo_issueTime!=rhs_.io_writeback_20_bits_debugInfo_issueTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_debugInfo_issueTime=0x%0h while the rhs_.io_writeback_20_bits_debugInfo_issueTime=0x%0h",this.io_writeback_20_bits_debugInfo_issueTime,rhs_.io_writeback_20_bits_debugInfo_issueTime),UVM_NONE)
        end

        if(this.io_writeback_20_bits_debugInfo_writebackTime!=rhs_.io_writeback_20_bits_debugInfo_writebackTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_debugInfo_writebackTime=0x%0h while the rhs_.io_writeback_20_bits_debugInfo_writebackTime=0x%0h",this.io_writeback_20_bits_debugInfo_writebackTime,rhs_.io_writeback_20_bits_debugInfo_writebackTime),UVM_NONE)
        end

        if(this.io_writeback_20_bits_debugInfo_runahead_checkpoint_id!=rhs_.io_writeback_20_bits_debugInfo_runahead_checkpoint_id) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_debugInfo_runahead_checkpoint_id=0x%0h while the rhs_.io_writeback_20_bits_debugInfo_runahead_checkpoint_id=0x%0h",this.io_writeback_20_bits_debugInfo_runahead_checkpoint_id,rhs_.io_writeback_20_bits_debugInfo_runahead_checkpoint_id),UVM_NONE)
        end

        if(this.io_writeback_20_bits_debugInfo_tlbFirstReqTime!=rhs_.io_writeback_20_bits_debugInfo_tlbFirstReqTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_debugInfo_tlbFirstReqTime=0x%0h while the rhs_.io_writeback_20_bits_debugInfo_tlbFirstReqTime=0x%0h",this.io_writeback_20_bits_debugInfo_tlbFirstReqTime,rhs_.io_writeback_20_bits_debugInfo_tlbFirstReqTime),UVM_NONE)
        end

        if(this.io_writeback_20_bits_debugInfo_tlbRespTime!=rhs_.io_writeback_20_bits_debugInfo_tlbRespTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_debugInfo_tlbRespTime=0x%0h while the rhs_.io_writeback_20_bits_debugInfo_tlbRespTime=0x%0h",this.io_writeback_20_bits_debugInfo_tlbRespTime,rhs_.io_writeback_20_bits_debugInfo_tlbRespTime),UVM_NONE)
        end

        if(this.io_writeback_20_bits_debug_seqNum!=rhs_.io_writeback_20_bits_debug_seqNum) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_20_bits_debug_seqNum=0x%0h while the rhs_.io_writeback_20_bits_debug_seqNum=0x%0h",this.io_writeback_20_bits_debug_seqNum,rhs_.io_writeback_20_bits_debug_seqNum),UVM_NONE)
        end

        if(this.io_writeback_19_valid!=rhs_.io_writeback_19_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_valid=0x%0h while the rhs_.io_writeback_19_valid=0x%0h",this.io_writeback_19_valid,rhs_.io_writeback_19_valid),UVM_NONE)
        end

        if(this.io_writeback_19_bits_data_0!=rhs_.io_writeback_19_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_data_0=0x%0h while the rhs_.io_writeback_19_bits_data_0=0x%0h",this.io_writeback_19_bits_data_0,rhs_.io_writeback_19_bits_data_0),UVM_NONE)
        end

        if(this.io_writeback_19_bits_pdest!=rhs_.io_writeback_19_bits_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_pdest=0x%0h while the rhs_.io_writeback_19_bits_pdest=0x%0h",this.io_writeback_19_bits_pdest,rhs_.io_writeback_19_bits_pdest),UVM_NONE)
        end

        if(this.io_writeback_19_bits_robIdx_flag!=rhs_.io_writeback_19_bits_robIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_robIdx_flag=0x%0h while the rhs_.io_writeback_19_bits_robIdx_flag=0x%0h",this.io_writeback_19_bits_robIdx_flag,rhs_.io_writeback_19_bits_robIdx_flag),UVM_NONE)
        end

        if(this.io_writeback_19_bits_robIdx_value!=rhs_.io_writeback_19_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_robIdx_value=0x%0h while the rhs_.io_writeback_19_bits_robIdx_value=0x%0h",this.io_writeback_19_bits_robIdx_value,rhs_.io_writeback_19_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_writeback_19_bits_intWen!=rhs_.io_writeback_19_bits_intWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_intWen=0x%0h while the rhs_.io_writeback_19_bits_intWen=0x%0h",this.io_writeback_19_bits_intWen,rhs_.io_writeback_19_bits_intWen),UVM_NONE)
        end

        if(this.io_writeback_19_bits_exceptionVec_0!=rhs_.io_writeback_19_bits_exceptionVec_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_exceptionVec_0=0x%0h while the rhs_.io_writeback_19_bits_exceptionVec_0=0x%0h",this.io_writeback_19_bits_exceptionVec_0,rhs_.io_writeback_19_bits_exceptionVec_0),UVM_NONE)
        end

        if(this.io_writeback_19_bits_exceptionVec_1!=rhs_.io_writeback_19_bits_exceptionVec_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_exceptionVec_1=0x%0h while the rhs_.io_writeback_19_bits_exceptionVec_1=0x%0h",this.io_writeback_19_bits_exceptionVec_1,rhs_.io_writeback_19_bits_exceptionVec_1),UVM_NONE)
        end

        if(this.io_writeback_19_bits_exceptionVec_2!=rhs_.io_writeback_19_bits_exceptionVec_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_exceptionVec_2=0x%0h while the rhs_.io_writeback_19_bits_exceptionVec_2=0x%0h",this.io_writeback_19_bits_exceptionVec_2,rhs_.io_writeback_19_bits_exceptionVec_2),UVM_NONE)
        end

        if(this.io_writeback_19_bits_exceptionVec_3!=rhs_.io_writeback_19_bits_exceptionVec_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_exceptionVec_3=0x%0h while the rhs_.io_writeback_19_bits_exceptionVec_3=0x%0h",this.io_writeback_19_bits_exceptionVec_3,rhs_.io_writeback_19_bits_exceptionVec_3),UVM_NONE)
        end

        if(this.io_writeback_19_bits_exceptionVec_4!=rhs_.io_writeback_19_bits_exceptionVec_4) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_exceptionVec_4=0x%0h while the rhs_.io_writeback_19_bits_exceptionVec_4=0x%0h",this.io_writeback_19_bits_exceptionVec_4,rhs_.io_writeback_19_bits_exceptionVec_4),UVM_NONE)
        end

        if(this.io_writeback_19_bits_exceptionVec_5!=rhs_.io_writeback_19_bits_exceptionVec_5) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_exceptionVec_5=0x%0h while the rhs_.io_writeback_19_bits_exceptionVec_5=0x%0h",this.io_writeback_19_bits_exceptionVec_5,rhs_.io_writeback_19_bits_exceptionVec_5),UVM_NONE)
        end

        if(this.io_writeback_19_bits_exceptionVec_6!=rhs_.io_writeback_19_bits_exceptionVec_6) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_exceptionVec_6=0x%0h while the rhs_.io_writeback_19_bits_exceptionVec_6=0x%0h",this.io_writeback_19_bits_exceptionVec_6,rhs_.io_writeback_19_bits_exceptionVec_6),UVM_NONE)
        end

        if(this.io_writeback_19_bits_exceptionVec_7!=rhs_.io_writeback_19_bits_exceptionVec_7) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_exceptionVec_7=0x%0h while the rhs_.io_writeback_19_bits_exceptionVec_7=0x%0h",this.io_writeback_19_bits_exceptionVec_7,rhs_.io_writeback_19_bits_exceptionVec_7),UVM_NONE)
        end

        if(this.io_writeback_19_bits_exceptionVec_8!=rhs_.io_writeback_19_bits_exceptionVec_8) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_exceptionVec_8=0x%0h while the rhs_.io_writeback_19_bits_exceptionVec_8=0x%0h",this.io_writeback_19_bits_exceptionVec_8,rhs_.io_writeback_19_bits_exceptionVec_8),UVM_NONE)
        end

        if(this.io_writeback_19_bits_exceptionVec_9!=rhs_.io_writeback_19_bits_exceptionVec_9) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_exceptionVec_9=0x%0h while the rhs_.io_writeback_19_bits_exceptionVec_9=0x%0h",this.io_writeback_19_bits_exceptionVec_9,rhs_.io_writeback_19_bits_exceptionVec_9),UVM_NONE)
        end

        if(this.io_writeback_19_bits_exceptionVec_10!=rhs_.io_writeback_19_bits_exceptionVec_10) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_exceptionVec_10=0x%0h while the rhs_.io_writeback_19_bits_exceptionVec_10=0x%0h",this.io_writeback_19_bits_exceptionVec_10,rhs_.io_writeback_19_bits_exceptionVec_10),UVM_NONE)
        end

        if(this.io_writeback_19_bits_exceptionVec_11!=rhs_.io_writeback_19_bits_exceptionVec_11) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_exceptionVec_11=0x%0h while the rhs_.io_writeback_19_bits_exceptionVec_11=0x%0h",this.io_writeback_19_bits_exceptionVec_11,rhs_.io_writeback_19_bits_exceptionVec_11),UVM_NONE)
        end

        if(this.io_writeback_19_bits_exceptionVec_12!=rhs_.io_writeback_19_bits_exceptionVec_12) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_exceptionVec_12=0x%0h while the rhs_.io_writeback_19_bits_exceptionVec_12=0x%0h",this.io_writeback_19_bits_exceptionVec_12,rhs_.io_writeback_19_bits_exceptionVec_12),UVM_NONE)
        end

        if(this.io_writeback_19_bits_exceptionVec_13!=rhs_.io_writeback_19_bits_exceptionVec_13) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_exceptionVec_13=0x%0h while the rhs_.io_writeback_19_bits_exceptionVec_13=0x%0h",this.io_writeback_19_bits_exceptionVec_13,rhs_.io_writeback_19_bits_exceptionVec_13),UVM_NONE)
        end

        if(this.io_writeback_19_bits_exceptionVec_14!=rhs_.io_writeback_19_bits_exceptionVec_14) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_exceptionVec_14=0x%0h while the rhs_.io_writeback_19_bits_exceptionVec_14=0x%0h",this.io_writeback_19_bits_exceptionVec_14,rhs_.io_writeback_19_bits_exceptionVec_14),UVM_NONE)
        end

        if(this.io_writeback_19_bits_exceptionVec_15!=rhs_.io_writeback_19_bits_exceptionVec_15) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_exceptionVec_15=0x%0h while the rhs_.io_writeback_19_bits_exceptionVec_15=0x%0h",this.io_writeback_19_bits_exceptionVec_15,rhs_.io_writeback_19_bits_exceptionVec_15),UVM_NONE)
        end

        if(this.io_writeback_19_bits_exceptionVec_16!=rhs_.io_writeback_19_bits_exceptionVec_16) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_exceptionVec_16=0x%0h while the rhs_.io_writeback_19_bits_exceptionVec_16=0x%0h",this.io_writeback_19_bits_exceptionVec_16,rhs_.io_writeback_19_bits_exceptionVec_16),UVM_NONE)
        end

        if(this.io_writeback_19_bits_exceptionVec_17!=rhs_.io_writeback_19_bits_exceptionVec_17) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_exceptionVec_17=0x%0h while the rhs_.io_writeback_19_bits_exceptionVec_17=0x%0h",this.io_writeback_19_bits_exceptionVec_17,rhs_.io_writeback_19_bits_exceptionVec_17),UVM_NONE)
        end

        if(this.io_writeback_19_bits_exceptionVec_18!=rhs_.io_writeback_19_bits_exceptionVec_18) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_exceptionVec_18=0x%0h while the rhs_.io_writeback_19_bits_exceptionVec_18=0x%0h",this.io_writeback_19_bits_exceptionVec_18,rhs_.io_writeback_19_bits_exceptionVec_18),UVM_NONE)
        end

        if(this.io_writeback_19_bits_exceptionVec_19!=rhs_.io_writeback_19_bits_exceptionVec_19) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_exceptionVec_19=0x%0h while the rhs_.io_writeback_19_bits_exceptionVec_19=0x%0h",this.io_writeback_19_bits_exceptionVec_19,rhs_.io_writeback_19_bits_exceptionVec_19),UVM_NONE)
        end

        if(this.io_writeback_19_bits_exceptionVec_20!=rhs_.io_writeback_19_bits_exceptionVec_20) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_exceptionVec_20=0x%0h while the rhs_.io_writeback_19_bits_exceptionVec_20=0x%0h",this.io_writeback_19_bits_exceptionVec_20,rhs_.io_writeback_19_bits_exceptionVec_20),UVM_NONE)
        end

        if(this.io_writeback_19_bits_exceptionVec_21!=rhs_.io_writeback_19_bits_exceptionVec_21) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_exceptionVec_21=0x%0h while the rhs_.io_writeback_19_bits_exceptionVec_21=0x%0h",this.io_writeback_19_bits_exceptionVec_21,rhs_.io_writeback_19_bits_exceptionVec_21),UVM_NONE)
        end

        if(this.io_writeback_19_bits_exceptionVec_22!=rhs_.io_writeback_19_bits_exceptionVec_22) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_exceptionVec_22=0x%0h while the rhs_.io_writeback_19_bits_exceptionVec_22=0x%0h",this.io_writeback_19_bits_exceptionVec_22,rhs_.io_writeback_19_bits_exceptionVec_22),UVM_NONE)
        end

        if(this.io_writeback_19_bits_exceptionVec_23!=rhs_.io_writeback_19_bits_exceptionVec_23) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_exceptionVec_23=0x%0h while the rhs_.io_writeback_19_bits_exceptionVec_23=0x%0h",this.io_writeback_19_bits_exceptionVec_23,rhs_.io_writeback_19_bits_exceptionVec_23),UVM_NONE)
        end

        if(this.io_writeback_19_bits_flushPipe!=rhs_.io_writeback_19_bits_flushPipe) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_flushPipe=0x%0h while the rhs_.io_writeback_19_bits_flushPipe=0x%0h",this.io_writeback_19_bits_flushPipe,rhs_.io_writeback_19_bits_flushPipe),UVM_NONE)
        end

        if(this.io_writeback_19_bits_sqIdx_flag!=rhs_.io_writeback_19_bits_sqIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_sqIdx_flag=0x%0h while the rhs_.io_writeback_19_bits_sqIdx_flag=0x%0h",this.io_writeback_19_bits_sqIdx_flag,rhs_.io_writeback_19_bits_sqIdx_flag),UVM_NONE)
        end

        if(this.io_writeback_19_bits_sqIdx_value!=rhs_.io_writeback_19_bits_sqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_sqIdx_value=0x%0h while the rhs_.io_writeback_19_bits_sqIdx_value=0x%0h",this.io_writeback_19_bits_sqIdx_value,rhs_.io_writeback_19_bits_sqIdx_value),UVM_NONE)
        end

        if(this.io_writeback_19_bits_trigger!=rhs_.io_writeback_19_bits_trigger) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_trigger=0x%0h while the rhs_.io_writeback_19_bits_trigger=0x%0h",this.io_writeback_19_bits_trigger,rhs_.io_writeback_19_bits_trigger),UVM_NONE)
        end

        if(this.io_writeback_19_bits_debug_isMMIO!=rhs_.io_writeback_19_bits_debug_isMMIO) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_debug_isMMIO=0x%0h while the rhs_.io_writeback_19_bits_debug_isMMIO=0x%0h",this.io_writeback_19_bits_debug_isMMIO,rhs_.io_writeback_19_bits_debug_isMMIO),UVM_NONE)
        end

        if(this.io_writeback_19_bits_debug_isNCIO!=rhs_.io_writeback_19_bits_debug_isNCIO) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_debug_isNCIO=0x%0h while the rhs_.io_writeback_19_bits_debug_isNCIO=0x%0h",this.io_writeback_19_bits_debug_isNCIO,rhs_.io_writeback_19_bits_debug_isNCIO),UVM_NONE)
        end

        if(this.io_writeback_19_bits_debug_isPerfCnt!=rhs_.io_writeback_19_bits_debug_isPerfCnt) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_debug_isPerfCnt=0x%0h while the rhs_.io_writeback_19_bits_debug_isPerfCnt=0x%0h",this.io_writeback_19_bits_debug_isPerfCnt,rhs_.io_writeback_19_bits_debug_isPerfCnt),UVM_NONE)
        end

        if(this.io_writeback_19_bits_debug_paddr!=rhs_.io_writeback_19_bits_debug_paddr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_debug_paddr=0x%0h while the rhs_.io_writeback_19_bits_debug_paddr=0x%0h",this.io_writeback_19_bits_debug_paddr,rhs_.io_writeback_19_bits_debug_paddr),UVM_NONE)
        end

        if(this.io_writeback_19_bits_debug_vaddr!=rhs_.io_writeback_19_bits_debug_vaddr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_debug_vaddr=0x%0h while the rhs_.io_writeback_19_bits_debug_vaddr=0x%0h",this.io_writeback_19_bits_debug_vaddr,rhs_.io_writeback_19_bits_debug_vaddr),UVM_NONE)
        end

        if(this.io_writeback_19_bits_debugInfo_eliminatedMove!=rhs_.io_writeback_19_bits_debugInfo_eliminatedMove) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_debugInfo_eliminatedMove=0x%0h while the rhs_.io_writeback_19_bits_debugInfo_eliminatedMove=0x%0h",this.io_writeback_19_bits_debugInfo_eliminatedMove,rhs_.io_writeback_19_bits_debugInfo_eliminatedMove),UVM_NONE)
        end

        if(this.io_writeback_19_bits_debugInfo_renameTime!=rhs_.io_writeback_19_bits_debugInfo_renameTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_debugInfo_renameTime=0x%0h while the rhs_.io_writeback_19_bits_debugInfo_renameTime=0x%0h",this.io_writeback_19_bits_debugInfo_renameTime,rhs_.io_writeback_19_bits_debugInfo_renameTime),UVM_NONE)
        end

        if(this.io_writeback_19_bits_debugInfo_dispatchTime!=rhs_.io_writeback_19_bits_debugInfo_dispatchTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_debugInfo_dispatchTime=0x%0h while the rhs_.io_writeback_19_bits_debugInfo_dispatchTime=0x%0h",this.io_writeback_19_bits_debugInfo_dispatchTime,rhs_.io_writeback_19_bits_debugInfo_dispatchTime),UVM_NONE)
        end

        if(this.io_writeback_19_bits_debugInfo_enqRsTime!=rhs_.io_writeback_19_bits_debugInfo_enqRsTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_debugInfo_enqRsTime=0x%0h while the rhs_.io_writeback_19_bits_debugInfo_enqRsTime=0x%0h",this.io_writeback_19_bits_debugInfo_enqRsTime,rhs_.io_writeback_19_bits_debugInfo_enqRsTime),UVM_NONE)
        end

        if(this.io_writeback_19_bits_debugInfo_selectTime!=rhs_.io_writeback_19_bits_debugInfo_selectTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_debugInfo_selectTime=0x%0h while the rhs_.io_writeback_19_bits_debugInfo_selectTime=0x%0h",this.io_writeback_19_bits_debugInfo_selectTime,rhs_.io_writeback_19_bits_debugInfo_selectTime),UVM_NONE)
        end

        if(this.io_writeback_19_bits_debugInfo_issueTime!=rhs_.io_writeback_19_bits_debugInfo_issueTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_debugInfo_issueTime=0x%0h while the rhs_.io_writeback_19_bits_debugInfo_issueTime=0x%0h",this.io_writeback_19_bits_debugInfo_issueTime,rhs_.io_writeback_19_bits_debugInfo_issueTime),UVM_NONE)
        end

        if(this.io_writeback_19_bits_debugInfo_writebackTime!=rhs_.io_writeback_19_bits_debugInfo_writebackTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_debugInfo_writebackTime=0x%0h while the rhs_.io_writeback_19_bits_debugInfo_writebackTime=0x%0h",this.io_writeback_19_bits_debugInfo_writebackTime,rhs_.io_writeback_19_bits_debugInfo_writebackTime),UVM_NONE)
        end

        if(this.io_writeback_19_bits_debugInfo_runahead_checkpoint_id!=rhs_.io_writeback_19_bits_debugInfo_runahead_checkpoint_id) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_debugInfo_runahead_checkpoint_id=0x%0h while the rhs_.io_writeback_19_bits_debugInfo_runahead_checkpoint_id=0x%0h",this.io_writeback_19_bits_debugInfo_runahead_checkpoint_id,rhs_.io_writeback_19_bits_debugInfo_runahead_checkpoint_id),UVM_NONE)
        end

        if(this.io_writeback_19_bits_debugInfo_tlbFirstReqTime!=rhs_.io_writeback_19_bits_debugInfo_tlbFirstReqTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_debugInfo_tlbFirstReqTime=0x%0h while the rhs_.io_writeback_19_bits_debugInfo_tlbFirstReqTime=0x%0h",this.io_writeback_19_bits_debugInfo_tlbFirstReqTime,rhs_.io_writeback_19_bits_debugInfo_tlbFirstReqTime),UVM_NONE)
        end

        if(this.io_writeback_19_bits_debugInfo_tlbRespTime!=rhs_.io_writeback_19_bits_debugInfo_tlbRespTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_debugInfo_tlbRespTime=0x%0h while the rhs_.io_writeback_19_bits_debugInfo_tlbRespTime=0x%0h",this.io_writeback_19_bits_debugInfo_tlbRespTime,rhs_.io_writeback_19_bits_debugInfo_tlbRespTime),UVM_NONE)
        end

        if(this.io_writeback_19_bits_debug_seqNum!=rhs_.io_writeback_19_bits_debug_seqNum) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_19_bits_debug_seqNum=0x%0h while the rhs_.io_writeback_19_bits_debug_seqNum=0x%0h",this.io_writeback_19_bits_debug_seqNum,rhs_.io_writeback_19_bits_debug_seqNum),UVM_NONE)
        end

        if(this.io_writeback_18_valid!=rhs_.io_writeback_18_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_valid=0x%0h while the rhs_.io_writeback_18_valid=0x%0h",this.io_writeback_18_valid,rhs_.io_writeback_18_valid),UVM_NONE)
        end

        if(this.io_writeback_18_bits_data_0!=rhs_.io_writeback_18_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_data_0=0x%0h while the rhs_.io_writeback_18_bits_data_0=0x%0h",this.io_writeback_18_bits_data_0,rhs_.io_writeback_18_bits_data_0),UVM_NONE)
        end

        if(this.io_writeback_18_bits_pdest!=rhs_.io_writeback_18_bits_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_pdest=0x%0h while the rhs_.io_writeback_18_bits_pdest=0x%0h",this.io_writeback_18_bits_pdest,rhs_.io_writeback_18_bits_pdest),UVM_NONE)
        end

        if(this.io_writeback_18_bits_robIdx_flag!=rhs_.io_writeback_18_bits_robIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_robIdx_flag=0x%0h while the rhs_.io_writeback_18_bits_robIdx_flag=0x%0h",this.io_writeback_18_bits_robIdx_flag,rhs_.io_writeback_18_bits_robIdx_flag),UVM_NONE)
        end

        if(this.io_writeback_18_bits_robIdx_value!=rhs_.io_writeback_18_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_robIdx_value=0x%0h while the rhs_.io_writeback_18_bits_robIdx_value=0x%0h",this.io_writeback_18_bits_robIdx_value,rhs_.io_writeback_18_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_writeback_18_bits_intWen!=rhs_.io_writeback_18_bits_intWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_intWen=0x%0h while the rhs_.io_writeback_18_bits_intWen=0x%0h",this.io_writeback_18_bits_intWen,rhs_.io_writeback_18_bits_intWen),UVM_NONE)
        end

        if(this.io_writeback_18_bits_exceptionVec_0!=rhs_.io_writeback_18_bits_exceptionVec_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_exceptionVec_0=0x%0h while the rhs_.io_writeback_18_bits_exceptionVec_0=0x%0h",this.io_writeback_18_bits_exceptionVec_0,rhs_.io_writeback_18_bits_exceptionVec_0),UVM_NONE)
        end

        if(this.io_writeback_18_bits_exceptionVec_1!=rhs_.io_writeback_18_bits_exceptionVec_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_exceptionVec_1=0x%0h while the rhs_.io_writeback_18_bits_exceptionVec_1=0x%0h",this.io_writeback_18_bits_exceptionVec_1,rhs_.io_writeback_18_bits_exceptionVec_1),UVM_NONE)
        end

        if(this.io_writeback_18_bits_exceptionVec_2!=rhs_.io_writeback_18_bits_exceptionVec_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_exceptionVec_2=0x%0h while the rhs_.io_writeback_18_bits_exceptionVec_2=0x%0h",this.io_writeback_18_bits_exceptionVec_2,rhs_.io_writeback_18_bits_exceptionVec_2),UVM_NONE)
        end

        if(this.io_writeback_18_bits_exceptionVec_3!=rhs_.io_writeback_18_bits_exceptionVec_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_exceptionVec_3=0x%0h while the rhs_.io_writeback_18_bits_exceptionVec_3=0x%0h",this.io_writeback_18_bits_exceptionVec_3,rhs_.io_writeback_18_bits_exceptionVec_3),UVM_NONE)
        end

        if(this.io_writeback_18_bits_exceptionVec_4!=rhs_.io_writeback_18_bits_exceptionVec_4) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_exceptionVec_4=0x%0h while the rhs_.io_writeback_18_bits_exceptionVec_4=0x%0h",this.io_writeback_18_bits_exceptionVec_4,rhs_.io_writeback_18_bits_exceptionVec_4),UVM_NONE)
        end

        if(this.io_writeback_18_bits_exceptionVec_5!=rhs_.io_writeback_18_bits_exceptionVec_5) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_exceptionVec_5=0x%0h while the rhs_.io_writeback_18_bits_exceptionVec_5=0x%0h",this.io_writeback_18_bits_exceptionVec_5,rhs_.io_writeback_18_bits_exceptionVec_5),UVM_NONE)
        end

        if(this.io_writeback_18_bits_exceptionVec_6!=rhs_.io_writeback_18_bits_exceptionVec_6) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_exceptionVec_6=0x%0h while the rhs_.io_writeback_18_bits_exceptionVec_6=0x%0h",this.io_writeback_18_bits_exceptionVec_6,rhs_.io_writeback_18_bits_exceptionVec_6),UVM_NONE)
        end

        if(this.io_writeback_18_bits_exceptionVec_7!=rhs_.io_writeback_18_bits_exceptionVec_7) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_exceptionVec_7=0x%0h while the rhs_.io_writeback_18_bits_exceptionVec_7=0x%0h",this.io_writeback_18_bits_exceptionVec_7,rhs_.io_writeback_18_bits_exceptionVec_7),UVM_NONE)
        end

        if(this.io_writeback_18_bits_exceptionVec_8!=rhs_.io_writeback_18_bits_exceptionVec_8) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_exceptionVec_8=0x%0h while the rhs_.io_writeback_18_bits_exceptionVec_8=0x%0h",this.io_writeback_18_bits_exceptionVec_8,rhs_.io_writeback_18_bits_exceptionVec_8),UVM_NONE)
        end

        if(this.io_writeback_18_bits_exceptionVec_9!=rhs_.io_writeback_18_bits_exceptionVec_9) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_exceptionVec_9=0x%0h while the rhs_.io_writeback_18_bits_exceptionVec_9=0x%0h",this.io_writeback_18_bits_exceptionVec_9,rhs_.io_writeback_18_bits_exceptionVec_9),UVM_NONE)
        end

        if(this.io_writeback_18_bits_exceptionVec_10!=rhs_.io_writeback_18_bits_exceptionVec_10) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_exceptionVec_10=0x%0h while the rhs_.io_writeback_18_bits_exceptionVec_10=0x%0h",this.io_writeback_18_bits_exceptionVec_10,rhs_.io_writeback_18_bits_exceptionVec_10),UVM_NONE)
        end

        if(this.io_writeback_18_bits_exceptionVec_11!=rhs_.io_writeback_18_bits_exceptionVec_11) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_exceptionVec_11=0x%0h while the rhs_.io_writeback_18_bits_exceptionVec_11=0x%0h",this.io_writeback_18_bits_exceptionVec_11,rhs_.io_writeback_18_bits_exceptionVec_11),UVM_NONE)
        end

        if(this.io_writeback_18_bits_exceptionVec_12!=rhs_.io_writeback_18_bits_exceptionVec_12) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_exceptionVec_12=0x%0h while the rhs_.io_writeback_18_bits_exceptionVec_12=0x%0h",this.io_writeback_18_bits_exceptionVec_12,rhs_.io_writeback_18_bits_exceptionVec_12),UVM_NONE)
        end

        if(this.io_writeback_18_bits_exceptionVec_13!=rhs_.io_writeback_18_bits_exceptionVec_13) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_exceptionVec_13=0x%0h while the rhs_.io_writeback_18_bits_exceptionVec_13=0x%0h",this.io_writeback_18_bits_exceptionVec_13,rhs_.io_writeback_18_bits_exceptionVec_13),UVM_NONE)
        end

        if(this.io_writeback_18_bits_exceptionVec_14!=rhs_.io_writeback_18_bits_exceptionVec_14) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_exceptionVec_14=0x%0h while the rhs_.io_writeback_18_bits_exceptionVec_14=0x%0h",this.io_writeback_18_bits_exceptionVec_14,rhs_.io_writeback_18_bits_exceptionVec_14),UVM_NONE)
        end

        if(this.io_writeback_18_bits_exceptionVec_15!=rhs_.io_writeback_18_bits_exceptionVec_15) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_exceptionVec_15=0x%0h while the rhs_.io_writeback_18_bits_exceptionVec_15=0x%0h",this.io_writeback_18_bits_exceptionVec_15,rhs_.io_writeback_18_bits_exceptionVec_15),UVM_NONE)
        end

        if(this.io_writeback_18_bits_exceptionVec_16!=rhs_.io_writeback_18_bits_exceptionVec_16) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_exceptionVec_16=0x%0h while the rhs_.io_writeback_18_bits_exceptionVec_16=0x%0h",this.io_writeback_18_bits_exceptionVec_16,rhs_.io_writeback_18_bits_exceptionVec_16),UVM_NONE)
        end

        if(this.io_writeback_18_bits_exceptionVec_17!=rhs_.io_writeback_18_bits_exceptionVec_17) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_exceptionVec_17=0x%0h while the rhs_.io_writeback_18_bits_exceptionVec_17=0x%0h",this.io_writeback_18_bits_exceptionVec_17,rhs_.io_writeback_18_bits_exceptionVec_17),UVM_NONE)
        end

        if(this.io_writeback_18_bits_exceptionVec_18!=rhs_.io_writeback_18_bits_exceptionVec_18) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_exceptionVec_18=0x%0h while the rhs_.io_writeback_18_bits_exceptionVec_18=0x%0h",this.io_writeback_18_bits_exceptionVec_18,rhs_.io_writeback_18_bits_exceptionVec_18),UVM_NONE)
        end

        if(this.io_writeback_18_bits_exceptionVec_19!=rhs_.io_writeback_18_bits_exceptionVec_19) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_exceptionVec_19=0x%0h while the rhs_.io_writeback_18_bits_exceptionVec_19=0x%0h",this.io_writeback_18_bits_exceptionVec_19,rhs_.io_writeback_18_bits_exceptionVec_19),UVM_NONE)
        end

        if(this.io_writeback_18_bits_exceptionVec_20!=rhs_.io_writeback_18_bits_exceptionVec_20) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_exceptionVec_20=0x%0h while the rhs_.io_writeback_18_bits_exceptionVec_20=0x%0h",this.io_writeback_18_bits_exceptionVec_20,rhs_.io_writeback_18_bits_exceptionVec_20),UVM_NONE)
        end

        if(this.io_writeback_18_bits_exceptionVec_21!=rhs_.io_writeback_18_bits_exceptionVec_21) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_exceptionVec_21=0x%0h while the rhs_.io_writeback_18_bits_exceptionVec_21=0x%0h",this.io_writeback_18_bits_exceptionVec_21,rhs_.io_writeback_18_bits_exceptionVec_21),UVM_NONE)
        end

        if(this.io_writeback_18_bits_exceptionVec_22!=rhs_.io_writeback_18_bits_exceptionVec_22) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_exceptionVec_22=0x%0h while the rhs_.io_writeback_18_bits_exceptionVec_22=0x%0h",this.io_writeback_18_bits_exceptionVec_22,rhs_.io_writeback_18_bits_exceptionVec_22),UVM_NONE)
        end

        if(this.io_writeback_18_bits_exceptionVec_23!=rhs_.io_writeback_18_bits_exceptionVec_23) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_exceptionVec_23=0x%0h while the rhs_.io_writeback_18_bits_exceptionVec_23=0x%0h",this.io_writeback_18_bits_exceptionVec_23,rhs_.io_writeback_18_bits_exceptionVec_23),UVM_NONE)
        end

        if(this.io_writeback_18_bits_flushPipe!=rhs_.io_writeback_18_bits_flushPipe) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_flushPipe=0x%0h while the rhs_.io_writeback_18_bits_flushPipe=0x%0h",this.io_writeback_18_bits_flushPipe,rhs_.io_writeback_18_bits_flushPipe),UVM_NONE)
        end

        if(this.io_writeback_18_bits_sqIdx_flag!=rhs_.io_writeback_18_bits_sqIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_sqIdx_flag=0x%0h while the rhs_.io_writeback_18_bits_sqIdx_flag=0x%0h",this.io_writeback_18_bits_sqIdx_flag,rhs_.io_writeback_18_bits_sqIdx_flag),UVM_NONE)
        end

        if(this.io_writeback_18_bits_sqIdx_value!=rhs_.io_writeback_18_bits_sqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_sqIdx_value=0x%0h while the rhs_.io_writeback_18_bits_sqIdx_value=0x%0h",this.io_writeback_18_bits_sqIdx_value,rhs_.io_writeback_18_bits_sqIdx_value),UVM_NONE)
        end

        if(this.io_writeback_18_bits_trigger!=rhs_.io_writeback_18_bits_trigger) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_trigger=0x%0h while the rhs_.io_writeback_18_bits_trigger=0x%0h",this.io_writeback_18_bits_trigger,rhs_.io_writeback_18_bits_trigger),UVM_NONE)
        end

        if(this.io_writeback_18_bits_debug_isMMIO!=rhs_.io_writeback_18_bits_debug_isMMIO) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_debug_isMMIO=0x%0h while the rhs_.io_writeback_18_bits_debug_isMMIO=0x%0h",this.io_writeback_18_bits_debug_isMMIO,rhs_.io_writeback_18_bits_debug_isMMIO),UVM_NONE)
        end

        if(this.io_writeback_18_bits_debug_isNCIO!=rhs_.io_writeback_18_bits_debug_isNCIO) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_debug_isNCIO=0x%0h while the rhs_.io_writeback_18_bits_debug_isNCIO=0x%0h",this.io_writeback_18_bits_debug_isNCIO,rhs_.io_writeback_18_bits_debug_isNCIO),UVM_NONE)
        end

        if(this.io_writeback_18_bits_debug_isPerfCnt!=rhs_.io_writeback_18_bits_debug_isPerfCnt) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_debug_isPerfCnt=0x%0h while the rhs_.io_writeback_18_bits_debug_isPerfCnt=0x%0h",this.io_writeback_18_bits_debug_isPerfCnt,rhs_.io_writeback_18_bits_debug_isPerfCnt),UVM_NONE)
        end

        if(this.io_writeback_18_bits_debug_paddr!=rhs_.io_writeback_18_bits_debug_paddr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_debug_paddr=0x%0h while the rhs_.io_writeback_18_bits_debug_paddr=0x%0h",this.io_writeback_18_bits_debug_paddr,rhs_.io_writeback_18_bits_debug_paddr),UVM_NONE)
        end

        if(this.io_writeback_18_bits_debug_vaddr!=rhs_.io_writeback_18_bits_debug_vaddr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_debug_vaddr=0x%0h while the rhs_.io_writeback_18_bits_debug_vaddr=0x%0h",this.io_writeback_18_bits_debug_vaddr,rhs_.io_writeback_18_bits_debug_vaddr),UVM_NONE)
        end

        if(this.io_writeback_18_bits_debugInfo_eliminatedMove!=rhs_.io_writeback_18_bits_debugInfo_eliminatedMove) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_debugInfo_eliminatedMove=0x%0h while the rhs_.io_writeback_18_bits_debugInfo_eliminatedMove=0x%0h",this.io_writeback_18_bits_debugInfo_eliminatedMove,rhs_.io_writeback_18_bits_debugInfo_eliminatedMove),UVM_NONE)
        end

        if(this.io_writeback_18_bits_debugInfo_renameTime!=rhs_.io_writeback_18_bits_debugInfo_renameTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_debugInfo_renameTime=0x%0h while the rhs_.io_writeback_18_bits_debugInfo_renameTime=0x%0h",this.io_writeback_18_bits_debugInfo_renameTime,rhs_.io_writeback_18_bits_debugInfo_renameTime),UVM_NONE)
        end

        if(this.io_writeback_18_bits_debugInfo_dispatchTime!=rhs_.io_writeback_18_bits_debugInfo_dispatchTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_debugInfo_dispatchTime=0x%0h while the rhs_.io_writeback_18_bits_debugInfo_dispatchTime=0x%0h",this.io_writeback_18_bits_debugInfo_dispatchTime,rhs_.io_writeback_18_bits_debugInfo_dispatchTime),UVM_NONE)
        end

        if(this.io_writeback_18_bits_debugInfo_enqRsTime!=rhs_.io_writeback_18_bits_debugInfo_enqRsTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_debugInfo_enqRsTime=0x%0h while the rhs_.io_writeback_18_bits_debugInfo_enqRsTime=0x%0h",this.io_writeback_18_bits_debugInfo_enqRsTime,rhs_.io_writeback_18_bits_debugInfo_enqRsTime),UVM_NONE)
        end

        if(this.io_writeback_18_bits_debugInfo_selectTime!=rhs_.io_writeback_18_bits_debugInfo_selectTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_debugInfo_selectTime=0x%0h while the rhs_.io_writeback_18_bits_debugInfo_selectTime=0x%0h",this.io_writeback_18_bits_debugInfo_selectTime,rhs_.io_writeback_18_bits_debugInfo_selectTime),UVM_NONE)
        end

        if(this.io_writeback_18_bits_debugInfo_issueTime!=rhs_.io_writeback_18_bits_debugInfo_issueTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_debugInfo_issueTime=0x%0h while the rhs_.io_writeback_18_bits_debugInfo_issueTime=0x%0h",this.io_writeback_18_bits_debugInfo_issueTime,rhs_.io_writeback_18_bits_debugInfo_issueTime),UVM_NONE)
        end

        if(this.io_writeback_18_bits_debugInfo_writebackTime!=rhs_.io_writeback_18_bits_debugInfo_writebackTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_debugInfo_writebackTime=0x%0h while the rhs_.io_writeback_18_bits_debugInfo_writebackTime=0x%0h",this.io_writeback_18_bits_debugInfo_writebackTime,rhs_.io_writeback_18_bits_debugInfo_writebackTime),UVM_NONE)
        end

        if(this.io_writeback_18_bits_debugInfo_runahead_checkpoint_id!=rhs_.io_writeback_18_bits_debugInfo_runahead_checkpoint_id) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_debugInfo_runahead_checkpoint_id=0x%0h while the rhs_.io_writeback_18_bits_debugInfo_runahead_checkpoint_id=0x%0h",this.io_writeback_18_bits_debugInfo_runahead_checkpoint_id,rhs_.io_writeback_18_bits_debugInfo_runahead_checkpoint_id),UVM_NONE)
        end

        if(this.io_writeback_18_bits_debugInfo_tlbFirstReqTime!=rhs_.io_writeback_18_bits_debugInfo_tlbFirstReqTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_debugInfo_tlbFirstReqTime=0x%0h while the rhs_.io_writeback_18_bits_debugInfo_tlbFirstReqTime=0x%0h",this.io_writeback_18_bits_debugInfo_tlbFirstReqTime,rhs_.io_writeback_18_bits_debugInfo_tlbFirstReqTime),UVM_NONE)
        end

        if(this.io_writeback_18_bits_debugInfo_tlbRespTime!=rhs_.io_writeback_18_bits_debugInfo_tlbRespTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_debugInfo_tlbRespTime=0x%0h while the rhs_.io_writeback_18_bits_debugInfo_tlbRespTime=0x%0h",this.io_writeback_18_bits_debugInfo_tlbRespTime,rhs_.io_writeback_18_bits_debugInfo_tlbRespTime),UVM_NONE)
        end

        if(this.io_writeback_18_bits_debug_seqNum!=rhs_.io_writeback_18_bits_debug_seqNum) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_18_bits_debug_seqNum=0x%0h while the rhs_.io_writeback_18_bits_debug_seqNum=0x%0h",this.io_writeback_18_bits_debug_seqNum,rhs_.io_writeback_18_bits_debug_seqNum),UVM_NONE)
        end

        if(this.io_writeback_17_valid!=rhs_.io_writeback_17_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_17_valid=0x%0h while the rhs_.io_writeback_17_valid=0x%0h",this.io_writeback_17_valid,rhs_.io_writeback_17_valid),UVM_NONE)
        end

        if(this.io_writeback_17_bits_data_0!=rhs_.io_writeback_17_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_17_bits_data_0=0x%0h while the rhs_.io_writeback_17_bits_data_0=0x%0h",this.io_writeback_17_bits_data_0,rhs_.io_writeback_17_bits_data_0),UVM_NONE)
        end

        if(this.io_writeback_17_bits_data_1!=rhs_.io_writeback_17_bits_data_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_17_bits_data_1=0x%0h while the rhs_.io_writeback_17_bits_data_1=0x%0h",this.io_writeback_17_bits_data_1,rhs_.io_writeback_17_bits_data_1),UVM_NONE)
        end

        if(this.io_writeback_17_bits_data_2!=rhs_.io_writeback_17_bits_data_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_17_bits_data_2=0x%0h while the rhs_.io_writeback_17_bits_data_2=0x%0h",this.io_writeback_17_bits_data_2,rhs_.io_writeback_17_bits_data_2),UVM_NONE)
        end

        if(this.io_writeback_17_bits_pdest!=rhs_.io_writeback_17_bits_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_17_bits_pdest=0x%0h while the rhs_.io_writeback_17_bits_pdest=0x%0h",this.io_writeback_17_bits_pdest,rhs_.io_writeback_17_bits_pdest),UVM_NONE)
        end

        if(this.io_writeback_17_bits_robIdx_flag!=rhs_.io_writeback_17_bits_robIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_17_bits_robIdx_flag=0x%0h while the rhs_.io_writeback_17_bits_robIdx_flag=0x%0h",this.io_writeback_17_bits_robIdx_flag,rhs_.io_writeback_17_bits_robIdx_flag),UVM_NONE)
        end

        if(this.io_writeback_17_bits_robIdx_value!=rhs_.io_writeback_17_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_17_bits_robIdx_value=0x%0h while the rhs_.io_writeback_17_bits_robIdx_value=0x%0h",this.io_writeback_17_bits_robIdx_value,rhs_.io_writeback_17_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_writeback_17_bits_vecWen!=rhs_.io_writeback_17_bits_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_17_bits_vecWen=0x%0h while the rhs_.io_writeback_17_bits_vecWen=0x%0h",this.io_writeback_17_bits_vecWen,rhs_.io_writeback_17_bits_vecWen),UVM_NONE)
        end

        if(this.io_writeback_17_bits_v0Wen!=rhs_.io_writeback_17_bits_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_17_bits_v0Wen=0x%0h while the rhs_.io_writeback_17_bits_v0Wen=0x%0h",this.io_writeback_17_bits_v0Wen,rhs_.io_writeback_17_bits_v0Wen),UVM_NONE)
        end

        if(this.io_writeback_17_bits_fflags!=rhs_.io_writeback_17_bits_fflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_17_bits_fflags=0x%0h while the rhs_.io_writeback_17_bits_fflags=0x%0h",this.io_writeback_17_bits_fflags,rhs_.io_writeback_17_bits_fflags),UVM_NONE)
        end

        if(this.io_writeback_17_bits_wflags!=rhs_.io_writeback_17_bits_wflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_17_bits_wflags=0x%0h while the rhs_.io_writeback_17_bits_wflags=0x%0h",this.io_writeback_17_bits_wflags,rhs_.io_writeback_17_bits_wflags),UVM_NONE)
        end

        if(this.io_writeback_17_bits_debugInfo_eliminatedMove!=rhs_.io_writeback_17_bits_debugInfo_eliminatedMove) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_17_bits_debugInfo_eliminatedMove=0x%0h while the rhs_.io_writeback_17_bits_debugInfo_eliminatedMove=0x%0h",this.io_writeback_17_bits_debugInfo_eliminatedMove,rhs_.io_writeback_17_bits_debugInfo_eliminatedMove),UVM_NONE)
        end

        if(this.io_writeback_17_bits_debugInfo_renameTime!=rhs_.io_writeback_17_bits_debugInfo_renameTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_17_bits_debugInfo_renameTime=0x%0h while the rhs_.io_writeback_17_bits_debugInfo_renameTime=0x%0h",this.io_writeback_17_bits_debugInfo_renameTime,rhs_.io_writeback_17_bits_debugInfo_renameTime),UVM_NONE)
        end

        if(this.io_writeback_17_bits_debugInfo_dispatchTime!=rhs_.io_writeback_17_bits_debugInfo_dispatchTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_17_bits_debugInfo_dispatchTime=0x%0h while the rhs_.io_writeback_17_bits_debugInfo_dispatchTime=0x%0h",this.io_writeback_17_bits_debugInfo_dispatchTime,rhs_.io_writeback_17_bits_debugInfo_dispatchTime),UVM_NONE)
        end

        if(this.io_writeback_17_bits_debugInfo_enqRsTime!=rhs_.io_writeback_17_bits_debugInfo_enqRsTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_17_bits_debugInfo_enqRsTime=0x%0h while the rhs_.io_writeback_17_bits_debugInfo_enqRsTime=0x%0h",this.io_writeback_17_bits_debugInfo_enqRsTime,rhs_.io_writeback_17_bits_debugInfo_enqRsTime),UVM_NONE)
        end

        if(this.io_writeback_17_bits_debugInfo_selectTime!=rhs_.io_writeback_17_bits_debugInfo_selectTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_17_bits_debugInfo_selectTime=0x%0h while the rhs_.io_writeback_17_bits_debugInfo_selectTime=0x%0h",this.io_writeback_17_bits_debugInfo_selectTime,rhs_.io_writeback_17_bits_debugInfo_selectTime),UVM_NONE)
        end

        if(this.io_writeback_17_bits_debugInfo_issueTime!=rhs_.io_writeback_17_bits_debugInfo_issueTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_17_bits_debugInfo_issueTime=0x%0h while the rhs_.io_writeback_17_bits_debugInfo_issueTime=0x%0h",this.io_writeback_17_bits_debugInfo_issueTime,rhs_.io_writeback_17_bits_debugInfo_issueTime),UVM_NONE)
        end

        if(this.io_writeback_17_bits_debugInfo_writebackTime!=rhs_.io_writeback_17_bits_debugInfo_writebackTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_17_bits_debugInfo_writebackTime=0x%0h while the rhs_.io_writeback_17_bits_debugInfo_writebackTime=0x%0h",this.io_writeback_17_bits_debugInfo_writebackTime,rhs_.io_writeback_17_bits_debugInfo_writebackTime),UVM_NONE)
        end

        if(this.io_writeback_17_bits_debugInfo_runahead_checkpoint_id!=rhs_.io_writeback_17_bits_debugInfo_runahead_checkpoint_id) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_17_bits_debugInfo_runahead_checkpoint_id=0x%0h while the rhs_.io_writeback_17_bits_debugInfo_runahead_checkpoint_id=0x%0h",this.io_writeback_17_bits_debugInfo_runahead_checkpoint_id,rhs_.io_writeback_17_bits_debugInfo_runahead_checkpoint_id),UVM_NONE)
        end

        if(this.io_writeback_17_bits_debugInfo_tlbFirstReqTime!=rhs_.io_writeback_17_bits_debugInfo_tlbFirstReqTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_17_bits_debugInfo_tlbFirstReqTime=0x%0h while the rhs_.io_writeback_17_bits_debugInfo_tlbFirstReqTime=0x%0h",this.io_writeback_17_bits_debugInfo_tlbFirstReqTime,rhs_.io_writeback_17_bits_debugInfo_tlbFirstReqTime),UVM_NONE)
        end

        if(this.io_writeback_17_bits_debugInfo_tlbRespTime!=rhs_.io_writeback_17_bits_debugInfo_tlbRespTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_17_bits_debugInfo_tlbRespTime=0x%0h while the rhs_.io_writeback_17_bits_debugInfo_tlbRespTime=0x%0h",this.io_writeback_17_bits_debugInfo_tlbRespTime,rhs_.io_writeback_17_bits_debugInfo_tlbRespTime),UVM_NONE)
        end

        if(this.io_writeback_17_bits_debug_seqNum!=rhs_.io_writeback_17_bits_debug_seqNum) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_17_bits_debug_seqNum=0x%0h while the rhs_.io_writeback_17_bits_debug_seqNum=0x%0h",this.io_writeback_17_bits_debug_seqNum,rhs_.io_writeback_17_bits_debug_seqNum),UVM_NONE)
        end

        if(this.io_writeback_16_valid!=rhs_.io_writeback_16_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_16_valid=0x%0h while the rhs_.io_writeback_16_valid=0x%0h",this.io_writeback_16_valid,rhs_.io_writeback_16_valid),UVM_NONE)
        end

        if(this.io_writeback_16_bits_data_0!=rhs_.io_writeback_16_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_16_bits_data_0=0x%0h while the rhs_.io_writeback_16_bits_data_0=0x%0h",this.io_writeback_16_bits_data_0,rhs_.io_writeback_16_bits_data_0),UVM_NONE)
        end

        if(this.io_writeback_16_bits_data_1!=rhs_.io_writeback_16_bits_data_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_16_bits_data_1=0x%0h while the rhs_.io_writeback_16_bits_data_1=0x%0h",this.io_writeback_16_bits_data_1,rhs_.io_writeback_16_bits_data_1),UVM_NONE)
        end

        if(this.io_writeback_16_bits_data_2!=rhs_.io_writeback_16_bits_data_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_16_bits_data_2=0x%0h while the rhs_.io_writeback_16_bits_data_2=0x%0h",this.io_writeback_16_bits_data_2,rhs_.io_writeback_16_bits_data_2),UVM_NONE)
        end

        if(this.io_writeback_16_bits_data_3!=rhs_.io_writeback_16_bits_data_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_16_bits_data_3=0x%0h while the rhs_.io_writeback_16_bits_data_3=0x%0h",this.io_writeback_16_bits_data_3,rhs_.io_writeback_16_bits_data_3),UVM_NONE)
        end

        if(this.io_writeback_16_bits_pdest!=rhs_.io_writeback_16_bits_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_16_bits_pdest=0x%0h while the rhs_.io_writeback_16_bits_pdest=0x%0h",this.io_writeback_16_bits_pdest,rhs_.io_writeback_16_bits_pdest),UVM_NONE)
        end

        if(this.io_writeback_16_bits_robIdx_flag!=rhs_.io_writeback_16_bits_robIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_16_bits_robIdx_flag=0x%0h while the rhs_.io_writeback_16_bits_robIdx_flag=0x%0h",this.io_writeback_16_bits_robIdx_flag,rhs_.io_writeback_16_bits_robIdx_flag),UVM_NONE)
        end

        if(this.io_writeback_16_bits_robIdx_value!=rhs_.io_writeback_16_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_16_bits_robIdx_value=0x%0h while the rhs_.io_writeback_16_bits_robIdx_value=0x%0h",this.io_writeback_16_bits_robIdx_value,rhs_.io_writeback_16_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_writeback_16_bits_fpWen!=rhs_.io_writeback_16_bits_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_16_bits_fpWen=0x%0h while the rhs_.io_writeback_16_bits_fpWen=0x%0h",this.io_writeback_16_bits_fpWen,rhs_.io_writeback_16_bits_fpWen),UVM_NONE)
        end

        if(this.io_writeback_16_bits_vecWen!=rhs_.io_writeback_16_bits_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_16_bits_vecWen=0x%0h while the rhs_.io_writeback_16_bits_vecWen=0x%0h",this.io_writeback_16_bits_vecWen,rhs_.io_writeback_16_bits_vecWen),UVM_NONE)
        end

        if(this.io_writeback_16_bits_v0Wen!=rhs_.io_writeback_16_bits_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_16_bits_v0Wen=0x%0h while the rhs_.io_writeback_16_bits_v0Wen=0x%0h",this.io_writeback_16_bits_v0Wen,rhs_.io_writeback_16_bits_v0Wen),UVM_NONE)
        end

        if(this.io_writeback_16_bits_fflags!=rhs_.io_writeback_16_bits_fflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_16_bits_fflags=0x%0h while the rhs_.io_writeback_16_bits_fflags=0x%0h",this.io_writeback_16_bits_fflags,rhs_.io_writeback_16_bits_fflags),UVM_NONE)
        end

        if(this.io_writeback_16_bits_wflags!=rhs_.io_writeback_16_bits_wflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_16_bits_wflags=0x%0h while the rhs_.io_writeback_16_bits_wflags=0x%0h",this.io_writeback_16_bits_wflags,rhs_.io_writeback_16_bits_wflags),UVM_NONE)
        end

        if(this.io_writeback_16_bits_debugInfo_eliminatedMove!=rhs_.io_writeback_16_bits_debugInfo_eliminatedMove) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_16_bits_debugInfo_eliminatedMove=0x%0h while the rhs_.io_writeback_16_bits_debugInfo_eliminatedMove=0x%0h",this.io_writeback_16_bits_debugInfo_eliminatedMove,rhs_.io_writeback_16_bits_debugInfo_eliminatedMove),UVM_NONE)
        end

        if(this.io_writeback_16_bits_debugInfo_renameTime!=rhs_.io_writeback_16_bits_debugInfo_renameTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_16_bits_debugInfo_renameTime=0x%0h while the rhs_.io_writeback_16_bits_debugInfo_renameTime=0x%0h",this.io_writeback_16_bits_debugInfo_renameTime,rhs_.io_writeback_16_bits_debugInfo_renameTime),UVM_NONE)
        end

        if(this.io_writeback_16_bits_debugInfo_dispatchTime!=rhs_.io_writeback_16_bits_debugInfo_dispatchTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_16_bits_debugInfo_dispatchTime=0x%0h while the rhs_.io_writeback_16_bits_debugInfo_dispatchTime=0x%0h",this.io_writeback_16_bits_debugInfo_dispatchTime,rhs_.io_writeback_16_bits_debugInfo_dispatchTime),UVM_NONE)
        end

        if(this.io_writeback_16_bits_debugInfo_enqRsTime!=rhs_.io_writeback_16_bits_debugInfo_enqRsTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_16_bits_debugInfo_enqRsTime=0x%0h while the rhs_.io_writeback_16_bits_debugInfo_enqRsTime=0x%0h",this.io_writeback_16_bits_debugInfo_enqRsTime,rhs_.io_writeback_16_bits_debugInfo_enqRsTime),UVM_NONE)
        end

        if(this.io_writeback_16_bits_debugInfo_selectTime!=rhs_.io_writeback_16_bits_debugInfo_selectTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_16_bits_debugInfo_selectTime=0x%0h while the rhs_.io_writeback_16_bits_debugInfo_selectTime=0x%0h",this.io_writeback_16_bits_debugInfo_selectTime,rhs_.io_writeback_16_bits_debugInfo_selectTime),UVM_NONE)
        end

        if(this.io_writeback_16_bits_debugInfo_issueTime!=rhs_.io_writeback_16_bits_debugInfo_issueTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_16_bits_debugInfo_issueTime=0x%0h while the rhs_.io_writeback_16_bits_debugInfo_issueTime=0x%0h",this.io_writeback_16_bits_debugInfo_issueTime,rhs_.io_writeback_16_bits_debugInfo_issueTime),UVM_NONE)
        end

        if(this.io_writeback_16_bits_debugInfo_writebackTime!=rhs_.io_writeback_16_bits_debugInfo_writebackTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_16_bits_debugInfo_writebackTime=0x%0h while the rhs_.io_writeback_16_bits_debugInfo_writebackTime=0x%0h",this.io_writeback_16_bits_debugInfo_writebackTime,rhs_.io_writeback_16_bits_debugInfo_writebackTime),UVM_NONE)
        end

        if(this.io_writeback_16_bits_debugInfo_runahead_checkpoint_id!=rhs_.io_writeback_16_bits_debugInfo_runahead_checkpoint_id) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_16_bits_debugInfo_runahead_checkpoint_id=0x%0h while the rhs_.io_writeback_16_bits_debugInfo_runahead_checkpoint_id=0x%0h",this.io_writeback_16_bits_debugInfo_runahead_checkpoint_id,rhs_.io_writeback_16_bits_debugInfo_runahead_checkpoint_id),UVM_NONE)
        end

        if(this.io_writeback_16_bits_debugInfo_tlbFirstReqTime!=rhs_.io_writeback_16_bits_debugInfo_tlbFirstReqTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_16_bits_debugInfo_tlbFirstReqTime=0x%0h while the rhs_.io_writeback_16_bits_debugInfo_tlbFirstReqTime=0x%0h",this.io_writeback_16_bits_debugInfo_tlbFirstReqTime,rhs_.io_writeback_16_bits_debugInfo_tlbFirstReqTime),UVM_NONE)
        end

        if(this.io_writeback_16_bits_debugInfo_tlbRespTime!=rhs_.io_writeback_16_bits_debugInfo_tlbRespTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_16_bits_debugInfo_tlbRespTime=0x%0h while the rhs_.io_writeback_16_bits_debugInfo_tlbRespTime=0x%0h",this.io_writeback_16_bits_debugInfo_tlbRespTime,rhs_.io_writeback_16_bits_debugInfo_tlbRespTime),UVM_NONE)
        end

        if(this.io_writeback_16_bits_debug_seqNum!=rhs_.io_writeback_16_bits_debug_seqNum) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_16_bits_debug_seqNum=0x%0h while the rhs_.io_writeback_16_bits_debug_seqNum=0x%0h",this.io_writeback_16_bits_debug_seqNum,rhs_.io_writeback_16_bits_debug_seqNum),UVM_NONE)
        end

        if(this.io_writeback_15_valid!=rhs_.io_writeback_15_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_15_valid=0x%0h while the rhs_.io_writeback_15_valid=0x%0h",this.io_writeback_15_valid,rhs_.io_writeback_15_valid),UVM_NONE)
        end

        if(this.io_writeback_15_bits_data_0!=rhs_.io_writeback_15_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_15_bits_data_0=0x%0h while the rhs_.io_writeback_15_bits_data_0=0x%0h",this.io_writeback_15_bits_data_0,rhs_.io_writeback_15_bits_data_0),UVM_NONE)
        end

        if(this.io_writeback_15_bits_data_1!=rhs_.io_writeback_15_bits_data_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_15_bits_data_1=0x%0h while the rhs_.io_writeback_15_bits_data_1=0x%0h",this.io_writeback_15_bits_data_1,rhs_.io_writeback_15_bits_data_1),UVM_NONE)
        end

        if(this.io_writeback_15_bits_data_2!=rhs_.io_writeback_15_bits_data_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_15_bits_data_2=0x%0h while the rhs_.io_writeback_15_bits_data_2=0x%0h",this.io_writeback_15_bits_data_2,rhs_.io_writeback_15_bits_data_2),UVM_NONE)
        end

        if(this.io_writeback_15_bits_pdest!=rhs_.io_writeback_15_bits_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_15_bits_pdest=0x%0h while the rhs_.io_writeback_15_bits_pdest=0x%0h",this.io_writeback_15_bits_pdest,rhs_.io_writeback_15_bits_pdest),UVM_NONE)
        end

        if(this.io_writeback_15_bits_robIdx_flag!=rhs_.io_writeback_15_bits_robIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_15_bits_robIdx_flag=0x%0h while the rhs_.io_writeback_15_bits_robIdx_flag=0x%0h",this.io_writeback_15_bits_robIdx_flag,rhs_.io_writeback_15_bits_robIdx_flag),UVM_NONE)
        end

        if(this.io_writeback_15_bits_robIdx_value!=rhs_.io_writeback_15_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_15_bits_robIdx_value=0x%0h while the rhs_.io_writeback_15_bits_robIdx_value=0x%0h",this.io_writeback_15_bits_robIdx_value,rhs_.io_writeback_15_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_writeback_15_bits_vecWen!=rhs_.io_writeback_15_bits_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_15_bits_vecWen=0x%0h while the rhs_.io_writeback_15_bits_vecWen=0x%0h",this.io_writeback_15_bits_vecWen,rhs_.io_writeback_15_bits_vecWen),UVM_NONE)
        end

        if(this.io_writeback_15_bits_v0Wen!=rhs_.io_writeback_15_bits_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_15_bits_v0Wen=0x%0h while the rhs_.io_writeback_15_bits_v0Wen=0x%0h",this.io_writeback_15_bits_v0Wen,rhs_.io_writeback_15_bits_v0Wen),UVM_NONE)
        end

        if(this.io_writeback_15_bits_fflags!=rhs_.io_writeback_15_bits_fflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_15_bits_fflags=0x%0h while the rhs_.io_writeback_15_bits_fflags=0x%0h",this.io_writeback_15_bits_fflags,rhs_.io_writeback_15_bits_fflags),UVM_NONE)
        end

        if(this.io_writeback_15_bits_wflags!=rhs_.io_writeback_15_bits_wflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_15_bits_wflags=0x%0h while the rhs_.io_writeback_15_bits_wflags=0x%0h",this.io_writeback_15_bits_wflags,rhs_.io_writeback_15_bits_wflags),UVM_NONE)
        end

        if(this.io_writeback_15_bits_vxsat!=rhs_.io_writeback_15_bits_vxsat) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_15_bits_vxsat=0x%0h while the rhs_.io_writeback_15_bits_vxsat=0x%0h",this.io_writeback_15_bits_vxsat,rhs_.io_writeback_15_bits_vxsat),UVM_NONE)
        end

        if(this.io_writeback_15_bits_debugInfo_eliminatedMove!=rhs_.io_writeback_15_bits_debugInfo_eliminatedMove) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_15_bits_debugInfo_eliminatedMove=0x%0h while the rhs_.io_writeback_15_bits_debugInfo_eliminatedMove=0x%0h",this.io_writeback_15_bits_debugInfo_eliminatedMove,rhs_.io_writeback_15_bits_debugInfo_eliminatedMove),UVM_NONE)
        end

        if(this.io_writeback_15_bits_debugInfo_renameTime!=rhs_.io_writeback_15_bits_debugInfo_renameTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_15_bits_debugInfo_renameTime=0x%0h while the rhs_.io_writeback_15_bits_debugInfo_renameTime=0x%0h",this.io_writeback_15_bits_debugInfo_renameTime,rhs_.io_writeback_15_bits_debugInfo_renameTime),UVM_NONE)
        end

        if(this.io_writeback_15_bits_debugInfo_dispatchTime!=rhs_.io_writeback_15_bits_debugInfo_dispatchTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_15_bits_debugInfo_dispatchTime=0x%0h while the rhs_.io_writeback_15_bits_debugInfo_dispatchTime=0x%0h",this.io_writeback_15_bits_debugInfo_dispatchTime,rhs_.io_writeback_15_bits_debugInfo_dispatchTime),UVM_NONE)
        end

        if(this.io_writeback_15_bits_debugInfo_enqRsTime!=rhs_.io_writeback_15_bits_debugInfo_enqRsTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_15_bits_debugInfo_enqRsTime=0x%0h while the rhs_.io_writeback_15_bits_debugInfo_enqRsTime=0x%0h",this.io_writeback_15_bits_debugInfo_enqRsTime,rhs_.io_writeback_15_bits_debugInfo_enqRsTime),UVM_NONE)
        end

        if(this.io_writeback_15_bits_debugInfo_selectTime!=rhs_.io_writeback_15_bits_debugInfo_selectTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_15_bits_debugInfo_selectTime=0x%0h while the rhs_.io_writeback_15_bits_debugInfo_selectTime=0x%0h",this.io_writeback_15_bits_debugInfo_selectTime,rhs_.io_writeback_15_bits_debugInfo_selectTime),UVM_NONE)
        end

        if(this.io_writeback_15_bits_debugInfo_issueTime!=rhs_.io_writeback_15_bits_debugInfo_issueTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_15_bits_debugInfo_issueTime=0x%0h while the rhs_.io_writeback_15_bits_debugInfo_issueTime=0x%0h",this.io_writeback_15_bits_debugInfo_issueTime,rhs_.io_writeback_15_bits_debugInfo_issueTime),UVM_NONE)
        end

        if(this.io_writeback_15_bits_debugInfo_writebackTime!=rhs_.io_writeback_15_bits_debugInfo_writebackTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_15_bits_debugInfo_writebackTime=0x%0h while the rhs_.io_writeback_15_bits_debugInfo_writebackTime=0x%0h",this.io_writeback_15_bits_debugInfo_writebackTime,rhs_.io_writeback_15_bits_debugInfo_writebackTime),UVM_NONE)
        end

        if(this.io_writeback_15_bits_debugInfo_runahead_checkpoint_id!=rhs_.io_writeback_15_bits_debugInfo_runahead_checkpoint_id) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_15_bits_debugInfo_runahead_checkpoint_id=0x%0h while the rhs_.io_writeback_15_bits_debugInfo_runahead_checkpoint_id=0x%0h",this.io_writeback_15_bits_debugInfo_runahead_checkpoint_id,rhs_.io_writeback_15_bits_debugInfo_runahead_checkpoint_id),UVM_NONE)
        end

        if(this.io_writeback_15_bits_debugInfo_tlbFirstReqTime!=rhs_.io_writeback_15_bits_debugInfo_tlbFirstReqTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_15_bits_debugInfo_tlbFirstReqTime=0x%0h while the rhs_.io_writeback_15_bits_debugInfo_tlbFirstReqTime=0x%0h",this.io_writeback_15_bits_debugInfo_tlbFirstReqTime,rhs_.io_writeback_15_bits_debugInfo_tlbFirstReqTime),UVM_NONE)
        end

        if(this.io_writeback_15_bits_debugInfo_tlbRespTime!=rhs_.io_writeback_15_bits_debugInfo_tlbRespTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_15_bits_debugInfo_tlbRespTime=0x%0h while the rhs_.io_writeback_15_bits_debugInfo_tlbRespTime=0x%0h",this.io_writeback_15_bits_debugInfo_tlbRespTime,rhs_.io_writeback_15_bits_debugInfo_tlbRespTime),UVM_NONE)
        end

        if(this.io_writeback_15_bits_debug_seqNum!=rhs_.io_writeback_15_bits_debug_seqNum) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_15_bits_debug_seqNum=0x%0h while the rhs_.io_writeback_15_bits_debug_seqNum=0x%0h",this.io_writeback_15_bits_debug_seqNum,rhs_.io_writeback_15_bits_debug_seqNum),UVM_NONE)
        end

        if(this.io_writeback_14_valid!=rhs_.io_writeback_14_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_valid=0x%0h while the rhs_.io_writeback_14_valid=0x%0h",this.io_writeback_14_valid,rhs_.io_writeback_14_valid),UVM_NONE)
        end

        if(this.io_writeback_14_bits_data_0!=rhs_.io_writeback_14_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_bits_data_0=0x%0h while the rhs_.io_writeback_14_bits_data_0=0x%0h",this.io_writeback_14_bits_data_0,rhs_.io_writeback_14_bits_data_0),UVM_NONE)
        end

        if(this.io_writeback_14_bits_data_1!=rhs_.io_writeback_14_bits_data_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_bits_data_1=0x%0h while the rhs_.io_writeback_14_bits_data_1=0x%0h",this.io_writeback_14_bits_data_1,rhs_.io_writeback_14_bits_data_1),UVM_NONE)
        end

        if(this.io_writeback_14_bits_data_2!=rhs_.io_writeback_14_bits_data_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_bits_data_2=0x%0h while the rhs_.io_writeback_14_bits_data_2=0x%0h",this.io_writeback_14_bits_data_2,rhs_.io_writeback_14_bits_data_2),UVM_NONE)
        end

        if(this.io_writeback_14_bits_data_3!=rhs_.io_writeback_14_bits_data_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_bits_data_3=0x%0h while the rhs_.io_writeback_14_bits_data_3=0x%0h",this.io_writeback_14_bits_data_3,rhs_.io_writeback_14_bits_data_3),UVM_NONE)
        end

        if(this.io_writeback_14_bits_data_4!=rhs_.io_writeback_14_bits_data_4) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_bits_data_4=0x%0h while the rhs_.io_writeback_14_bits_data_4=0x%0h",this.io_writeback_14_bits_data_4,rhs_.io_writeback_14_bits_data_4),UVM_NONE)
        end

        if(this.io_writeback_14_bits_data_5!=rhs_.io_writeback_14_bits_data_5) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_bits_data_5=0x%0h while the rhs_.io_writeback_14_bits_data_5=0x%0h",this.io_writeback_14_bits_data_5,rhs_.io_writeback_14_bits_data_5),UVM_NONE)
        end

        if(this.io_writeback_14_bits_pdest!=rhs_.io_writeback_14_bits_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_bits_pdest=0x%0h while the rhs_.io_writeback_14_bits_pdest=0x%0h",this.io_writeback_14_bits_pdest,rhs_.io_writeback_14_bits_pdest),UVM_NONE)
        end

        if(this.io_writeback_14_bits_robIdx_flag!=rhs_.io_writeback_14_bits_robIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_bits_robIdx_flag=0x%0h while the rhs_.io_writeback_14_bits_robIdx_flag=0x%0h",this.io_writeback_14_bits_robIdx_flag,rhs_.io_writeback_14_bits_robIdx_flag),UVM_NONE)
        end

        if(this.io_writeback_14_bits_robIdx_value!=rhs_.io_writeback_14_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_bits_robIdx_value=0x%0h while the rhs_.io_writeback_14_bits_robIdx_value=0x%0h",this.io_writeback_14_bits_robIdx_value,rhs_.io_writeback_14_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_writeback_14_bits_intWen!=rhs_.io_writeback_14_bits_intWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_bits_intWen=0x%0h while the rhs_.io_writeback_14_bits_intWen=0x%0h",this.io_writeback_14_bits_intWen,rhs_.io_writeback_14_bits_intWen),UVM_NONE)
        end

        if(this.io_writeback_14_bits_fpWen!=rhs_.io_writeback_14_bits_fpWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_bits_fpWen=0x%0h while the rhs_.io_writeback_14_bits_fpWen=0x%0h",this.io_writeback_14_bits_fpWen,rhs_.io_writeback_14_bits_fpWen),UVM_NONE)
        end

        if(this.io_writeback_14_bits_vecWen!=rhs_.io_writeback_14_bits_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_bits_vecWen=0x%0h while the rhs_.io_writeback_14_bits_vecWen=0x%0h",this.io_writeback_14_bits_vecWen,rhs_.io_writeback_14_bits_vecWen),UVM_NONE)
        end

        if(this.io_writeback_14_bits_v0Wen!=rhs_.io_writeback_14_bits_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_bits_v0Wen=0x%0h while the rhs_.io_writeback_14_bits_v0Wen=0x%0h",this.io_writeback_14_bits_v0Wen,rhs_.io_writeback_14_bits_v0Wen),UVM_NONE)
        end

        if(this.io_writeback_14_bits_vlWen!=rhs_.io_writeback_14_bits_vlWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_bits_vlWen=0x%0h while the rhs_.io_writeback_14_bits_vlWen=0x%0h",this.io_writeback_14_bits_vlWen,rhs_.io_writeback_14_bits_vlWen),UVM_NONE)
        end

        if(this.io_writeback_14_bits_fflags!=rhs_.io_writeback_14_bits_fflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_bits_fflags=0x%0h while the rhs_.io_writeback_14_bits_fflags=0x%0h",this.io_writeback_14_bits_fflags,rhs_.io_writeback_14_bits_fflags),UVM_NONE)
        end

        if(this.io_writeback_14_bits_wflags!=rhs_.io_writeback_14_bits_wflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_bits_wflags=0x%0h while the rhs_.io_writeback_14_bits_wflags=0x%0h",this.io_writeback_14_bits_wflags,rhs_.io_writeback_14_bits_wflags),UVM_NONE)
        end

        if(this.io_writeback_14_bits_exceptionVec_2!=rhs_.io_writeback_14_bits_exceptionVec_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_bits_exceptionVec_2=0x%0h while the rhs_.io_writeback_14_bits_exceptionVec_2=0x%0h",this.io_writeback_14_bits_exceptionVec_2,rhs_.io_writeback_14_bits_exceptionVec_2),UVM_NONE)
        end

        if(this.io_writeback_14_bits_debugInfo_eliminatedMove!=rhs_.io_writeback_14_bits_debugInfo_eliminatedMove) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_bits_debugInfo_eliminatedMove=0x%0h while the rhs_.io_writeback_14_bits_debugInfo_eliminatedMove=0x%0h",this.io_writeback_14_bits_debugInfo_eliminatedMove,rhs_.io_writeback_14_bits_debugInfo_eliminatedMove),UVM_NONE)
        end

        if(this.io_writeback_14_bits_debugInfo_renameTime!=rhs_.io_writeback_14_bits_debugInfo_renameTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_bits_debugInfo_renameTime=0x%0h while the rhs_.io_writeback_14_bits_debugInfo_renameTime=0x%0h",this.io_writeback_14_bits_debugInfo_renameTime,rhs_.io_writeback_14_bits_debugInfo_renameTime),UVM_NONE)
        end

        if(this.io_writeback_14_bits_debugInfo_dispatchTime!=rhs_.io_writeback_14_bits_debugInfo_dispatchTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_bits_debugInfo_dispatchTime=0x%0h while the rhs_.io_writeback_14_bits_debugInfo_dispatchTime=0x%0h",this.io_writeback_14_bits_debugInfo_dispatchTime,rhs_.io_writeback_14_bits_debugInfo_dispatchTime),UVM_NONE)
        end

        if(this.io_writeback_14_bits_debugInfo_enqRsTime!=rhs_.io_writeback_14_bits_debugInfo_enqRsTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_bits_debugInfo_enqRsTime=0x%0h while the rhs_.io_writeback_14_bits_debugInfo_enqRsTime=0x%0h",this.io_writeback_14_bits_debugInfo_enqRsTime,rhs_.io_writeback_14_bits_debugInfo_enqRsTime),UVM_NONE)
        end

        if(this.io_writeback_14_bits_debugInfo_selectTime!=rhs_.io_writeback_14_bits_debugInfo_selectTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_bits_debugInfo_selectTime=0x%0h while the rhs_.io_writeback_14_bits_debugInfo_selectTime=0x%0h",this.io_writeback_14_bits_debugInfo_selectTime,rhs_.io_writeback_14_bits_debugInfo_selectTime),UVM_NONE)
        end

        if(this.io_writeback_14_bits_debugInfo_issueTime!=rhs_.io_writeback_14_bits_debugInfo_issueTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_bits_debugInfo_issueTime=0x%0h while the rhs_.io_writeback_14_bits_debugInfo_issueTime=0x%0h",this.io_writeback_14_bits_debugInfo_issueTime,rhs_.io_writeback_14_bits_debugInfo_issueTime),UVM_NONE)
        end

        if(this.io_writeback_14_bits_debugInfo_writebackTime!=rhs_.io_writeback_14_bits_debugInfo_writebackTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_bits_debugInfo_writebackTime=0x%0h while the rhs_.io_writeback_14_bits_debugInfo_writebackTime=0x%0h",this.io_writeback_14_bits_debugInfo_writebackTime,rhs_.io_writeback_14_bits_debugInfo_writebackTime),UVM_NONE)
        end

        if(this.io_writeback_14_bits_debugInfo_runahead_checkpoint_id!=rhs_.io_writeback_14_bits_debugInfo_runahead_checkpoint_id) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_bits_debugInfo_runahead_checkpoint_id=0x%0h while the rhs_.io_writeback_14_bits_debugInfo_runahead_checkpoint_id=0x%0h",this.io_writeback_14_bits_debugInfo_runahead_checkpoint_id,rhs_.io_writeback_14_bits_debugInfo_runahead_checkpoint_id),UVM_NONE)
        end

        if(this.io_writeback_14_bits_debugInfo_tlbFirstReqTime!=rhs_.io_writeback_14_bits_debugInfo_tlbFirstReqTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_bits_debugInfo_tlbFirstReqTime=0x%0h while the rhs_.io_writeback_14_bits_debugInfo_tlbFirstReqTime=0x%0h",this.io_writeback_14_bits_debugInfo_tlbFirstReqTime,rhs_.io_writeback_14_bits_debugInfo_tlbFirstReqTime),UVM_NONE)
        end

        if(this.io_writeback_14_bits_debugInfo_tlbRespTime!=rhs_.io_writeback_14_bits_debugInfo_tlbRespTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_bits_debugInfo_tlbRespTime=0x%0h while the rhs_.io_writeback_14_bits_debugInfo_tlbRespTime=0x%0h",this.io_writeback_14_bits_debugInfo_tlbRespTime,rhs_.io_writeback_14_bits_debugInfo_tlbRespTime),UVM_NONE)
        end

        if(this.io_writeback_14_bits_debug_seqNum!=rhs_.io_writeback_14_bits_debug_seqNum) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_14_bits_debug_seqNum=0x%0h while the rhs_.io_writeback_14_bits_debug_seqNum=0x%0h",this.io_writeback_14_bits_debug_seqNum,rhs_.io_writeback_14_bits_debug_seqNum),UVM_NONE)
        end

        if(this.io_writeback_13_valid!=rhs_.io_writeback_13_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_13_valid=0x%0h while the rhs_.io_writeback_13_valid=0x%0h",this.io_writeback_13_valid,rhs_.io_writeback_13_valid),UVM_NONE)
        end

        if(this.io_writeback_13_bits_data_0!=rhs_.io_writeback_13_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_13_bits_data_0=0x%0h while the rhs_.io_writeback_13_bits_data_0=0x%0h",this.io_writeback_13_bits_data_0,rhs_.io_writeback_13_bits_data_0),UVM_NONE)
        end

        if(this.io_writeback_13_bits_data_1!=rhs_.io_writeback_13_bits_data_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_13_bits_data_1=0x%0h while the rhs_.io_writeback_13_bits_data_1=0x%0h",this.io_writeback_13_bits_data_1,rhs_.io_writeback_13_bits_data_1),UVM_NONE)
        end

        if(this.io_writeback_13_bits_data_2!=rhs_.io_writeback_13_bits_data_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_13_bits_data_2=0x%0h while the rhs_.io_writeback_13_bits_data_2=0x%0h",this.io_writeback_13_bits_data_2,rhs_.io_writeback_13_bits_data_2),UVM_NONE)
        end

        if(this.io_writeback_13_bits_pdest!=rhs_.io_writeback_13_bits_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_13_bits_pdest=0x%0h while the rhs_.io_writeback_13_bits_pdest=0x%0h",this.io_writeback_13_bits_pdest,rhs_.io_writeback_13_bits_pdest),UVM_NONE)
        end

        if(this.io_writeback_13_bits_robIdx_flag!=rhs_.io_writeback_13_bits_robIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_13_bits_robIdx_flag=0x%0h while the rhs_.io_writeback_13_bits_robIdx_flag=0x%0h",this.io_writeback_13_bits_robIdx_flag,rhs_.io_writeback_13_bits_robIdx_flag),UVM_NONE)
        end

        if(this.io_writeback_13_bits_robIdx_value!=rhs_.io_writeback_13_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_13_bits_robIdx_value=0x%0h while the rhs_.io_writeback_13_bits_robIdx_value=0x%0h",this.io_writeback_13_bits_robIdx_value,rhs_.io_writeback_13_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_writeback_13_bits_vecWen!=rhs_.io_writeback_13_bits_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_13_bits_vecWen=0x%0h while the rhs_.io_writeback_13_bits_vecWen=0x%0h",this.io_writeback_13_bits_vecWen,rhs_.io_writeback_13_bits_vecWen),UVM_NONE)
        end

        if(this.io_writeback_13_bits_v0Wen!=rhs_.io_writeback_13_bits_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_13_bits_v0Wen=0x%0h while the rhs_.io_writeback_13_bits_v0Wen=0x%0h",this.io_writeback_13_bits_v0Wen,rhs_.io_writeback_13_bits_v0Wen),UVM_NONE)
        end

        if(this.io_writeback_13_bits_fflags!=rhs_.io_writeback_13_bits_fflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_13_bits_fflags=0x%0h while the rhs_.io_writeback_13_bits_fflags=0x%0h",this.io_writeback_13_bits_fflags,rhs_.io_writeback_13_bits_fflags),UVM_NONE)
        end

        if(this.io_writeback_13_bits_wflags!=rhs_.io_writeback_13_bits_wflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_13_bits_wflags=0x%0h while the rhs_.io_writeback_13_bits_wflags=0x%0h",this.io_writeback_13_bits_wflags,rhs_.io_writeback_13_bits_wflags),UVM_NONE)
        end

        if(this.io_writeback_13_bits_vxsat!=rhs_.io_writeback_13_bits_vxsat) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_13_bits_vxsat=0x%0h while the rhs_.io_writeback_13_bits_vxsat=0x%0h",this.io_writeback_13_bits_vxsat,rhs_.io_writeback_13_bits_vxsat),UVM_NONE)
        end

        if(this.io_writeback_13_bits_exceptionVec_2!=rhs_.io_writeback_13_bits_exceptionVec_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_13_bits_exceptionVec_2=0x%0h while the rhs_.io_writeback_13_bits_exceptionVec_2=0x%0h",this.io_writeback_13_bits_exceptionVec_2,rhs_.io_writeback_13_bits_exceptionVec_2),UVM_NONE)
        end

        if(this.io_writeback_13_bits_debugInfo_eliminatedMove!=rhs_.io_writeback_13_bits_debugInfo_eliminatedMove) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_13_bits_debugInfo_eliminatedMove=0x%0h while the rhs_.io_writeback_13_bits_debugInfo_eliminatedMove=0x%0h",this.io_writeback_13_bits_debugInfo_eliminatedMove,rhs_.io_writeback_13_bits_debugInfo_eliminatedMove),UVM_NONE)
        end

        if(this.io_writeback_13_bits_debugInfo_renameTime!=rhs_.io_writeback_13_bits_debugInfo_renameTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_13_bits_debugInfo_renameTime=0x%0h while the rhs_.io_writeback_13_bits_debugInfo_renameTime=0x%0h",this.io_writeback_13_bits_debugInfo_renameTime,rhs_.io_writeback_13_bits_debugInfo_renameTime),UVM_NONE)
        end

        if(this.io_writeback_13_bits_debugInfo_dispatchTime!=rhs_.io_writeback_13_bits_debugInfo_dispatchTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_13_bits_debugInfo_dispatchTime=0x%0h while the rhs_.io_writeback_13_bits_debugInfo_dispatchTime=0x%0h",this.io_writeback_13_bits_debugInfo_dispatchTime,rhs_.io_writeback_13_bits_debugInfo_dispatchTime),UVM_NONE)
        end

        if(this.io_writeback_13_bits_debugInfo_enqRsTime!=rhs_.io_writeback_13_bits_debugInfo_enqRsTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_13_bits_debugInfo_enqRsTime=0x%0h while the rhs_.io_writeback_13_bits_debugInfo_enqRsTime=0x%0h",this.io_writeback_13_bits_debugInfo_enqRsTime,rhs_.io_writeback_13_bits_debugInfo_enqRsTime),UVM_NONE)
        end

        if(this.io_writeback_13_bits_debugInfo_selectTime!=rhs_.io_writeback_13_bits_debugInfo_selectTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_13_bits_debugInfo_selectTime=0x%0h while the rhs_.io_writeback_13_bits_debugInfo_selectTime=0x%0h",this.io_writeback_13_bits_debugInfo_selectTime,rhs_.io_writeback_13_bits_debugInfo_selectTime),UVM_NONE)
        end

        if(this.io_writeback_13_bits_debugInfo_issueTime!=rhs_.io_writeback_13_bits_debugInfo_issueTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_13_bits_debugInfo_issueTime=0x%0h while the rhs_.io_writeback_13_bits_debugInfo_issueTime=0x%0h",this.io_writeback_13_bits_debugInfo_issueTime,rhs_.io_writeback_13_bits_debugInfo_issueTime),UVM_NONE)
        end

        if(this.io_writeback_13_bits_debugInfo_writebackTime!=rhs_.io_writeback_13_bits_debugInfo_writebackTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_13_bits_debugInfo_writebackTime=0x%0h while the rhs_.io_writeback_13_bits_debugInfo_writebackTime=0x%0h",this.io_writeback_13_bits_debugInfo_writebackTime,rhs_.io_writeback_13_bits_debugInfo_writebackTime),UVM_NONE)
        end

        if(this.io_writeback_13_bits_debugInfo_runahead_checkpoint_id!=rhs_.io_writeback_13_bits_debugInfo_runahead_checkpoint_id) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_13_bits_debugInfo_runahead_checkpoint_id=0x%0h while the rhs_.io_writeback_13_bits_debugInfo_runahead_checkpoint_id=0x%0h",this.io_writeback_13_bits_debugInfo_runahead_checkpoint_id,rhs_.io_writeback_13_bits_debugInfo_runahead_checkpoint_id),UVM_NONE)
        end

        if(this.io_writeback_13_bits_debugInfo_tlbFirstReqTime!=rhs_.io_writeback_13_bits_debugInfo_tlbFirstReqTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_13_bits_debugInfo_tlbFirstReqTime=0x%0h while the rhs_.io_writeback_13_bits_debugInfo_tlbFirstReqTime=0x%0h",this.io_writeback_13_bits_debugInfo_tlbFirstReqTime,rhs_.io_writeback_13_bits_debugInfo_tlbFirstReqTime),UVM_NONE)
        end

        if(this.io_writeback_13_bits_debugInfo_tlbRespTime!=rhs_.io_writeback_13_bits_debugInfo_tlbRespTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_13_bits_debugInfo_tlbRespTime=0x%0h while the rhs_.io_writeback_13_bits_debugInfo_tlbRespTime=0x%0h",this.io_writeback_13_bits_debugInfo_tlbRespTime,rhs_.io_writeback_13_bits_debugInfo_tlbRespTime),UVM_NONE)
        end

        if(this.io_writeback_13_bits_debug_seqNum!=rhs_.io_writeback_13_bits_debug_seqNum) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_13_bits_debug_seqNum=0x%0h while the rhs_.io_writeback_13_bits_debug_seqNum=0x%0h",this.io_writeback_13_bits_debug_seqNum,rhs_.io_writeback_13_bits_debug_seqNum),UVM_NONE)
        end

        if(this.io_writeback_7_valid!=rhs_.io_writeback_7_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_valid=0x%0h while the rhs_.io_writeback_7_valid=0x%0h",this.io_writeback_7_valid,rhs_.io_writeback_7_valid),UVM_NONE)
        end

        if(this.io_writeback_7_bits_data_0!=rhs_.io_writeback_7_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_data_0=0x%0h while the rhs_.io_writeback_7_bits_data_0=0x%0h",this.io_writeback_7_bits_data_0,rhs_.io_writeback_7_bits_data_0),UVM_NONE)
        end

        if(this.io_writeback_7_bits_data_1!=rhs_.io_writeback_7_bits_data_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_data_1=0x%0h while the rhs_.io_writeback_7_bits_data_1=0x%0h",this.io_writeback_7_bits_data_1,rhs_.io_writeback_7_bits_data_1),UVM_NONE)
        end

        if(this.io_writeback_7_bits_pdest!=rhs_.io_writeback_7_bits_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_pdest=0x%0h while the rhs_.io_writeback_7_bits_pdest=0x%0h",this.io_writeback_7_bits_pdest,rhs_.io_writeback_7_bits_pdest),UVM_NONE)
        end

        if(this.io_writeback_7_bits_robIdx_flag!=rhs_.io_writeback_7_bits_robIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_robIdx_flag=0x%0h while the rhs_.io_writeback_7_bits_robIdx_flag=0x%0h",this.io_writeback_7_bits_robIdx_flag,rhs_.io_writeback_7_bits_robIdx_flag),UVM_NONE)
        end

        if(this.io_writeback_7_bits_robIdx_value!=rhs_.io_writeback_7_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_robIdx_value=0x%0h while the rhs_.io_writeback_7_bits_robIdx_value=0x%0h",this.io_writeback_7_bits_robIdx_value,rhs_.io_writeback_7_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_writeback_7_bits_intWen!=rhs_.io_writeback_7_bits_intWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_intWen=0x%0h while the rhs_.io_writeback_7_bits_intWen=0x%0h",this.io_writeback_7_bits_intWen,rhs_.io_writeback_7_bits_intWen),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_valid!=rhs_.io_writeback_7_bits_redirect_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_valid=0x%0h while the rhs_.io_writeback_7_bits_redirect_valid=0x%0h",this.io_writeback_7_bits_redirect_valid,rhs_.io_writeback_7_bits_redirect_valid),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_isRVC!=rhs_.io_writeback_7_bits_redirect_bits_isRVC) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_isRVC=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_isRVC=0x%0h",this.io_writeback_7_bits_redirect_bits_isRVC,rhs_.io_writeback_7_bits_redirect_bits_isRVC),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_robIdx_flag!=rhs_.io_writeback_7_bits_redirect_bits_robIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_robIdx_flag=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_robIdx_flag=0x%0h",this.io_writeback_7_bits_redirect_bits_robIdx_flag,rhs_.io_writeback_7_bits_redirect_bits_robIdx_flag),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_robIdx_value!=rhs_.io_writeback_7_bits_redirect_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_robIdx_value=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_robIdx_value=0x%0h",this.io_writeback_7_bits_redirect_bits_robIdx_value,rhs_.io_writeback_7_bits_redirect_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_ftqIdx_flag!=rhs_.io_writeback_7_bits_redirect_bits_ftqIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_ftqIdx_flag=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_ftqIdx_flag=0x%0h",this.io_writeback_7_bits_redirect_bits_ftqIdx_flag,rhs_.io_writeback_7_bits_redirect_bits_ftqIdx_flag),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_ftqIdx_value!=rhs_.io_writeback_7_bits_redirect_bits_ftqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_ftqIdx_value=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_ftqIdx_value=0x%0h",this.io_writeback_7_bits_redirect_bits_ftqIdx_value,rhs_.io_writeback_7_bits_redirect_bits_ftqIdx_value),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_ftqOffset!=rhs_.io_writeback_7_bits_redirect_bits_ftqOffset) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_ftqOffset=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_ftqOffset=0x%0h",this.io_writeback_7_bits_redirect_bits_ftqOffset,rhs_.io_writeback_7_bits_redirect_bits_ftqOffset),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_level!=rhs_.io_writeback_7_bits_redirect_bits_level) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_level=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_level=0x%0h",this.io_writeback_7_bits_redirect_bits_level,rhs_.io_writeback_7_bits_redirect_bits_level),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_interrupt!=rhs_.io_writeback_7_bits_redirect_bits_interrupt) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_interrupt=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_interrupt=0x%0h",this.io_writeback_7_bits_redirect_bits_interrupt,rhs_.io_writeback_7_bits_redirect_bits_interrupt),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_pc!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_pc) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_pc=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_pc=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_pc,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_pc),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_ssp!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_ssp) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_ssp=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_ssp=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_ssp,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_ssp),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_sctr!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_sctr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_sctr=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_sctr=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_sctr,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_sctr),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_ghr!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_ghr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_ghr=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_ghr=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_ghr,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_ghr),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_target!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_target) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_target=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_target=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_target,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_target),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_taken!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_taken) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_taken=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_taken=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_taken,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_taken),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_shift!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_shift) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_shift=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_shift=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_shift,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_shift),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF!=rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF=0x%0h",this.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF,rhs_.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_fullTarget!=rhs_.io_writeback_7_bits_redirect_bits_fullTarget) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_fullTarget=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_fullTarget=0x%0h",this.io_writeback_7_bits_redirect_bits_fullTarget,rhs_.io_writeback_7_bits_redirect_bits_fullTarget),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_stFtqIdx_flag!=rhs_.io_writeback_7_bits_redirect_bits_stFtqIdx_flag) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_stFtqIdx_flag=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_stFtqIdx_flag=0x%0h",this.io_writeback_7_bits_redirect_bits_stFtqIdx_flag,rhs_.io_writeback_7_bits_redirect_bits_stFtqIdx_flag),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_stFtqIdx_value!=rhs_.io_writeback_7_bits_redirect_bits_stFtqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_stFtqIdx_value=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_stFtqIdx_value=0x%0h",this.io_writeback_7_bits_redirect_bits_stFtqIdx_value,rhs_.io_writeback_7_bits_redirect_bits_stFtqIdx_value),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_stFtqOffset!=rhs_.io_writeback_7_bits_redirect_bits_stFtqOffset) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_stFtqOffset=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_stFtqOffset=0x%0h",this.io_writeback_7_bits_redirect_bits_stFtqOffset,rhs_.io_writeback_7_bits_redirect_bits_stFtqOffset),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id!=rhs_.io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id=0x%0h",this.io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id,rhs_.io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_debugIsCtrl!=rhs_.io_writeback_7_bits_redirect_bits_debugIsCtrl) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_debugIsCtrl=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_debugIsCtrl=0x%0h",this.io_writeback_7_bits_redirect_bits_debugIsCtrl,rhs_.io_writeback_7_bits_redirect_bits_debugIsCtrl),UVM_NONE)
        end

        if(this.io_writeback_7_bits_redirect_bits_debugIsMemVio!=rhs_.io_writeback_7_bits_redirect_bits_debugIsMemVio) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_redirect_bits_debugIsMemVio=0x%0h while the rhs_.io_writeback_7_bits_redirect_bits_debugIsMemVio=0x%0h",this.io_writeback_7_bits_redirect_bits_debugIsMemVio,rhs_.io_writeback_7_bits_redirect_bits_debugIsMemVio),UVM_NONE)
        end

        if(this.io_writeback_7_bits_exceptionVec_2!=rhs_.io_writeback_7_bits_exceptionVec_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_exceptionVec_2=0x%0h while the rhs_.io_writeback_7_bits_exceptionVec_2=0x%0h",this.io_writeback_7_bits_exceptionVec_2,rhs_.io_writeback_7_bits_exceptionVec_2),UVM_NONE)
        end

        if(this.io_writeback_7_bits_exceptionVec_3!=rhs_.io_writeback_7_bits_exceptionVec_3) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_exceptionVec_3=0x%0h while the rhs_.io_writeback_7_bits_exceptionVec_3=0x%0h",this.io_writeback_7_bits_exceptionVec_3,rhs_.io_writeback_7_bits_exceptionVec_3),UVM_NONE)
        end

        if(this.io_writeback_7_bits_exceptionVec_8!=rhs_.io_writeback_7_bits_exceptionVec_8) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_exceptionVec_8=0x%0h while the rhs_.io_writeback_7_bits_exceptionVec_8=0x%0h",this.io_writeback_7_bits_exceptionVec_8,rhs_.io_writeback_7_bits_exceptionVec_8),UVM_NONE)
        end

        if(this.io_writeback_7_bits_exceptionVec_9!=rhs_.io_writeback_7_bits_exceptionVec_9) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_exceptionVec_9=0x%0h while the rhs_.io_writeback_7_bits_exceptionVec_9=0x%0h",this.io_writeback_7_bits_exceptionVec_9,rhs_.io_writeback_7_bits_exceptionVec_9),UVM_NONE)
        end

        if(this.io_writeback_7_bits_exceptionVec_10!=rhs_.io_writeback_7_bits_exceptionVec_10) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_exceptionVec_10=0x%0h while the rhs_.io_writeback_7_bits_exceptionVec_10=0x%0h",this.io_writeback_7_bits_exceptionVec_10,rhs_.io_writeback_7_bits_exceptionVec_10),UVM_NONE)
        end

        if(this.io_writeback_7_bits_exceptionVec_11!=rhs_.io_writeback_7_bits_exceptionVec_11) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_exceptionVec_11=0x%0h while the rhs_.io_writeback_7_bits_exceptionVec_11=0x%0h",this.io_writeback_7_bits_exceptionVec_11,rhs_.io_writeback_7_bits_exceptionVec_11),UVM_NONE)
        end

        if(this.io_writeback_7_bits_exceptionVec_22!=rhs_.io_writeback_7_bits_exceptionVec_22) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_exceptionVec_22=0x%0h while the rhs_.io_writeback_7_bits_exceptionVec_22=0x%0h",this.io_writeback_7_bits_exceptionVec_22,rhs_.io_writeback_7_bits_exceptionVec_22),UVM_NONE)
        end

        if(this.io_writeback_7_bits_flushPipe!=rhs_.io_writeback_7_bits_flushPipe) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_flushPipe=0x%0h while the rhs_.io_writeback_7_bits_flushPipe=0x%0h",this.io_writeback_7_bits_flushPipe,rhs_.io_writeback_7_bits_flushPipe),UVM_NONE)
        end

        if(this.io_writeback_7_bits_predecodeInfo_valid!=rhs_.io_writeback_7_bits_predecodeInfo_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_predecodeInfo_valid=0x%0h while the rhs_.io_writeback_7_bits_predecodeInfo_valid=0x%0h",this.io_writeback_7_bits_predecodeInfo_valid,rhs_.io_writeback_7_bits_predecodeInfo_valid),UVM_NONE)
        end

        if(this.io_writeback_7_bits_predecodeInfo_isRVC!=rhs_.io_writeback_7_bits_predecodeInfo_isRVC) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_predecodeInfo_isRVC=0x%0h while the rhs_.io_writeback_7_bits_predecodeInfo_isRVC=0x%0h",this.io_writeback_7_bits_predecodeInfo_isRVC,rhs_.io_writeback_7_bits_predecodeInfo_isRVC),UVM_NONE)
        end

        if(this.io_writeback_7_bits_predecodeInfo_brType!=rhs_.io_writeback_7_bits_predecodeInfo_brType) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_predecodeInfo_brType=0x%0h while the rhs_.io_writeback_7_bits_predecodeInfo_brType=0x%0h",this.io_writeback_7_bits_predecodeInfo_brType,rhs_.io_writeback_7_bits_predecodeInfo_brType),UVM_NONE)
        end

        if(this.io_writeback_7_bits_predecodeInfo_isCall!=rhs_.io_writeback_7_bits_predecodeInfo_isCall) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_predecodeInfo_isCall=0x%0h while the rhs_.io_writeback_7_bits_predecodeInfo_isCall=0x%0h",this.io_writeback_7_bits_predecodeInfo_isCall,rhs_.io_writeback_7_bits_predecodeInfo_isCall),UVM_NONE)
        end

        if(this.io_writeback_7_bits_predecodeInfo_isRet!=rhs_.io_writeback_7_bits_predecodeInfo_isRet) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_predecodeInfo_isRet=0x%0h while the rhs_.io_writeback_7_bits_predecodeInfo_isRet=0x%0h",this.io_writeback_7_bits_predecodeInfo_isRet,rhs_.io_writeback_7_bits_predecodeInfo_isRet),UVM_NONE)
        end

        if(this.io_writeback_7_bits_debug_isPerfCnt!=rhs_.io_writeback_7_bits_debug_isPerfCnt) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_debug_isPerfCnt=0x%0h while the rhs_.io_writeback_7_bits_debug_isPerfCnt=0x%0h",this.io_writeback_7_bits_debug_isPerfCnt,rhs_.io_writeback_7_bits_debug_isPerfCnt),UVM_NONE)
        end

        if(this.io_writeback_7_bits_debugInfo_eliminatedMove!=rhs_.io_writeback_7_bits_debugInfo_eliminatedMove) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_debugInfo_eliminatedMove=0x%0h while the rhs_.io_writeback_7_bits_debugInfo_eliminatedMove=0x%0h",this.io_writeback_7_bits_debugInfo_eliminatedMove,rhs_.io_writeback_7_bits_debugInfo_eliminatedMove),UVM_NONE)
        end

        if(this.io_writeback_7_bits_debugInfo_renameTime!=rhs_.io_writeback_7_bits_debugInfo_renameTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_debugInfo_renameTime=0x%0h while the rhs_.io_writeback_7_bits_debugInfo_renameTime=0x%0h",this.io_writeback_7_bits_debugInfo_renameTime,rhs_.io_writeback_7_bits_debugInfo_renameTime),UVM_NONE)
        end

        if(this.io_writeback_7_bits_debugInfo_dispatchTime!=rhs_.io_writeback_7_bits_debugInfo_dispatchTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_debugInfo_dispatchTime=0x%0h while the rhs_.io_writeback_7_bits_debugInfo_dispatchTime=0x%0h",this.io_writeback_7_bits_debugInfo_dispatchTime,rhs_.io_writeback_7_bits_debugInfo_dispatchTime),UVM_NONE)
        end

        if(this.io_writeback_7_bits_debugInfo_enqRsTime!=rhs_.io_writeback_7_bits_debugInfo_enqRsTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_debugInfo_enqRsTime=0x%0h while the rhs_.io_writeback_7_bits_debugInfo_enqRsTime=0x%0h",this.io_writeback_7_bits_debugInfo_enqRsTime,rhs_.io_writeback_7_bits_debugInfo_enqRsTime),UVM_NONE)
        end

        if(this.io_writeback_7_bits_debugInfo_selectTime!=rhs_.io_writeback_7_bits_debugInfo_selectTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_debugInfo_selectTime=0x%0h while the rhs_.io_writeback_7_bits_debugInfo_selectTime=0x%0h",this.io_writeback_7_bits_debugInfo_selectTime,rhs_.io_writeback_7_bits_debugInfo_selectTime),UVM_NONE)
        end

        if(this.io_writeback_7_bits_debugInfo_issueTime!=rhs_.io_writeback_7_bits_debugInfo_issueTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_debugInfo_issueTime=0x%0h while the rhs_.io_writeback_7_bits_debugInfo_issueTime=0x%0h",this.io_writeback_7_bits_debugInfo_issueTime,rhs_.io_writeback_7_bits_debugInfo_issueTime),UVM_NONE)
        end

        if(this.io_writeback_7_bits_debugInfo_writebackTime!=rhs_.io_writeback_7_bits_debugInfo_writebackTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_debugInfo_writebackTime=0x%0h while the rhs_.io_writeback_7_bits_debugInfo_writebackTime=0x%0h",this.io_writeback_7_bits_debugInfo_writebackTime,rhs_.io_writeback_7_bits_debugInfo_writebackTime),UVM_NONE)
        end

        if(this.io_writeback_7_bits_debugInfo_runahead_checkpoint_id!=rhs_.io_writeback_7_bits_debugInfo_runahead_checkpoint_id) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_debugInfo_runahead_checkpoint_id=0x%0h while the rhs_.io_writeback_7_bits_debugInfo_runahead_checkpoint_id=0x%0h",this.io_writeback_7_bits_debugInfo_runahead_checkpoint_id,rhs_.io_writeback_7_bits_debugInfo_runahead_checkpoint_id),UVM_NONE)
        end

        if(this.io_writeback_7_bits_debugInfo_tlbFirstReqTime!=rhs_.io_writeback_7_bits_debugInfo_tlbFirstReqTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_debugInfo_tlbFirstReqTime=0x%0h while the rhs_.io_writeback_7_bits_debugInfo_tlbFirstReqTime=0x%0h",this.io_writeback_7_bits_debugInfo_tlbFirstReqTime,rhs_.io_writeback_7_bits_debugInfo_tlbFirstReqTime),UVM_NONE)
        end

        if(this.io_writeback_7_bits_debugInfo_tlbRespTime!=rhs_.io_writeback_7_bits_debugInfo_tlbRespTime) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_debugInfo_tlbRespTime=0x%0h while the rhs_.io_writeback_7_bits_debugInfo_tlbRespTime=0x%0h",this.io_writeback_7_bits_debugInfo_tlbRespTime,rhs_.io_writeback_7_bits_debugInfo_tlbRespTime),UVM_NONE)
        end

        if(this.io_writeback_7_bits_debug_seqNum!=rhs_.io_writeback_7_bits_debug_seqNum) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_7_bits_debug_seqNum=0x%0h while the rhs_.io_writeback_7_bits_debug_seqNum=0x%0h",this.io_writeback_7_bits_debug_seqNum,rhs_.io_writeback_7_bits_debug_seqNum),UVM_NONE)
        end

        if(this.io_writeback_5_valid!=rhs_.io_writeback_5_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_5_valid=0x%0h while the rhs_.io_writeback_5_valid=0x%0h",this.io_writeback_5_valid,rhs_.io_writeback_5_valid),UVM_NONE)
        end

        if(this.io_writeback_5_bits_redirect_valid!=rhs_.io_writeback_5_bits_redirect_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_5_bits_redirect_valid=0x%0h while the rhs_.io_writeback_5_bits_redirect_valid=0x%0h",this.io_writeback_5_bits_redirect_valid,rhs_.io_writeback_5_bits_redirect_valid),UVM_NONE)
        end

        if(this.io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred!=rhs_.io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred=0x%0h while the rhs_.io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred=0x%0h",this.io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred,rhs_.io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred),UVM_NONE)
        end

        if(this.io_writeback_3_valid!=rhs_.io_writeback_3_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_3_valid=0x%0h while the rhs_.io_writeback_3_valid=0x%0h",this.io_writeback_3_valid,rhs_.io_writeback_3_valid),UVM_NONE)
        end

        if(this.io_writeback_3_bits_redirect_valid!=rhs_.io_writeback_3_bits_redirect_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_3_bits_redirect_valid=0x%0h while the rhs_.io_writeback_3_bits_redirect_valid=0x%0h",this.io_writeback_3_bits_redirect_valid,rhs_.io_writeback_3_bits_redirect_valid),UVM_NONE)
        end

        if(this.io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred!=rhs_.io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred=0x%0h while the rhs_.io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred=0x%0h",this.io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred,rhs_.io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred),UVM_NONE)
        end

        if(this.io_writeback_1_valid!=rhs_.io_writeback_1_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_1_valid=0x%0h while the rhs_.io_writeback_1_valid=0x%0h",this.io_writeback_1_valid,rhs_.io_writeback_1_valid),UVM_NONE)
        end

        if(this.io_writeback_1_bits_redirect_valid!=rhs_.io_writeback_1_bits_redirect_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_1_bits_redirect_valid=0x%0h while the rhs_.io_writeback_1_bits_redirect_valid=0x%0h",this.io_writeback_1_bits_redirect_valid,rhs_.io_writeback_1_bits_redirect_valid),UVM_NONE)
        end

        if(this.io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred!=rhs_.io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred=0x%0h while the rhs_.io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred=0x%0h",this.io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred,rhs_.io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred),UVM_NONE)
        end

        if(this.io_exuWriteback_26_valid!=rhs_.io_exuWriteback_26_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_26_valid=0x%0h while the rhs_.io_exuWriteback_26_valid=0x%0h",this.io_exuWriteback_26_valid,rhs_.io_exuWriteback_26_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_26_bits_robIdx_value!=rhs_.io_exuWriteback_26_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_26_bits_robIdx_value=0x%0h while the rhs_.io_exuWriteback_26_bits_robIdx_value=0x%0h",this.io_exuWriteback_26_bits_robIdx_value,rhs_.io_exuWriteback_26_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_25_valid!=rhs_.io_exuWriteback_25_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_25_valid=0x%0h while the rhs_.io_exuWriteback_25_valid=0x%0h",this.io_exuWriteback_25_valid,rhs_.io_exuWriteback_25_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_25_bits_robIdx_value!=rhs_.io_exuWriteback_25_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_25_bits_robIdx_value=0x%0h while the rhs_.io_exuWriteback_25_bits_robIdx_value=0x%0h",this.io_exuWriteback_25_bits_robIdx_value,rhs_.io_exuWriteback_25_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_24_valid!=rhs_.io_exuWriteback_24_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_24_valid=0x%0h while the rhs_.io_exuWriteback_24_valid=0x%0h",this.io_exuWriteback_24_valid,rhs_.io_exuWriteback_24_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_24_bits_data_0!=rhs_.io_exuWriteback_24_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_24_bits_data_0=0x%0h while the rhs_.io_exuWriteback_24_bits_data_0=0x%0h",this.io_exuWriteback_24_bits_data_0,rhs_.io_exuWriteback_24_bits_data_0),UVM_NONE)
        end

        if(this.io_exuWriteback_24_bits_pdest!=rhs_.io_exuWriteback_24_bits_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_24_bits_pdest=0x%0h while the rhs_.io_exuWriteback_24_bits_pdest=0x%0h",this.io_exuWriteback_24_bits_pdest,rhs_.io_exuWriteback_24_bits_pdest),UVM_NONE)
        end

        if(this.io_exuWriteback_24_bits_robIdx_value!=rhs_.io_exuWriteback_24_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_24_bits_robIdx_value=0x%0h while the rhs_.io_exuWriteback_24_bits_robIdx_value=0x%0h",this.io_exuWriteback_24_bits_robIdx_value,rhs_.io_exuWriteback_24_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_24_bits_vecWen!=rhs_.io_exuWriteback_24_bits_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_24_bits_vecWen=0x%0h while the rhs_.io_exuWriteback_24_bits_vecWen=0x%0h",this.io_exuWriteback_24_bits_vecWen,rhs_.io_exuWriteback_24_bits_vecWen),UVM_NONE)
        end

        if(this.io_exuWriteback_24_bits_v0Wen!=rhs_.io_exuWriteback_24_bits_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_24_bits_v0Wen=0x%0h while the rhs_.io_exuWriteback_24_bits_v0Wen=0x%0h",this.io_exuWriteback_24_bits_v0Wen,rhs_.io_exuWriteback_24_bits_v0Wen),UVM_NONE)
        end

        if(this.io_exuWriteback_24_bits_vls_vdIdx!=rhs_.io_exuWriteback_24_bits_vls_vdIdx) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_24_bits_vls_vdIdx=0x%0h while the rhs_.io_exuWriteback_24_bits_vls_vdIdx=0x%0h",this.io_exuWriteback_24_bits_vls_vdIdx,rhs_.io_exuWriteback_24_bits_vls_vdIdx),UVM_NONE)
        end

        if(this.io_exuWriteback_24_bits_debug_isMMIO!=rhs_.io_exuWriteback_24_bits_debug_isMMIO) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_24_bits_debug_isMMIO=0x%0h while the rhs_.io_exuWriteback_24_bits_debug_isMMIO=0x%0h",this.io_exuWriteback_24_bits_debug_isMMIO,rhs_.io_exuWriteback_24_bits_debug_isMMIO),UVM_NONE)
        end

        if(this.io_exuWriteback_24_bits_debug_isNCIO!=rhs_.io_exuWriteback_24_bits_debug_isNCIO) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_24_bits_debug_isNCIO=0x%0h while the rhs_.io_exuWriteback_24_bits_debug_isNCIO=0x%0h",this.io_exuWriteback_24_bits_debug_isNCIO,rhs_.io_exuWriteback_24_bits_debug_isNCIO),UVM_NONE)
        end

        if(this.io_exuWriteback_24_bits_debug_isPerfCnt!=rhs_.io_exuWriteback_24_bits_debug_isPerfCnt) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_24_bits_debug_isPerfCnt=0x%0h while the rhs_.io_exuWriteback_24_bits_debug_isPerfCnt=0x%0h",this.io_exuWriteback_24_bits_debug_isPerfCnt,rhs_.io_exuWriteback_24_bits_debug_isPerfCnt),UVM_NONE)
        end

        if(this.io_exuWriteback_24_bits_debug_paddr!=rhs_.io_exuWriteback_24_bits_debug_paddr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_24_bits_debug_paddr=0x%0h while the rhs_.io_exuWriteback_24_bits_debug_paddr=0x%0h",this.io_exuWriteback_24_bits_debug_paddr,rhs_.io_exuWriteback_24_bits_debug_paddr),UVM_NONE)
        end

        if(this.io_exuWriteback_23_valid!=rhs_.io_exuWriteback_23_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_23_valid=0x%0h while the rhs_.io_exuWriteback_23_valid=0x%0h",this.io_exuWriteback_23_valid,rhs_.io_exuWriteback_23_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_23_bits_data_0!=rhs_.io_exuWriteback_23_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_23_bits_data_0=0x%0h while the rhs_.io_exuWriteback_23_bits_data_0=0x%0h",this.io_exuWriteback_23_bits_data_0,rhs_.io_exuWriteback_23_bits_data_0),UVM_NONE)
        end

        if(this.io_exuWriteback_23_bits_pdest!=rhs_.io_exuWriteback_23_bits_pdest) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_23_bits_pdest=0x%0h while the rhs_.io_exuWriteback_23_bits_pdest=0x%0h",this.io_exuWriteback_23_bits_pdest,rhs_.io_exuWriteback_23_bits_pdest),UVM_NONE)
        end

        if(this.io_exuWriteback_23_bits_robIdx_value!=rhs_.io_exuWriteback_23_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_23_bits_robIdx_value=0x%0h while the rhs_.io_exuWriteback_23_bits_robIdx_value=0x%0h",this.io_exuWriteback_23_bits_robIdx_value,rhs_.io_exuWriteback_23_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_23_bits_vecWen!=rhs_.io_exuWriteback_23_bits_vecWen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_23_bits_vecWen=0x%0h while the rhs_.io_exuWriteback_23_bits_vecWen=0x%0h",this.io_exuWriteback_23_bits_vecWen,rhs_.io_exuWriteback_23_bits_vecWen),UVM_NONE)
        end

        if(this.io_exuWriteback_23_bits_v0Wen!=rhs_.io_exuWriteback_23_bits_v0Wen) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_23_bits_v0Wen=0x%0h while the rhs_.io_exuWriteback_23_bits_v0Wen=0x%0h",this.io_exuWriteback_23_bits_v0Wen,rhs_.io_exuWriteback_23_bits_v0Wen),UVM_NONE)
        end

        if(this.io_exuWriteback_23_bits_vls_vdIdx!=rhs_.io_exuWriteback_23_bits_vls_vdIdx) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_23_bits_vls_vdIdx=0x%0h while the rhs_.io_exuWriteback_23_bits_vls_vdIdx=0x%0h",this.io_exuWriteback_23_bits_vls_vdIdx,rhs_.io_exuWriteback_23_bits_vls_vdIdx),UVM_NONE)
        end

        if(this.io_exuWriteback_23_bits_debug_isMMIO!=rhs_.io_exuWriteback_23_bits_debug_isMMIO) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_23_bits_debug_isMMIO=0x%0h while the rhs_.io_exuWriteback_23_bits_debug_isMMIO=0x%0h",this.io_exuWriteback_23_bits_debug_isMMIO,rhs_.io_exuWriteback_23_bits_debug_isMMIO),UVM_NONE)
        end

        if(this.io_exuWriteback_23_bits_debug_isNCIO!=rhs_.io_exuWriteback_23_bits_debug_isNCIO) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_23_bits_debug_isNCIO=0x%0h while the rhs_.io_exuWriteback_23_bits_debug_isNCIO=0x%0h",this.io_exuWriteback_23_bits_debug_isNCIO,rhs_.io_exuWriteback_23_bits_debug_isNCIO),UVM_NONE)
        end

        if(this.io_exuWriteback_23_bits_debug_isPerfCnt!=rhs_.io_exuWriteback_23_bits_debug_isPerfCnt) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_23_bits_debug_isPerfCnt=0x%0h while the rhs_.io_exuWriteback_23_bits_debug_isPerfCnt=0x%0h",this.io_exuWriteback_23_bits_debug_isPerfCnt,rhs_.io_exuWriteback_23_bits_debug_isPerfCnt),UVM_NONE)
        end

        if(this.io_exuWriteback_23_bits_debug_paddr!=rhs_.io_exuWriteback_23_bits_debug_paddr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_23_bits_debug_paddr=0x%0h while the rhs_.io_exuWriteback_23_bits_debug_paddr=0x%0h",this.io_exuWriteback_23_bits_debug_paddr,rhs_.io_exuWriteback_23_bits_debug_paddr),UVM_NONE)
        end

        if(this.io_exuWriteback_22_valid!=rhs_.io_exuWriteback_22_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_22_valid=0x%0h while the rhs_.io_exuWriteback_22_valid=0x%0h",this.io_exuWriteback_22_valid,rhs_.io_exuWriteback_22_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_22_bits_data_0!=rhs_.io_exuWriteback_22_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_22_bits_data_0=0x%0h while the rhs_.io_exuWriteback_22_bits_data_0=0x%0h",this.io_exuWriteback_22_bits_data_0,rhs_.io_exuWriteback_22_bits_data_0),UVM_NONE)
        end

        if(this.io_exuWriteback_22_bits_robIdx_value!=rhs_.io_exuWriteback_22_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_22_bits_robIdx_value=0x%0h while the rhs_.io_exuWriteback_22_bits_robIdx_value=0x%0h",this.io_exuWriteback_22_bits_robIdx_value,rhs_.io_exuWriteback_22_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_22_bits_lqIdx_value!=rhs_.io_exuWriteback_22_bits_lqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_22_bits_lqIdx_value=0x%0h while the rhs_.io_exuWriteback_22_bits_lqIdx_value=0x%0h",this.io_exuWriteback_22_bits_lqIdx_value,rhs_.io_exuWriteback_22_bits_lqIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_22_bits_debug_isMMIO!=rhs_.io_exuWriteback_22_bits_debug_isMMIO) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_22_bits_debug_isMMIO=0x%0h while the rhs_.io_exuWriteback_22_bits_debug_isMMIO=0x%0h",this.io_exuWriteback_22_bits_debug_isMMIO,rhs_.io_exuWriteback_22_bits_debug_isMMIO),UVM_NONE)
        end

        if(this.io_exuWriteback_22_bits_debug_isNCIO!=rhs_.io_exuWriteback_22_bits_debug_isNCIO) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_22_bits_debug_isNCIO=0x%0h while the rhs_.io_exuWriteback_22_bits_debug_isNCIO=0x%0h",this.io_exuWriteback_22_bits_debug_isNCIO,rhs_.io_exuWriteback_22_bits_debug_isNCIO),UVM_NONE)
        end

        if(this.io_exuWriteback_22_bits_debug_isPerfCnt!=rhs_.io_exuWriteback_22_bits_debug_isPerfCnt) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_22_bits_debug_isPerfCnt=0x%0h while the rhs_.io_exuWriteback_22_bits_debug_isPerfCnt=0x%0h",this.io_exuWriteback_22_bits_debug_isPerfCnt,rhs_.io_exuWriteback_22_bits_debug_isPerfCnt),UVM_NONE)
        end

        if(this.io_exuWriteback_22_bits_debug_paddr!=rhs_.io_exuWriteback_22_bits_debug_paddr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_22_bits_debug_paddr=0x%0h while the rhs_.io_exuWriteback_22_bits_debug_paddr=0x%0h",this.io_exuWriteback_22_bits_debug_paddr,rhs_.io_exuWriteback_22_bits_debug_paddr),UVM_NONE)
        end

        if(this.io_exuWriteback_21_valid!=rhs_.io_exuWriteback_21_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_21_valid=0x%0h while the rhs_.io_exuWriteback_21_valid=0x%0h",this.io_exuWriteback_21_valid,rhs_.io_exuWriteback_21_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_21_bits_data_0!=rhs_.io_exuWriteback_21_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_21_bits_data_0=0x%0h while the rhs_.io_exuWriteback_21_bits_data_0=0x%0h",this.io_exuWriteback_21_bits_data_0,rhs_.io_exuWriteback_21_bits_data_0),UVM_NONE)
        end

        if(this.io_exuWriteback_21_bits_robIdx_value!=rhs_.io_exuWriteback_21_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_21_bits_robIdx_value=0x%0h while the rhs_.io_exuWriteback_21_bits_robIdx_value=0x%0h",this.io_exuWriteback_21_bits_robIdx_value,rhs_.io_exuWriteback_21_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_21_bits_lqIdx_value!=rhs_.io_exuWriteback_21_bits_lqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_21_bits_lqIdx_value=0x%0h while the rhs_.io_exuWriteback_21_bits_lqIdx_value=0x%0h",this.io_exuWriteback_21_bits_lqIdx_value,rhs_.io_exuWriteback_21_bits_lqIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_21_bits_debug_isMMIO!=rhs_.io_exuWriteback_21_bits_debug_isMMIO) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_21_bits_debug_isMMIO=0x%0h while the rhs_.io_exuWriteback_21_bits_debug_isMMIO=0x%0h",this.io_exuWriteback_21_bits_debug_isMMIO,rhs_.io_exuWriteback_21_bits_debug_isMMIO),UVM_NONE)
        end

        if(this.io_exuWriteback_21_bits_debug_isNCIO!=rhs_.io_exuWriteback_21_bits_debug_isNCIO) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_21_bits_debug_isNCIO=0x%0h while the rhs_.io_exuWriteback_21_bits_debug_isNCIO=0x%0h",this.io_exuWriteback_21_bits_debug_isNCIO,rhs_.io_exuWriteback_21_bits_debug_isNCIO),UVM_NONE)
        end

        if(this.io_exuWriteback_21_bits_debug_isPerfCnt!=rhs_.io_exuWriteback_21_bits_debug_isPerfCnt) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_21_bits_debug_isPerfCnt=0x%0h while the rhs_.io_exuWriteback_21_bits_debug_isPerfCnt=0x%0h",this.io_exuWriteback_21_bits_debug_isPerfCnt,rhs_.io_exuWriteback_21_bits_debug_isPerfCnt),UVM_NONE)
        end

        if(this.io_exuWriteback_21_bits_debug_paddr!=rhs_.io_exuWriteback_21_bits_debug_paddr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_21_bits_debug_paddr=0x%0h while the rhs_.io_exuWriteback_21_bits_debug_paddr=0x%0h",this.io_exuWriteback_21_bits_debug_paddr,rhs_.io_exuWriteback_21_bits_debug_paddr),UVM_NONE)
        end

        if(this.io_exuWriteback_20_valid!=rhs_.io_exuWriteback_20_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_20_valid=0x%0h while the rhs_.io_exuWriteback_20_valid=0x%0h",this.io_exuWriteback_20_valid,rhs_.io_exuWriteback_20_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_20_bits_data_0!=rhs_.io_exuWriteback_20_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_20_bits_data_0=0x%0h while the rhs_.io_exuWriteback_20_bits_data_0=0x%0h",this.io_exuWriteback_20_bits_data_0,rhs_.io_exuWriteback_20_bits_data_0),UVM_NONE)
        end

        if(this.io_exuWriteback_20_bits_robIdx_value!=rhs_.io_exuWriteback_20_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_20_bits_robIdx_value=0x%0h while the rhs_.io_exuWriteback_20_bits_robIdx_value=0x%0h",this.io_exuWriteback_20_bits_robIdx_value,rhs_.io_exuWriteback_20_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_20_bits_lqIdx_value!=rhs_.io_exuWriteback_20_bits_lqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_20_bits_lqIdx_value=0x%0h while the rhs_.io_exuWriteback_20_bits_lqIdx_value=0x%0h",this.io_exuWriteback_20_bits_lqIdx_value,rhs_.io_exuWriteback_20_bits_lqIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_20_bits_debug_isMMIO!=rhs_.io_exuWriteback_20_bits_debug_isMMIO) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_20_bits_debug_isMMIO=0x%0h while the rhs_.io_exuWriteback_20_bits_debug_isMMIO=0x%0h",this.io_exuWriteback_20_bits_debug_isMMIO,rhs_.io_exuWriteback_20_bits_debug_isMMIO),UVM_NONE)
        end

        if(this.io_exuWriteback_20_bits_debug_isNCIO!=rhs_.io_exuWriteback_20_bits_debug_isNCIO) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_20_bits_debug_isNCIO=0x%0h while the rhs_.io_exuWriteback_20_bits_debug_isNCIO=0x%0h",this.io_exuWriteback_20_bits_debug_isNCIO,rhs_.io_exuWriteback_20_bits_debug_isNCIO),UVM_NONE)
        end

        if(this.io_exuWriteback_20_bits_debug_isPerfCnt!=rhs_.io_exuWriteback_20_bits_debug_isPerfCnt) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_20_bits_debug_isPerfCnt=0x%0h while the rhs_.io_exuWriteback_20_bits_debug_isPerfCnt=0x%0h",this.io_exuWriteback_20_bits_debug_isPerfCnt,rhs_.io_exuWriteback_20_bits_debug_isPerfCnt),UVM_NONE)
        end

        if(this.io_exuWriteback_20_bits_debug_paddr!=rhs_.io_exuWriteback_20_bits_debug_paddr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_20_bits_debug_paddr=0x%0h while the rhs_.io_exuWriteback_20_bits_debug_paddr=0x%0h",this.io_exuWriteback_20_bits_debug_paddr,rhs_.io_exuWriteback_20_bits_debug_paddr),UVM_NONE)
        end

        if(this.io_exuWriteback_19_valid!=rhs_.io_exuWriteback_19_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_19_valid=0x%0h while the rhs_.io_exuWriteback_19_valid=0x%0h",this.io_exuWriteback_19_valid,rhs_.io_exuWriteback_19_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_19_bits_data_0!=rhs_.io_exuWriteback_19_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_19_bits_data_0=0x%0h while the rhs_.io_exuWriteback_19_bits_data_0=0x%0h",this.io_exuWriteback_19_bits_data_0,rhs_.io_exuWriteback_19_bits_data_0),UVM_NONE)
        end

        if(this.io_exuWriteback_19_bits_robIdx_value!=rhs_.io_exuWriteback_19_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_19_bits_robIdx_value=0x%0h while the rhs_.io_exuWriteback_19_bits_robIdx_value=0x%0h",this.io_exuWriteback_19_bits_robIdx_value,rhs_.io_exuWriteback_19_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_19_bits_sqIdx_value!=rhs_.io_exuWriteback_19_bits_sqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_19_bits_sqIdx_value=0x%0h while the rhs_.io_exuWriteback_19_bits_sqIdx_value=0x%0h",this.io_exuWriteback_19_bits_sqIdx_value,rhs_.io_exuWriteback_19_bits_sqIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_19_bits_debug_isMMIO!=rhs_.io_exuWriteback_19_bits_debug_isMMIO) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_19_bits_debug_isMMIO=0x%0h while the rhs_.io_exuWriteback_19_bits_debug_isMMIO=0x%0h",this.io_exuWriteback_19_bits_debug_isMMIO,rhs_.io_exuWriteback_19_bits_debug_isMMIO),UVM_NONE)
        end

        if(this.io_exuWriteback_19_bits_debug_isNCIO!=rhs_.io_exuWriteback_19_bits_debug_isNCIO) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_19_bits_debug_isNCIO=0x%0h while the rhs_.io_exuWriteback_19_bits_debug_isNCIO=0x%0h",this.io_exuWriteback_19_bits_debug_isNCIO,rhs_.io_exuWriteback_19_bits_debug_isNCIO),UVM_NONE)
        end

        if(this.io_exuWriteback_19_bits_debug_isPerfCnt!=rhs_.io_exuWriteback_19_bits_debug_isPerfCnt) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_19_bits_debug_isPerfCnt=0x%0h while the rhs_.io_exuWriteback_19_bits_debug_isPerfCnt=0x%0h",this.io_exuWriteback_19_bits_debug_isPerfCnt,rhs_.io_exuWriteback_19_bits_debug_isPerfCnt),UVM_NONE)
        end

        if(this.io_exuWriteback_19_bits_debug_paddr!=rhs_.io_exuWriteback_19_bits_debug_paddr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_19_bits_debug_paddr=0x%0h while the rhs_.io_exuWriteback_19_bits_debug_paddr=0x%0h",this.io_exuWriteback_19_bits_debug_paddr,rhs_.io_exuWriteback_19_bits_debug_paddr),UVM_NONE)
        end

        if(this.io_exuWriteback_18_valid!=rhs_.io_exuWriteback_18_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_18_valid=0x%0h while the rhs_.io_exuWriteback_18_valid=0x%0h",this.io_exuWriteback_18_valid,rhs_.io_exuWriteback_18_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_18_bits_data_0!=rhs_.io_exuWriteback_18_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_18_bits_data_0=0x%0h while the rhs_.io_exuWriteback_18_bits_data_0=0x%0h",this.io_exuWriteback_18_bits_data_0,rhs_.io_exuWriteback_18_bits_data_0),UVM_NONE)
        end

        if(this.io_exuWriteback_18_bits_robIdx_value!=rhs_.io_exuWriteback_18_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_18_bits_robIdx_value=0x%0h while the rhs_.io_exuWriteback_18_bits_robIdx_value=0x%0h",this.io_exuWriteback_18_bits_robIdx_value,rhs_.io_exuWriteback_18_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_18_bits_sqIdx_value!=rhs_.io_exuWriteback_18_bits_sqIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_18_bits_sqIdx_value=0x%0h while the rhs_.io_exuWriteback_18_bits_sqIdx_value=0x%0h",this.io_exuWriteback_18_bits_sqIdx_value,rhs_.io_exuWriteback_18_bits_sqIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_18_bits_debug_isMMIO!=rhs_.io_exuWriteback_18_bits_debug_isMMIO) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_18_bits_debug_isMMIO=0x%0h while the rhs_.io_exuWriteback_18_bits_debug_isMMIO=0x%0h",this.io_exuWriteback_18_bits_debug_isMMIO,rhs_.io_exuWriteback_18_bits_debug_isMMIO),UVM_NONE)
        end

        if(this.io_exuWriteback_18_bits_debug_isNCIO!=rhs_.io_exuWriteback_18_bits_debug_isNCIO) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_18_bits_debug_isNCIO=0x%0h while the rhs_.io_exuWriteback_18_bits_debug_isNCIO=0x%0h",this.io_exuWriteback_18_bits_debug_isNCIO,rhs_.io_exuWriteback_18_bits_debug_isNCIO),UVM_NONE)
        end

        if(this.io_exuWriteback_18_bits_debug_isPerfCnt!=rhs_.io_exuWriteback_18_bits_debug_isPerfCnt) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_18_bits_debug_isPerfCnt=0x%0h while the rhs_.io_exuWriteback_18_bits_debug_isPerfCnt=0x%0h",this.io_exuWriteback_18_bits_debug_isPerfCnt,rhs_.io_exuWriteback_18_bits_debug_isPerfCnt),UVM_NONE)
        end

        if(this.io_exuWriteback_18_bits_debug_paddr!=rhs_.io_exuWriteback_18_bits_debug_paddr) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_18_bits_debug_paddr=0x%0h while the rhs_.io_exuWriteback_18_bits_debug_paddr=0x%0h",this.io_exuWriteback_18_bits_debug_paddr,rhs_.io_exuWriteback_18_bits_debug_paddr),UVM_NONE)
        end

        if(this.io_exuWriteback_17_valid!=rhs_.io_exuWriteback_17_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_17_valid=0x%0h while the rhs_.io_exuWriteback_17_valid=0x%0h",this.io_exuWriteback_17_valid,rhs_.io_exuWriteback_17_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_17_bits_data_0!=rhs_.io_exuWriteback_17_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_17_bits_data_0=0x%0h while the rhs_.io_exuWriteback_17_bits_data_0=0x%0h",this.io_exuWriteback_17_bits_data_0,rhs_.io_exuWriteback_17_bits_data_0),UVM_NONE)
        end

        if(this.io_exuWriteback_17_bits_robIdx_value!=rhs_.io_exuWriteback_17_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_17_bits_robIdx_value=0x%0h while the rhs_.io_exuWriteback_17_bits_robIdx_value=0x%0h",this.io_exuWriteback_17_bits_robIdx_value,rhs_.io_exuWriteback_17_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_17_bits_fflags!=rhs_.io_exuWriteback_17_bits_fflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_17_bits_fflags=0x%0h while the rhs_.io_exuWriteback_17_bits_fflags=0x%0h",this.io_exuWriteback_17_bits_fflags,rhs_.io_exuWriteback_17_bits_fflags),UVM_NONE)
        end

        if(this.io_exuWriteback_17_bits_wflags!=rhs_.io_exuWriteback_17_bits_wflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_17_bits_wflags=0x%0h while the rhs_.io_exuWriteback_17_bits_wflags=0x%0h",this.io_exuWriteback_17_bits_wflags,rhs_.io_exuWriteback_17_bits_wflags),UVM_NONE)
        end

        if(this.io_exuWriteback_16_valid!=rhs_.io_exuWriteback_16_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_16_valid=0x%0h while the rhs_.io_exuWriteback_16_valid=0x%0h",this.io_exuWriteback_16_valid,rhs_.io_exuWriteback_16_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_16_bits_data_0!=rhs_.io_exuWriteback_16_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_16_bits_data_0=0x%0h while the rhs_.io_exuWriteback_16_bits_data_0=0x%0h",this.io_exuWriteback_16_bits_data_0,rhs_.io_exuWriteback_16_bits_data_0),UVM_NONE)
        end

        if(this.io_exuWriteback_16_bits_robIdx_value!=rhs_.io_exuWriteback_16_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_16_bits_robIdx_value=0x%0h while the rhs_.io_exuWriteback_16_bits_robIdx_value=0x%0h",this.io_exuWriteback_16_bits_robIdx_value,rhs_.io_exuWriteback_16_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_16_bits_fflags!=rhs_.io_exuWriteback_16_bits_fflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_16_bits_fflags=0x%0h while the rhs_.io_exuWriteback_16_bits_fflags=0x%0h",this.io_exuWriteback_16_bits_fflags,rhs_.io_exuWriteback_16_bits_fflags),UVM_NONE)
        end

        if(this.io_exuWriteback_16_bits_wflags!=rhs_.io_exuWriteback_16_bits_wflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_16_bits_wflags=0x%0h while the rhs_.io_exuWriteback_16_bits_wflags=0x%0h",this.io_exuWriteback_16_bits_wflags,rhs_.io_exuWriteback_16_bits_wflags),UVM_NONE)
        end

        if(this.io_exuWriteback_15_valid!=rhs_.io_exuWriteback_15_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_15_valid=0x%0h while the rhs_.io_exuWriteback_15_valid=0x%0h",this.io_exuWriteback_15_valid,rhs_.io_exuWriteback_15_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_15_bits_data_0!=rhs_.io_exuWriteback_15_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_15_bits_data_0=0x%0h while the rhs_.io_exuWriteback_15_bits_data_0=0x%0h",this.io_exuWriteback_15_bits_data_0,rhs_.io_exuWriteback_15_bits_data_0),UVM_NONE)
        end

        if(this.io_exuWriteback_15_bits_robIdx_value!=rhs_.io_exuWriteback_15_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_15_bits_robIdx_value=0x%0h while the rhs_.io_exuWriteback_15_bits_robIdx_value=0x%0h",this.io_exuWriteback_15_bits_robIdx_value,rhs_.io_exuWriteback_15_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_15_bits_fflags!=rhs_.io_exuWriteback_15_bits_fflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_15_bits_fflags=0x%0h while the rhs_.io_exuWriteback_15_bits_fflags=0x%0h",this.io_exuWriteback_15_bits_fflags,rhs_.io_exuWriteback_15_bits_fflags),UVM_NONE)
        end

        if(this.io_exuWriteback_15_bits_wflags!=rhs_.io_exuWriteback_15_bits_wflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_15_bits_wflags=0x%0h while the rhs_.io_exuWriteback_15_bits_wflags=0x%0h",this.io_exuWriteback_15_bits_wflags,rhs_.io_exuWriteback_15_bits_wflags),UVM_NONE)
        end

        if(this.io_exuWriteback_15_bits_vxsat!=rhs_.io_exuWriteback_15_bits_vxsat) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_15_bits_vxsat=0x%0h while the rhs_.io_exuWriteback_15_bits_vxsat=0x%0h",this.io_exuWriteback_15_bits_vxsat,rhs_.io_exuWriteback_15_bits_vxsat),UVM_NONE)
        end

        if(this.io_exuWriteback_14_valid!=rhs_.io_exuWriteback_14_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_14_valid=0x%0h while the rhs_.io_exuWriteback_14_valid=0x%0h",this.io_exuWriteback_14_valid,rhs_.io_exuWriteback_14_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_14_bits_data_0!=rhs_.io_exuWriteback_14_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_14_bits_data_0=0x%0h while the rhs_.io_exuWriteback_14_bits_data_0=0x%0h",this.io_exuWriteback_14_bits_data_0,rhs_.io_exuWriteback_14_bits_data_0),UVM_NONE)
        end

        if(this.io_exuWriteback_14_bits_robIdx_value!=rhs_.io_exuWriteback_14_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_14_bits_robIdx_value=0x%0h while the rhs_.io_exuWriteback_14_bits_robIdx_value=0x%0h",this.io_exuWriteback_14_bits_robIdx_value,rhs_.io_exuWriteback_14_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_14_bits_fflags!=rhs_.io_exuWriteback_14_bits_fflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_14_bits_fflags=0x%0h while the rhs_.io_exuWriteback_14_bits_fflags=0x%0h",this.io_exuWriteback_14_bits_fflags,rhs_.io_exuWriteback_14_bits_fflags),UVM_NONE)
        end

        if(this.io_exuWriteback_14_bits_wflags!=rhs_.io_exuWriteback_14_bits_wflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_14_bits_wflags=0x%0h while the rhs_.io_exuWriteback_14_bits_wflags=0x%0h",this.io_exuWriteback_14_bits_wflags,rhs_.io_exuWriteback_14_bits_wflags),UVM_NONE)
        end

        if(this.io_exuWriteback_13_valid!=rhs_.io_exuWriteback_13_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_13_valid=0x%0h while the rhs_.io_exuWriteback_13_valid=0x%0h",this.io_exuWriteback_13_valid,rhs_.io_exuWriteback_13_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_13_bits_data_0!=rhs_.io_exuWriteback_13_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_13_bits_data_0=0x%0h while the rhs_.io_exuWriteback_13_bits_data_0=0x%0h",this.io_exuWriteback_13_bits_data_0,rhs_.io_exuWriteback_13_bits_data_0),UVM_NONE)
        end

        if(this.io_exuWriteback_13_bits_robIdx_value!=rhs_.io_exuWriteback_13_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_13_bits_robIdx_value=0x%0h while the rhs_.io_exuWriteback_13_bits_robIdx_value=0x%0h",this.io_exuWriteback_13_bits_robIdx_value,rhs_.io_exuWriteback_13_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_13_bits_fflags!=rhs_.io_exuWriteback_13_bits_fflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_13_bits_fflags=0x%0h while the rhs_.io_exuWriteback_13_bits_fflags=0x%0h",this.io_exuWriteback_13_bits_fflags,rhs_.io_exuWriteback_13_bits_fflags),UVM_NONE)
        end

        if(this.io_exuWriteback_13_bits_wflags!=rhs_.io_exuWriteback_13_bits_wflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_13_bits_wflags=0x%0h while the rhs_.io_exuWriteback_13_bits_wflags=0x%0h",this.io_exuWriteback_13_bits_wflags,rhs_.io_exuWriteback_13_bits_wflags),UVM_NONE)
        end

        if(this.io_exuWriteback_13_bits_vxsat!=rhs_.io_exuWriteback_13_bits_vxsat) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_13_bits_vxsat=0x%0h while the rhs_.io_exuWriteback_13_bits_vxsat=0x%0h",this.io_exuWriteback_13_bits_vxsat,rhs_.io_exuWriteback_13_bits_vxsat),UVM_NONE)
        end

        if(this.io_exuWriteback_12_valid!=rhs_.io_exuWriteback_12_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_12_valid=0x%0h while the rhs_.io_exuWriteback_12_valid=0x%0h",this.io_exuWriteback_12_valid,rhs_.io_exuWriteback_12_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_12_bits_data_0!=rhs_.io_exuWriteback_12_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_12_bits_data_0=0x%0h while the rhs_.io_exuWriteback_12_bits_data_0=0x%0h",this.io_exuWriteback_12_bits_data_0,rhs_.io_exuWriteback_12_bits_data_0),UVM_NONE)
        end

        if(this.io_exuWriteback_12_bits_robIdx_value!=rhs_.io_exuWriteback_12_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_12_bits_robIdx_value=0x%0h while the rhs_.io_exuWriteback_12_bits_robIdx_value=0x%0h",this.io_exuWriteback_12_bits_robIdx_value,rhs_.io_exuWriteback_12_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_12_bits_fflags!=rhs_.io_exuWriteback_12_bits_fflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_12_bits_fflags=0x%0h while the rhs_.io_exuWriteback_12_bits_fflags=0x%0h",this.io_exuWriteback_12_bits_fflags,rhs_.io_exuWriteback_12_bits_fflags),UVM_NONE)
        end

        if(this.io_exuWriteback_12_bits_wflags!=rhs_.io_exuWriteback_12_bits_wflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_12_bits_wflags=0x%0h while the rhs_.io_exuWriteback_12_bits_wflags=0x%0h",this.io_exuWriteback_12_bits_wflags,rhs_.io_exuWriteback_12_bits_wflags),UVM_NONE)
        end

        if(this.io_exuWriteback_11_valid!=rhs_.io_exuWriteback_11_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_11_valid=0x%0h while the rhs_.io_exuWriteback_11_valid=0x%0h",this.io_exuWriteback_11_valid,rhs_.io_exuWriteback_11_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_11_bits_data_0!=rhs_.io_exuWriteback_11_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_11_bits_data_0=0x%0h while the rhs_.io_exuWriteback_11_bits_data_0=0x%0h",this.io_exuWriteback_11_bits_data_0,rhs_.io_exuWriteback_11_bits_data_0),UVM_NONE)
        end

        if(this.io_exuWriteback_11_bits_robIdx_value!=rhs_.io_exuWriteback_11_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_11_bits_robIdx_value=0x%0h while the rhs_.io_exuWriteback_11_bits_robIdx_value=0x%0h",this.io_exuWriteback_11_bits_robIdx_value,rhs_.io_exuWriteback_11_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_11_bits_fflags!=rhs_.io_exuWriteback_11_bits_fflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_11_bits_fflags=0x%0h while the rhs_.io_exuWriteback_11_bits_fflags=0x%0h",this.io_exuWriteback_11_bits_fflags,rhs_.io_exuWriteback_11_bits_fflags),UVM_NONE)
        end

        if(this.io_exuWriteback_11_bits_wflags!=rhs_.io_exuWriteback_11_bits_wflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_11_bits_wflags=0x%0h while the rhs_.io_exuWriteback_11_bits_wflags=0x%0h",this.io_exuWriteback_11_bits_wflags,rhs_.io_exuWriteback_11_bits_wflags),UVM_NONE)
        end

        if(this.io_exuWriteback_10_valid!=rhs_.io_exuWriteback_10_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_10_valid=0x%0h while the rhs_.io_exuWriteback_10_valid=0x%0h",this.io_exuWriteback_10_valid,rhs_.io_exuWriteback_10_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_10_bits_data_0!=rhs_.io_exuWriteback_10_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_10_bits_data_0=0x%0h while the rhs_.io_exuWriteback_10_bits_data_0=0x%0h",this.io_exuWriteback_10_bits_data_0,rhs_.io_exuWriteback_10_bits_data_0),UVM_NONE)
        end

        if(this.io_exuWriteback_10_bits_robIdx_value!=rhs_.io_exuWriteback_10_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_10_bits_robIdx_value=0x%0h while the rhs_.io_exuWriteback_10_bits_robIdx_value=0x%0h",this.io_exuWriteback_10_bits_robIdx_value,rhs_.io_exuWriteback_10_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_10_bits_fflags!=rhs_.io_exuWriteback_10_bits_fflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_10_bits_fflags=0x%0h while the rhs_.io_exuWriteback_10_bits_fflags=0x%0h",this.io_exuWriteback_10_bits_fflags,rhs_.io_exuWriteback_10_bits_fflags),UVM_NONE)
        end

        if(this.io_exuWriteback_10_bits_wflags!=rhs_.io_exuWriteback_10_bits_wflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_10_bits_wflags=0x%0h while the rhs_.io_exuWriteback_10_bits_wflags=0x%0h",this.io_exuWriteback_10_bits_wflags,rhs_.io_exuWriteback_10_bits_wflags),UVM_NONE)
        end

        if(this.io_exuWriteback_9_valid!=rhs_.io_exuWriteback_9_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_9_valid=0x%0h while the rhs_.io_exuWriteback_9_valid=0x%0h",this.io_exuWriteback_9_valid,rhs_.io_exuWriteback_9_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_9_bits_data_0!=rhs_.io_exuWriteback_9_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_9_bits_data_0=0x%0h while the rhs_.io_exuWriteback_9_bits_data_0=0x%0h",this.io_exuWriteback_9_bits_data_0,rhs_.io_exuWriteback_9_bits_data_0),UVM_NONE)
        end

        if(this.io_exuWriteback_9_bits_robIdx_value!=rhs_.io_exuWriteback_9_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_9_bits_robIdx_value=0x%0h while the rhs_.io_exuWriteback_9_bits_robIdx_value=0x%0h",this.io_exuWriteback_9_bits_robIdx_value,rhs_.io_exuWriteback_9_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_9_bits_fflags!=rhs_.io_exuWriteback_9_bits_fflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_9_bits_fflags=0x%0h while the rhs_.io_exuWriteback_9_bits_fflags=0x%0h",this.io_exuWriteback_9_bits_fflags,rhs_.io_exuWriteback_9_bits_fflags),UVM_NONE)
        end

        if(this.io_exuWriteback_9_bits_wflags!=rhs_.io_exuWriteback_9_bits_wflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_9_bits_wflags=0x%0h while the rhs_.io_exuWriteback_9_bits_wflags=0x%0h",this.io_exuWriteback_9_bits_wflags,rhs_.io_exuWriteback_9_bits_wflags),UVM_NONE)
        end

        if(this.io_exuWriteback_8_valid!=rhs_.io_exuWriteback_8_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_8_valid=0x%0h while the rhs_.io_exuWriteback_8_valid=0x%0h",this.io_exuWriteback_8_valid,rhs_.io_exuWriteback_8_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_8_bits_data_0!=rhs_.io_exuWriteback_8_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_8_bits_data_0=0x%0h while the rhs_.io_exuWriteback_8_bits_data_0=0x%0h",this.io_exuWriteback_8_bits_data_0,rhs_.io_exuWriteback_8_bits_data_0),UVM_NONE)
        end

        if(this.io_exuWriteback_8_bits_robIdx_value!=rhs_.io_exuWriteback_8_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_8_bits_robIdx_value=0x%0h while the rhs_.io_exuWriteback_8_bits_robIdx_value=0x%0h",this.io_exuWriteback_8_bits_robIdx_value,rhs_.io_exuWriteback_8_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_8_bits_fflags!=rhs_.io_exuWriteback_8_bits_fflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_8_bits_fflags=0x%0h while the rhs_.io_exuWriteback_8_bits_fflags=0x%0h",this.io_exuWriteback_8_bits_fflags,rhs_.io_exuWriteback_8_bits_fflags),UVM_NONE)
        end

        if(this.io_exuWriteback_8_bits_wflags!=rhs_.io_exuWriteback_8_bits_wflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_8_bits_wflags=0x%0h while the rhs_.io_exuWriteback_8_bits_wflags=0x%0h",this.io_exuWriteback_8_bits_wflags,rhs_.io_exuWriteback_8_bits_wflags),UVM_NONE)
        end

        if(this.io_exuWriteback_7_valid!=rhs_.io_exuWriteback_7_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_7_valid=0x%0h while the rhs_.io_exuWriteback_7_valid=0x%0h",this.io_exuWriteback_7_valid,rhs_.io_exuWriteback_7_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_7_bits_data_0!=rhs_.io_exuWriteback_7_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_7_bits_data_0=0x%0h while the rhs_.io_exuWriteback_7_bits_data_0=0x%0h",this.io_exuWriteback_7_bits_data_0,rhs_.io_exuWriteback_7_bits_data_0),UVM_NONE)
        end

        if(this.io_exuWriteback_7_bits_robIdx_value!=rhs_.io_exuWriteback_7_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_7_bits_robIdx_value=0x%0h while the rhs_.io_exuWriteback_7_bits_robIdx_value=0x%0h",this.io_exuWriteback_7_bits_robIdx_value,rhs_.io_exuWriteback_7_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_7_bits_debug_isPerfCnt!=rhs_.io_exuWriteback_7_bits_debug_isPerfCnt) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_7_bits_debug_isPerfCnt=0x%0h while the rhs_.io_exuWriteback_7_bits_debug_isPerfCnt=0x%0h",this.io_exuWriteback_7_bits_debug_isPerfCnt,rhs_.io_exuWriteback_7_bits_debug_isPerfCnt),UVM_NONE)
        end

        if(this.io_exuWriteback_6_valid!=rhs_.io_exuWriteback_6_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_6_valid=0x%0h while the rhs_.io_exuWriteback_6_valid=0x%0h",this.io_exuWriteback_6_valid,rhs_.io_exuWriteback_6_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_6_bits_data_0!=rhs_.io_exuWriteback_6_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_6_bits_data_0=0x%0h while the rhs_.io_exuWriteback_6_bits_data_0=0x%0h",this.io_exuWriteback_6_bits_data_0,rhs_.io_exuWriteback_6_bits_data_0),UVM_NONE)
        end

        if(this.io_exuWriteback_6_bits_robIdx_value!=rhs_.io_exuWriteback_6_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_6_bits_robIdx_value=0x%0h while the rhs_.io_exuWriteback_6_bits_robIdx_value=0x%0h",this.io_exuWriteback_6_bits_robIdx_value,rhs_.io_exuWriteback_6_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_5_valid!=rhs_.io_exuWriteback_5_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_5_valid=0x%0h while the rhs_.io_exuWriteback_5_valid=0x%0h",this.io_exuWriteback_5_valid,rhs_.io_exuWriteback_5_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_5_bits_data_0!=rhs_.io_exuWriteback_5_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_5_bits_data_0=0x%0h while the rhs_.io_exuWriteback_5_bits_data_0=0x%0h",this.io_exuWriteback_5_bits_data_0,rhs_.io_exuWriteback_5_bits_data_0),UVM_NONE)
        end

        if(this.io_exuWriteback_5_bits_robIdx_value!=rhs_.io_exuWriteback_5_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_5_bits_robIdx_value=0x%0h while the rhs_.io_exuWriteback_5_bits_robIdx_value=0x%0h",this.io_exuWriteback_5_bits_robIdx_value,rhs_.io_exuWriteback_5_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_5_bits_redirect_valid!=rhs_.io_exuWriteback_5_bits_redirect_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_5_bits_redirect_valid=0x%0h while the rhs_.io_exuWriteback_5_bits_redirect_valid=0x%0h",this.io_exuWriteback_5_bits_redirect_valid,rhs_.io_exuWriteback_5_bits_redirect_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken!=rhs_.io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken=0x%0h while the rhs_.io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken=0x%0h",this.io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken,rhs_.io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken),UVM_NONE)
        end

        if(this.io_exuWriteback_5_bits_fflags!=rhs_.io_exuWriteback_5_bits_fflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_5_bits_fflags=0x%0h while the rhs_.io_exuWriteback_5_bits_fflags=0x%0h",this.io_exuWriteback_5_bits_fflags,rhs_.io_exuWriteback_5_bits_fflags),UVM_NONE)
        end

        if(this.io_exuWriteback_5_bits_wflags!=rhs_.io_exuWriteback_5_bits_wflags) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_5_bits_wflags=0x%0h while the rhs_.io_exuWriteback_5_bits_wflags=0x%0h",this.io_exuWriteback_5_bits_wflags,rhs_.io_exuWriteback_5_bits_wflags),UVM_NONE)
        end

        if(this.io_exuWriteback_4_valid!=rhs_.io_exuWriteback_4_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_4_valid=0x%0h while the rhs_.io_exuWriteback_4_valid=0x%0h",this.io_exuWriteback_4_valid,rhs_.io_exuWriteback_4_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_4_bits_data_0!=rhs_.io_exuWriteback_4_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_4_bits_data_0=0x%0h while the rhs_.io_exuWriteback_4_bits_data_0=0x%0h",this.io_exuWriteback_4_bits_data_0,rhs_.io_exuWriteback_4_bits_data_0),UVM_NONE)
        end

        if(this.io_exuWriteback_4_bits_robIdx_value!=rhs_.io_exuWriteback_4_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_4_bits_robIdx_value=0x%0h while the rhs_.io_exuWriteback_4_bits_robIdx_value=0x%0h",this.io_exuWriteback_4_bits_robIdx_value,rhs_.io_exuWriteback_4_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_3_valid!=rhs_.io_exuWriteback_3_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_3_valid=0x%0h while the rhs_.io_exuWriteback_3_valid=0x%0h",this.io_exuWriteback_3_valid,rhs_.io_exuWriteback_3_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_3_bits_data_0!=rhs_.io_exuWriteback_3_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_3_bits_data_0=0x%0h while the rhs_.io_exuWriteback_3_bits_data_0=0x%0h",this.io_exuWriteback_3_bits_data_0,rhs_.io_exuWriteback_3_bits_data_0),UVM_NONE)
        end

        if(this.io_exuWriteback_3_bits_robIdx_value!=rhs_.io_exuWriteback_3_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_3_bits_robIdx_value=0x%0h while the rhs_.io_exuWriteback_3_bits_robIdx_value=0x%0h",this.io_exuWriteback_3_bits_robIdx_value,rhs_.io_exuWriteback_3_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_3_bits_redirect_valid!=rhs_.io_exuWriteback_3_bits_redirect_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_3_bits_redirect_valid=0x%0h while the rhs_.io_exuWriteback_3_bits_redirect_valid=0x%0h",this.io_exuWriteback_3_bits_redirect_valid,rhs_.io_exuWriteback_3_bits_redirect_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken!=rhs_.io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken=0x%0h while the rhs_.io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken=0x%0h",this.io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken,rhs_.io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken),UVM_NONE)
        end

        if(this.io_exuWriteback_2_valid!=rhs_.io_exuWriteback_2_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_2_valid=0x%0h while the rhs_.io_exuWriteback_2_valid=0x%0h",this.io_exuWriteback_2_valid,rhs_.io_exuWriteback_2_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_2_bits_data_0!=rhs_.io_exuWriteback_2_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_2_bits_data_0=0x%0h while the rhs_.io_exuWriteback_2_bits_data_0=0x%0h",this.io_exuWriteback_2_bits_data_0,rhs_.io_exuWriteback_2_bits_data_0),UVM_NONE)
        end

        if(this.io_exuWriteback_2_bits_robIdx_value!=rhs_.io_exuWriteback_2_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_2_bits_robIdx_value=0x%0h while the rhs_.io_exuWriteback_2_bits_robIdx_value=0x%0h",this.io_exuWriteback_2_bits_robIdx_value,rhs_.io_exuWriteback_2_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_1_valid!=rhs_.io_exuWriteback_1_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_1_valid=0x%0h while the rhs_.io_exuWriteback_1_valid=0x%0h",this.io_exuWriteback_1_valid,rhs_.io_exuWriteback_1_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_1_bits_data_0!=rhs_.io_exuWriteback_1_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_1_bits_data_0=0x%0h while the rhs_.io_exuWriteback_1_bits_data_0=0x%0h",this.io_exuWriteback_1_bits_data_0,rhs_.io_exuWriteback_1_bits_data_0),UVM_NONE)
        end

        if(this.io_exuWriteback_1_bits_robIdx_value!=rhs_.io_exuWriteback_1_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_1_bits_robIdx_value=0x%0h while the rhs_.io_exuWriteback_1_bits_robIdx_value=0x%0h",this.io_exuWriteback_1_bits_robIdx_value,rhs_.io_exuWriteback_1_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_exuWriteback_1_bits_redirect_valid!=rhs_.io_exuWriteback_1_bits_redirect_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_1_bits_redirect_valid=0x%0h while the rhs_.io_exuWriteback_1_bits_redirect_valid=0x%0h",this.io_exuWriteback_1_bits_redirect_valid,rhs_.io_exuWriteback_1_bits_redirect_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken!=rhs_.io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken=0x%0h while the rhs_.io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken=0x%0h",this.io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken,rhs_.io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken),UVM_NONE)
        end

        if(this.io_exuWriteback_0_valid!=rhs_.io_exuWriteback_0_valid) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_0_valid=0x%0h while the rhs_.io_exuWriteback_0_valid=0x%0h",this.io_exuWriteback_0_valid,rhs_.io_exuWriteback_0_valid),UVM_NONE)
        end

        if(this.io_exuWriteback_0_bits_data_0!=rhs_.io_exuWriteback_0_bits_data_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_0_bits_data_0=0x%0h while the rhs_.io_exuWriteback_0_bits_data_0=0x%0h",this.io_exuWriteback_0_bits_data_0,rhs_.io_exuWriteback_0_bits_data_0),UVM_NONE)
        end

        if(this.io_exuWriteback_0_bits_robIdx_value!=rhs_.io_exuWriteback_0_bits_robIdx_value) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_exuWriteback_0_bits_robIdx_value=0x%0h while the rhs_.io_exuWriteback_0_bits_robIdx_value=0x%0h",this.io_exuWriteback_0_bits_robIdx_value,rhs_.io_exuWriteback_0_bits_robIdx_value),UVM_NONE)
        end

        if(this.io_writebackNums_0_bits!=rhs_.io_writebackNums_0_bits) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNums_0_bits=0x%0h while the rhs_.io_writebackNums_0_bits=0x%0h",this.io_writebackNums_0_bits,rhs_.io_writebackNums_0_bits),UVM_NONE)
        end

        if(this.io_writebackNums_1_bits!=rhs_.io_writebackNums_1_bits) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNums_1_bits=0x%0h while the rhs_.io_writebackNums_1_bits=0x%0h",this.io_writebackNums_1_bits,rhs_.io_writebackNums_1_bits),UVM_NONE)
        end

        if(this.io_writebackNums_2_bits!=rhs_.io_writebackNums_2_bits) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNums_2_bits=0x%0h while the rhs_.io_writebackNums_2_bits=0x%0h",this.io_writebackNums_2_bits,rhs_.io_writebackNums_2_bits),UVM_NONE)
        end

        if(this.io_writebackNums_3_bits!=rhs_.io_writebackNums_3_bits) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNums_3_bits=0x%0h while the rhs_.io_writebackNums_3_bits=0x%0h",this.io_writebackNums_3_bits,rhs_.io_writebackNums_3_bits),UVM_NONE)
        end

        if(this.io_writebackNums_4_bits!=rhs_.io_writebackNums_4_bits) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNums_4_bits=0x%0h while the rhs_.io_writebackNums_4_bits=0x%0h",this.io_writebackNums_4_bits,rhs_.io_writebackNums_4_bits),UVM_NONE)
        end

        if(this.io_writebackNums_5_bits!=rhs_.io_writebackNums_5_bits) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNums_5_bits=0x%0h while the rhs_.io_writebackNums_5_bits=0x%0h",this.io_writebackNums_5_bits,rhs_.io_writebackNums_5_bits),UVM_NONE)
        end

        if(this.io_writebackNums_6_bits!=rhs_.io_writebackNums_6_bits) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNums_6_bits=0x%0h while the rhs_.io_writebackNums_6_bits=0x%0h",this.io_writebackNums_6_bits,rhs_.io_writebackNums_6_bits),UVM_NONE)
        end

        if(this.io_writebackNums_7_bits!=rhs_.io_writebackNums_7_bits) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNums_7_bits=0x%0h while the rhs_.io_writebackNums_7_bits=0x%0h",this.io_writebackNums_7_bits,rhs_.io_writebackNums_7_bits),UVM_NONE)
        end

        if(this.io_writebackNums_8_bits!=rhs_.io_writebackNums_8_bits) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNums_8_bits=0x%0h while the rhs_.io_writebackNums_8_bits=0x%0h",this.io_writebackNums_8_bits,rhs_.io_writebackNums_8_bits),UVM_NONE)
        end

        if(this.io_writebackNums_9_bits!=rhs_.io_writebackNums_9_bits) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNums_9_bits=0x%0h while the rhs_.io_writebackNums_9_bits=0x%0h",this.io_writebackNums_9_bits,rhs_.io_writebackNums_9_bits),UVM_NONE)
        end

        if(this.io_writebackNums_10_bits!=rhs_.io_writebackNums_10_bits) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNums_10_bits=0x%0h while the rhs_.io_writebackNums_10_bits=0x%0h",this.io_writebackNums_10_bits,rhs_.io_writebackNums_10_bits),UVM_NONE)
        end

        if(this.io_writebackNums_11_bits!=rhs_.io_writebackNums_11_bits) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNums_11_bits=0x%0h while the rhs_.io_writebackNums_11_bits=0x%0h",this.io_writebackNums_11_bits,rhs_.io_writebackNums_11_bits),UVM_NONE)
        end

        if(this.io_writebackNums_12_bits!=rhs_.io_writebackNums_12_bits) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNums_12_bits=0x%0h while the rhs_.io_writebackNums_12_bits=0x%0h",this.io_writebackNums_12_bits,rhs_.io_writebackNums_12_bits),UVM_NONE)
        end

        if(this.io_writebackNums_13_bits!=rhs_.io_writebackNums_13_bits) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNums_13_bits=0x%0h while the rhs_.io_writebackNums_13_bits=0x%0h",this.io_writebackNums_13_bits,rhs_.io_writebackNums_13_bits),UVM_NONE)
        end

        if(this.io_writebackNums_14_bits!=rhs_.io_writebackNums_14_bits) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNums_14_bits=0x%0h while the rhs_.io_writebackNums_14_bits=0x%0h",this.io_writebackNums_14_bits,rhs_.io_writebackNums_14_bits),UVM_NONE)
        end

        if(this.io_writebackNums_15_bits!=rhs_.io_writebackNums_15_bits) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNums_15_bits=0x%0h while the rhs_.io_writebackNums_15_bits=0x%0h",this.io_writebackNums_15_bits,rhs_.io_writebackNums_15_bits),UVM_NONE)
        end

        if(this.io_writebackNums_16_bits!=rhs_.io_writebackNums_16_bits) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNums_16_bits=0x%0h while the rhs_.io_writebackNums_16_bits=0x%0h",this.io_writebackNums_16_bits,rhs_.io_writebackNums_16_bits),UVM_NONE)
        end

        if(this.io_writebackNums_17_bits!=rhs_.io_writebackNums_17_bits) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNums_17_bits=0x%0h while the rhs_.io_writebackNums_17_bits=0x%0h",this.io_writebackNums_17_bits,rhs_.io_writebackNums_17_bits),UVM_NONE)
        end

        if(this.io_writebackNums_18_bits!=rhs_.io_writebackNums_18_bits) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNums_18_bits=0x%0h while the rhs_.io_writebackNums_18_bits=0x%0h",this.io_writebackNums_18_bits,rhs_.io_writebackNums_18_bits),UVM_NONE)
        end

        if(this.io_writebackNums_19_bits!=rhs_.io_writebackNums_19_bits) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNums_19_bits=0x%0h while the rhs_.io_writebackNums_19_bits=0x%0h",this.io_writebackNums_19_bits,rhs_.io_writebackNums_19_bits),UVM_NONE)
        end

        if(this.io_writebackNums_20_bits!=rhs_.io_writebackNums_20_bits) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNums_20_bits=0x%0h while the rhs_.io_writebackNums_20_bits=0x%0h",this.io_writebackNums_20_bits,rhs_.io_writebackNums_20_bits),UVM_NONE)
        end

        if(this.io_writebackNums_21_bits!=rhs_.io_writebackNums_21_bits) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNums_21_bits=0x%0h while the rhs_.io_writebackNums_21_bits=0x%0h",this.io_writebackNums_21_bits,rhs_.io_writebackNums_21_bits),UVM_NONE)
        end

        if(this.io_writebackNums_22_bits!=rhs_.io_writebackNums_22_bits) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNums_22_bits=0x%0h while the rhs_.io_writebackNums_22_bits=0x%0h",this.io_writebackNums_22_bits,rhs_.io_writebackNums_22_bits),UVM_NONE)
        end

        if(this.io_writebackNums_23_bits!=rhs_.io_writebackNums_23_bits) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNums_23_bits=0x%0h while the rhs_.io_writebackNums_23_bits=0x%0h",this.io_writebackNums_23_bits,rhs_.io_writebackNums_23_bits),UVM_NONE)
        end

        if(this.io_writebackNums_24_bits!=rhs_.io_writebackNums_24_bits) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNums_24_bits=0x%0h while the rhs_.io_writebackNums_24_bits=0x%0h",this.io_writebackNums_24_bits,rhs_.io_writebackNums_24_bits),UVM_NONE)
        end

        if(this.io_writebackNeedFlush_0!=rhs_.io_writebackNeedFlush_0) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNeedFlush_0=0x%0h while the rhs_.io_writebackNeedFlush_0=0x%0h",this.io_writebackNeedFlush_0,rhs_.io_writebackNeedFlush_0),UVM_NONE)
        end

        if(this.io_writebackNeedFlush_1!=rhs_.io_writebackNeedFlush_1) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNeedFlush_1=0x%0h while the rhs_.io_writebackNeedFlush_1=0x%0h",this.io_writebackNeedFlush_1,rhs_.io_writebackNeedFlush_1),UVM_NONE)
        end

        if(this.io_writebackNeedFlush_2!=rhs_.io_writebackNeedFlush_2) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNeedFlush_2=0x%0h while the rhs_.io_writebackNeedFlush_2=0x%0h",this.io_writebackNeedFlush_2,rhs_.io_writebackNeedFlush_2),UVM_NONE)
        end

        if(this.io_writebackNeedFlush_6!=rhs_.io_writebackNeedFlush_6) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNeedFlush_6=0x%0h while the rhs_.io_writebackNeedFlush_6=0x%0h",this.io_writebackNeedFlush_6,rhs_.io_writebackNeedFlush_6),UVM_NONE)
        end

        if(this.io_writebackNeedFlush_7!=rhs_.io_writebackNeedFlush_7) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNeedFlush_7=0x%0h while the rhs_.io_writebackNeedFlush_7=0x%0h",this.io_writebackNeedFlush_7,rhs_.io_writebackNeedFlush_7),UVM_NONE)
        end

        if(this.io_writebackNeedFlush_8!=rhs_.io_writebackNeedFlush_8) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNeedFlush_8=0x%0h while the rhs_.io_writebackNeedFlush_8=0x%0h",this.io_writebackNeedFlush_8,rhs_.io_writebackNeedFlush_8),UVM_NONE)
        end

        if(this.io_writebackNeedFlush_9!=rhs_.io_writebackNeedFlush_9) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNeedFlush_9=0x%0h while the rhs_.io_writebackNeedFlush_9=0x%0h",this.io_writebackNeedFlush_9,rhs_.io_writebackNeedFlush_9),UVM_NONE)
        end

        if(this.io_writebackNeedFlush_10!=rhs_.io_writebackNeedFlush_10) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNeedFlush_10=0x%0h while the rhs_.io_writebackNeedFlush_10=0x%0h",this.io_writebackNeedFlush_10,rhs_.io_writebackNeedFlush_10),UVM_NONE)
        end

        if(this.io_writebackNeedFlush_11!=rhs_.io_writebackNeedFlush_11) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNeedFlush_11=0x%0h while the rhs_.io_writebackNeedFlush_11=0x%0h",this.io_writebackNeedFlush_11,rhs_.io_writebackNeedFlush_11),UVM_NONE)
        end

        if(this.io_writebackNeedFlush_12!=rhs_.io_writebackNeedFlush_12) begin
            super_result = 0;
            `uvm_info(get_type_name(),$sformatf("compare fail for this.io_writebackNeedFlush_12=0x%0h while the rhs_.io_writebackNeedFlush_12=0x%0h",this.io_writebackNeedFlush_12,rhs_.io_writebackNeedFlush_12),UVM_NONE)
        end

    end
    return super_result;
endfunction:compare

`endif


//=========================================================
//File name    : rename_in_connect.sv
//Author       : nanyunhao
//Module name  : rename_in_connect
//Discribution : rename_in_connect : rename_in Interface connection macro
//Date         : 2026-01-22
//=========================================================
`ifndef RENAME_IN_CONNECT__SV
`define RENAME_IN_CONNECT__SV

`define ROB__RENAME_IN_CONNECT(U_IF_NAME,AGENT_PATH,RTL_PATH) \
    rename_in_agent_interface  U_IF_NAME (clk,tc_if.rst_n); \
    initial begin \
        uvm_config_db#(virtual rename_in_agent_interface)::set(null,`"*AGENT_PATH*`", "vif", U_IF_NAME); \
    end \
    `ifdef ROB_UT \
    initial begin \
        force RTL_PATH.clock = U_IF_NAME.clock; \
        force RTL_PATH.reset = U_IF_NAME.reset; \
        force RTL_PATH.io_hartId = U_IF_NAME.io_hartId; \
        force RTL_PATH.io_enq_req_0_valid = U_IF_NAME.io_enq_req_0_valid; \
        force RTL_PATH.io_enq_req_0_bits_instr = U_IF_NAME.io_enq_req_0_bits_instr; \
        force RTL_PATH.io_enq_req_0_bits_pc = U_IF_NAME.io_enq_req_0_bits_pc; \
        force RTL_PATH.io_enq_req_0_bits_exceptionVec_0 = U_IF_NAME.io_enq_req_0_bits_exceptionVec_0; \
        force RTL_PATH.io_enq_req_0_bits_exceptionVec_1 = U_IF_NAME.io_enq_req_0_bits_exceptionVec_1; \
        force RTL_PATH.io_enq_req_0_bits_exceptionVec_2 = U_IF_NAME.io_enq_req_0_bits_exceptionVec_2; \
        force RTL_PATH.io_enq_req_0_bits_exceptionVec_3 = U_IF_NAME.io_enq_req_0_bits_exceptionVec_3; \
        force RTL_PATH.io_enq_req_0_bits_exceptionVec_12 = U_IF_NAME.io_enq_req_0_bits_exceptionVec_12; \
        force RTL_PATH.io_enq_req_0_bits_exceptionVec_20 = U_IF_NAME.io_enq_req_0_bits_exceptionVec_20; \
        force RTL_PATH.io_enq_req_0_bits_exceptionVec_22 = U_IF_NAME.io_enq_req_0_bits_exceptionVec_22; \
        force RTL_PATH.io_enq_req_0_bits_isFetchMalAddr = U_IF_NAME.io_enq_req_0_bits_isFetchMalAddr; \
        force RTL_PATH.io_enq_req_0_bits_hasException = U_IF_NAME.io_enq_req_0_bits_hasException; \
        force RTL_PATH.io_enq_req_0_bits_trigger = U_IF_NAME.io_enq_req_0_bits_trigger; \
        force RTL_PATH.io_enq_req_0_bits_preDecodeInfo_isRVC = U_IF_NAME.io_enq_req_0_bits_preDecodeInfo_isRVC; \
        force RTL_PATH.io_enq_req_0_bits_crossPageIPFFix = U_IF_NAME.io_enq_req_0_bits_crossPageIPFFix; \
        force RTL_PATH.io_enq_req_0_bits_ftqPtr_flag = U_IF_NAME.io_enq_req_0_bits_ftqPtr_flag; \
        force RTL_PATH.io_enq_req_0_bits_ftqPtr_value = U_IF_NAME.io_enq_req_0_bits_ftqPtr_value; \
        force RTL_PATH.io_enq_req_0_bits_ftqOffset = U_IF_NAME.io_enq_req_0_bits_ftqOffset; \
        force RTL_PATH.io_enq_req_0_bits_ldest = U_IF_NAME.io_enq_req_0_bits_ldest; \
        force RTL_PATH.io_enq_req_0_bits_fuType = U_IF_NAME.io_enq_req_0_bits_fuType; \
        force RTL_PATH.io_enq_req_0_bits_fuOpType = U_IF_NAME.io_enq_req_0_bits_fuOpType; \
        force RTL_PATH.io_enq_req_0_bits_rfWen = U_IF_NAME.io_enq_req_0_bits_rfWen; \
        force RTL_PATH.io_enq_req_0_bits_fpWen = U_IF_NAME.io_enq_req_0_bits_fpWen; \
        force RTL_PATH.io_enq_req_0_bits_vecWen = U_IF_NAME.io_enq_req_0_bits_vecWen; \
        force RTL_PATH.io_enq_req_0_bits_v0Wen = U_IF_NAME.io_enq_req_0_bits_v0Wen; \
        force RTL_PATH.io_enq_req_0_bits_vlWen = U_IF_NAME.io_enq_req_0_bits_vlWen; \
        force RTL_PATH.io_enq_req_0_bits_isXSTrap = U_IF_NAME.io_enq_req_0_bits_isXSTrap; \
        force RTL_PATH.io_enq_req_0_bits_waitForward = U_IF_NAME.io_enq_req_0_bits_waitForward; \
        force RTL_PATH.io_enq_req_0_bits_blockBackward = U_IF_NAME.io_enq_req_0_bits_blockBackward; \
        force RTL_PATH.io_enq_req_0_bits_flushPipe = U_IF_NAME.io_enq_req_0_bits_flushPipe; \
        force RTL_PATH.io_enq_req_0_bits_vpu_vill = U_IF_NAME.io_enq_req_0_bits_vpu_vill; \
        force RTL_PATH.io_enq_req_0_bits_vpu_vma = U_IF_NAME.io_enq_req_0_bits_vpu_vma; \
        force RTL_PATH.io_enq_req_0_bits_vpu_vta = U_IF_NAME.io_enq_req_0_bits_vpu_vta; \
        force RTL_PATH.io_enq_req_0_bits_vpu_vsew = U_IF_NAME.io_enq_req_0_bits_vpu_vsew; \
        force RTL_PATH.io_enq_req_0_bits_vpu_vlmul = U_IF_NAME.io_enq_req_0_bits_vpu_vlmul; \
        force RTL_PATH.io_enq_req_0_bits_vpu_specVill = U_IF_NAME.io_enq_req_0_bits_vpu_specVill; \
        force RTL_PATH.io_enq_req_0_bits_vpu_specVma = U_IF_NAME.io_enq_req_0_bits_vpu_specVma; \
        force RTL_PATH.io_enq_req_0_bits_vpu_specVta = U_IF_NAME.io_enq_req_0_bits_vpu_specVta; \
        force RTL_PATH.io_enq_req_0_bits_vpu_specVsew = U_IF_NAME.io_enq_req_0_bits_vpu_specVsew; \
        force RTL_PATH.io_enq_req_0_bits_vpu_specVlmul = U_IF_NAME.io_enq_req_0_bits_vpu_specVlmul; \
        force RTL_PATH.io_enq_req_0_bits_vlsInstr = U_IF_NAME.io_enq_req_0_bits_vlsInstr; \
        force RTL_PATH.io_enq_req_0_bits_wfflags = U_IF_NAME.io_enq_req_0_bits_wfflags; \
        force RTL_PATH.io_enq_req_0_bits_isMove = U_IF_NAME.io_enq_req_0_bits_isMove; \
        force RTL_PATH.io_enq_req_0_bits_isVset = U_IF_NAME.io_enq_req_0_bits_isVset; \
        force RTL_PATH.io_enq_req_0_bits_firstUop = U_IF_NAME.io_enq_req_0_bits_firstUop; \
        force RTL_PATH.io_enq_req_0_bits_lastUop = U_IF_NAME.io_enq_req_0_bits_lastUop; \
        force RTL_PATH.io_enq_req_0_bits_numWB = U_IF_NAME.io_enq_req_0_bits_numWB; \
        force RTL_PATH.io_enq_req_0_bits_commitType = U_IF_NAME.io_enq_req_0_bits_commitType; \
        force RTL_PATH.io_enq_req_0_bits_pdest = U_IF_NAME.io_enq_req_0_bits_pdest; \
        force RTL_PATH.io_enq_req_0_bits_robIdx_flag = U_IF_NAME.io_enq_req_0_bits_robIdx_flag; \
        force RTL_PATH.io_enq_req_0_bits_robIdx_value = U_IF_NAME.io_enq_req_0_bits_robIdx_value; \
        force RTL_PATH.io_enq_req_0_bits_instrSize = U_IF_NAME.io_enq_req_0_bits_instrSize; \
        force RTL_PATH.io_enq_req_0_bits_dirtyFs = U_IF_NAME.io_enq_req_0_bits_dirtyFs; \
        force RTL_PATH.io_enq_req_0_bits_dirtyVs = U_IF_NAME.io_enq_req_0_bits_dirtyVs; \
        force RTL_PATH.io_enq_req_0_bits_traceBlockInPipe_itype = U_IF_NAME.io_enq_req_0_bits_traceBlockInPipe_itype; \
        force RTL_PATH.io_enq_req_0_bits_traceBlockInPipe_iretire = U_IF_NAME.io_enq_req_0_bits_traceBlockInPipe_iretire; \
        force RTL_PATH.io_enq_req_0_bits_traceBlockInPipe_ilastsize = U_IF_NAME.io_enq_req_0_bits_traceBlockInPipe_ilastsize; \
        force RTL_PATH.io_enq_req_0_bits_eliminatedMove = U_IF_NAME.io_enq_req_0_bits_eliminatedMove; \
        force RTL_PATH.io_enq_req_0_bits_snapshot = U_IF_NAME.io_enq_req_0_bits_snapshot; \
        force RTL_PATH.io_enq_req_0_bits_lqIdx_value = U_IF_NAME.io_enq_req_0_bits_lqIdx_value; \
        force RTL_PATH.io_enq_req_0_bits_sqIdx_value = U_IF_NAME.io_enq_req_0_bits_sqIdx_value; \
        force RTL_PATH.io_enq_req_0_bits_singleStep = U_IF_NAME.io_enq_req_0_bits_singleStep; \
        force RTL_PATH.io_enq_req_0_bits_debug_sim_trig = U_IF_NAME.io_enq_req_0_bits_debug_sim_trig; \
        force RTL_PATH.io_enq_req_1_valid = U_IF_NAME.io_enq_req_1_valid; \
        force RTL_PATH.io_enq_req_1_bits_instr = U_IF_NAME.io_enq_req_1_bits_instr; \
        force RTL_PATH.io_enq_req_1_bits_pc = U_IF_NAME.io_enq_req_1_bits_pc; \
        force RTL_PATH.io_enq_req_1_bits_exceptionVec_0 = U_IF_NAME.io_enq_req_1_bits_exceptionVec_0; \
        force RTL_PATH.io_enq_req_1_bits_exceptionVec_1 = U_IF_NAME.io_enq_req_1_bits_exceptionVec_1; \
        force RTL_PATH.io_enq_req_1_bits_exceptionVec_2 = U_IF_NAME.io_enq_req_1_bits_exceptionVec_2; \
        force RTL_PATH.io_enq_req_1_bits_exceptionVec_3 = U_IF_NAME.io_enq_req_1_bits_exceptionVec_3; \
        force RTL_PATH.io_enq_req_1_bits_exceptionVec_12 = U_IF_NAME.io_enq_req_1_bits_exceptionVec_12; \
        force RTL_PATH.io_enq_req_1_bits_exceptionVec_20 = U_IF_NAME.io_enq_req_1_bits_exceptionVec_20; \
        force RTL_PATH.io_enq_req_1_bits_exceptionVec_22 = U_IF_NAME.io_enq_req_1_bits_exceptionVec_22; \
        force RTL_PATH.io_enq_req_1_bits_isFetchMalAddr = U_IF_NAME.io_enq_req_1_bits_isFetchMalAddr; \
        force RTL_PATH.io_enq_req_1_bits_hasException = U_IF_NAME.io_enq_req_1_bits_hasException; \
        force RTL_PATH.io_enq_req_1_bits_trigger = U_IF_NAME.io_enq_req_1_bits_trigger; \
        force RTL_PATH.io_enq_req_1_bits_preDecodeInfo_isRVC = U_IF_NAME.io_enq_req_1_bits_preDecodeInfo_isRVC; \
        force RTL_PATH.io_enq_req_1_bits_crossPageIPFFix = U_IF_NAME.io_enq_req_1_bits_crossPageIPFFix; \
        force RTL_PATH.io_enq_req_1_bits_ftqPtr_flag = U_IF_NAME.io_enq_req_1_bits_ftqPtr_flag; \
        force RTL_PATH.io_enq_req_1_bits_ftqPtr_value = U_IF_NAME.io_enq_req_1_bits_ftqPtr_value; \
        force RTL_PATH.io_enq_req_1_bits_ftqOffset = U_IF_NAME.io_enq_req_1_bits_ftqOffset; \
        force RTL_PATH.io_enq_req_1_bits_ldest = U_IF_NAME.io_enq_req_1_bits_ldest; \
        force RTL_PATH.io_enq_req_1_bits_fuType = U_IF_NAME.io_enq_req_1_bits_fuType; \
        force RTL_PATH.io_enq_req_1_bits_fuOpType = U_IF_NAME.io_enq_req_1_bits_fuOpType; \
        force RTL_PATH.io_enq_req_1_bits_rfWen = U_IF_NAME.io_enq_req_1_bits_rfWen; \
        force RTL_PATH.io_enq_req_1_bits_fpWen = U_IF_NAME.io_enq_req_1_bits_fpWen; \
        force RTL_PATH.io_enq_req_1_bits_vecWen = U_IF_NAME.io_enq_req_1_bits_vecWen; \
        force RTL_PATH.io_enq_req_1_bits_v0Wen = U_IF_NAME.io_enq_req_1_bits_v0Wen; \
        force RTL_PATH.io_enq_req_1_bits_vlWen = U_IF_NAME.io_enq_req_1_bits_vlWen; \
        force RTL_PATH.io_enq_req_1_bits_isXSTrap = U_IF_NAME.io_enq_req_1_bits_isXSTrap; \
        force RTL_PATH.io_enq_req_1_bits_waitForward = U_IF_NAME.io_enq_req_1_bits_waitForward; \
        force RTL_PATH.io_enq_req_1_bits_blockBackward = U_IF_NAME.io_enq_req_1_bits_blockBackward; \
        force RTL_PATH.io_enq_req_1_bits_flushPipe = U_IF_NAME.io_enq_req_1_bits_flushPipe; \
        force RTL_PATH.io_enq_req_1_bits_vpu_vill = U_IF_NAME.io_enq_req_1_bits_vpu_vill; \
        force RTL_PATH.io_enq_req_1_bits_vpu_vma = U_IF_NAME.io_enq_req_1_bits_vpu_vma; \
        force RTL_PATH.io_enq_req_1_bits_vpu_vta = U_IF_NAME.io_enq_req_1_bits_vpu_vta; \
        force RTL_PATH.io_enq_req_1_bits_vpu_vsew = U_IF_NAME.io_enq_req_1_bits_vpu_vsew; \
        force RTL_PATH.io_enq_req_1_bits_vpu_vlmul = U_IF_NAME.io_enq_req_1_bits_vpu_vlmul; \
        force RTL_PATH.io_enq_req_1_bits_vpu_specVill = U_IF_NAME.io_enq_req_1_bits_vpu_specVill; \
        force RTL_PATH.io_enq_req_1_bits_vpu_specVma = U_IF_NAME.io_enq_req_1_bits_vpu_specVma; \
        force RTL_PATH.io_enq_req_1_bits_vpu_specVta = U_IF_NAME.io_enq_req_1_bits_vpu_specVta; \
        force RTL_PATH.io_enq_req_1_bits_vpu_specVsew = U_IF_NAME.io_enq_req_1_bits_vpu_specVsew; \
        force RTL_PATH.io_enq_req_1_bits_vpu_specVlmul = U_IF_NAME.io_enq_req_1_bits_vpu_specVlmul; \
        force RTL_PATH.io_enq_req_1_bits_vlsInstr = U_IF_NAME.io_enq_req_1_bits_vlsInstr; \
        force RTL_PATH.io_enq_req_1_bits_wfflags = U_IF_NAME.io_enq_req_1_bits_wfflags; \
        force RTL_PATH.io_enq_req_1_bits_isMove = U_IF_NAME.io_enq_req_1_bits_isMove; \
        force RTL_PATH.io_enq_req_1_bits_isVset = U_IF_NAME.io_enq_req_1_bits_isVset; \
        force RTL_PATH.io_enq_req_1_bits_firstUop = U_IF_NAME.io_enq_req_1_bits_firstUop; \
        force RTL_PATH.io_enq_req_1_bits_lastUop = U_IF_NAME.io_enq_req_1_bits_lastUop; \
        force RTL_PATH.io_enq_req_1_bits_numWB = U_IF_NAME.io_enq_req_1_bits_numWB; \
        force RTL_PATH.io_enq_req_1_bits_commitType = U_IF_NAME.io_enq_req_1_bits_commitType; \
        force RTL_PATH.io_enq_req_1_bits_pdest = U_IF_NAME.io_enq_req_1_bits_pdest; \
        force RTL_PATH.io_enq_req_1_bits_robIdx_flag = U_IF_NAME.io_enq_req_1_bits_robIdx_flag; \
        force RTL_PATH.io_enq_req_1_bits_robIdx_value = U_IF_NAME.io_enq_req_1_bits_robIdx_value; \
        force RTL_PATH.io_enq_req_1_bits_instrSize = U_IF_NAME.io_enq_req_1_bits_instrSize; \
        force RTL_PATH.io_enq_req_1_bits_dirtyFs = U_IF_NAME.io_enq_req_1_bits_dirtyFs; \
        force RTL_PATH.io_enq_req_1_bits_dirtyVs = U_IF_NAME.io_enq_req_1_bits_dirtyVs; \
        force RTL_PATH.io_enq_req_1_bits_traceBlockInPipe_itype = U_IF_NAME.io_enq_req_1_bits_traceBlockInPipe_itype; \
        force RTL_PATH.io_enq_req_1_bits_traceBlockInPipe_iretire = U_IF_NAME.io_enq_req_1_bits_traceBlockInPipe_iretire; \
        force RTL_PATH.io_enq_req_1_bits_traceBlockInPipe_ilastsize = U_IF_NAME.io_enq_req_1_bits_traceBlockInPipe_ilastsize; \
        force RTL_PATH.io_enq_req_1_bits_eliminatedMove = U_IF_NAME.io_enq_req_1_bits_eliminatedMove; \
        force RTL_PATH.io_enq_req_1_bits_snapshot = U_IF_NAME.io_enq_req_1_bits_snapshot; \
        force RTL_PATH.io_enq_req_1_bits_lqIdx_value = U_IF_NAME.io_enq_req_1_bits_lqIdx_value; \
        force RTL_PATH.io_enq_req_1_bits_sqIdx_value = U_IF_NAME.io_enq_req_1_bits_sqIdx_value; \
        force RTL_PATH.io_enq_req_1_bits_singleStep = U_IF_NAME.io_enq_req_1_bits_singleStep; \
        force RTL_PATH.io_enq_req_1_bits_debug_sim_trig = U_IF_NAME.io_enq_req_1_bits_debug_sim_trig; \
        force RTL_PATH.io_enq_req_2_valid = U_IF_NAME.io_enq_req_2_valid; \
        force RTL_PATH.io_enq_req_2_bits_instr = U_IF_NAME.io_enq_req_2_bits_instr; \
        force RTL_PATH.io_enq_req_2_bits_pc = U_IF_NAME.io_enq_req_2_bits_pc; \
        force RTL_PATH.io_enq_req_2_bits_exceptionVec_0 = U_IF_NAME.io_enq_req_2_bits_exceptionVec_0; \
        force RTL_PATH.io_enq_req_2_bits_exceptionVec_1 = U_IF_NAME.io_enq_req_2_bits_exceptionVec_1; \
        force RTL_PATH.io_enq_req_2_bits_exceptionVec_2 = U_IF_NAME.io_enq_req_2_bits_exceptionVec_2; \
        force RTL_PATH.io_enq_req_2_bits_exceptionVec_3 = U_IF_NAME.io_enq_req_2_bits_exceptionVec_3; \
        force RTL_PATH.io_enq_req_2_bits_exceptionVec_12 = U_IF_NAME.io_enq_req_2_bits_exceptionVec_12; \
        force RTL_PATH.io_enq_req_2_bits_exceptionVec_20 = U_IF_NAME.io_enq_req_2_bits_exceptionVec_20; \
        force RTL_PATH.io_enq_req_2_bits_exceptionVec_22 = U_IF_NAME.io_enq_req_2_bits_exceptionVec_22; \
        force RTL_PATH.io_enq_req_2_bits_isFetchMalAddr = U_IF_NAME.io_enq_req_2_bits_isFetchMalAddr; \
        force RTL_PATH.io_enq_req_2_bits_hasException = U_IF_NAME.io_enq_req_2_bits_hasException; \
        force RTL_PATH.io_enq_req_2_bits_trigger = U_IF_NAME.io_enq_req_2_bits_trigger; \
        force RTL_PATH.io_enq_req_2_bits_preDecodeInfo_isRVC = U_IF_NAME.io_enq_req_2_bits_preDecodeInfo_isRVC; \
        force RTL_PATH.io_enq_req_2_bits_crossPageIPFFix = U_IF_NAME.io_enq_req_2_bits_crossPageIPFFix; \
        force RTL_PATH.io_enq_req_2_bits_ftqPtr_flag = U_IF_NAME.io_enq_req_2_bits_ftqPtr_flag; \
        force RTL_PATH.io_enq_req_2_bits_ftqPtr_value = U_IF_NAME.io_enq_req_2_bits_ftqPtr_value; \
        force RTL_PATH.io_enq_req_2_bits_ftqOffset = U_IF_NAME.io_enq_req_2_bits_ftqOffset; \
        force RTL_PATH.io_enq_req_2_bits_ldest = U_IF_NAME.io_enq_req_2_bits_ldest; \
        force RTL_PATH.io_enq_req_2_bits_fuType = U_IF_NAME.io_enq_req_2_bits_fuType; \
        force RTL_PATH.io_enq_req_2_bits_fuOpType = U_IF_NAME.io_enq_req_2_bits_fuOpType; \
        force RTL_PATH.io_enq_req_2_bits_rfWen = U_IF_NAME.io_enq_req_2_bits_rfWen; \
        force RTL_PATH.io_enq_req_2_bits_fpWen = U_IF_NAME.io_enq_req_2_bits_fpWen; \
        force RTL_PATH.io_enq_req_2_bits_vecWen = U_IF_NAME.io_enq_req_2_bits_vecWen; \
        force RTL_PATH.io_enq_req_2_bits_v0Wen = U_IF_NAME.io_enq_req_2_bits_v0Wen; \
        force RTL_PATH.io_enq_req_2_bits_vlWen = U_IF_NAME.io_enq_req_2_bits_vlWen; \
        force RTL_PATH.io_enq_req_2_bits_isXSTrap = U_IF_NAME.io_enq_req_2_bits_isXSTrap; \
        force RTL_PATH.io_enq_req_2_bits_waitForward = U_IF_NAME.io_enq_req_2_bits_waitForward; \
        force RTL_PATH.io_enq_req_2_bits_blockBackward = U_IF_NAME.io_enq_req_2_bits_blockBackward; \
        force RTL_PATH.io_enq_req_2_bits_flushPipe = U_IF_NAME.io_enq_req_2_bits_flushPipe; \
        force RTL_PATH.io_enq_req_2_bits_vpu_vill = U_IF_NAME.io_enq_req_2_bits_vpu_vill; \
        force RTL_PATH.io_enq_req_2_bits_vpu_vma = U_IF_NAME.io_enq_req_2_bits_vpu_vma; \
        force RTL_PATH.io_enq_req_2_bits_vpu_vta = U_IF_NAME.io_enq_req_2_bits_vpu_vta; \
        force RTL_PATH.io_enq_req_2_bits_vpu_vsew = U_IF_NAME.io_enq_req_2_bits_vpu_vsew; \
        force RTL_PATH.io_enq_req_2_bits_vpu_vlmul = U_IF_NAME.io_enq_req_2_bits_vpu_vlmul; \
        force RTL_PATH.io_enq_req_2_bits_vpu_specVill = U_IF_NAME.io_enq_req_2_bits_vpu_specVill; \
        force RTL_PATH.io_enq_req_2_bits_vpu_specVma = U_IF_NAME.io_enq_req_2_bits_vpu_specVma; \
        force RTL_PATH.io_enq_req_2_bits_vpu_specVta = U_IF_NAME.io_enq_req_2_bits_vpu_specVta; \
        force RTL_PATH.io_enq_req_2_bits_vpu_specVsew = U_IF_NAME.io_enq_req_2_bits_vpu_specVsew; \
        force RTL_PATH.io_enq_req_2_bits_vpu_specVlmul = U_IF_NAME.io_enq_req_2_bits_vpu_specVlmul; \
        force RTL_PATH.io_enq_req_2_bits_vlsInstr = U_IF_NAME.io_enq_req_2_bits_vlsInstr; \
        force RTL_PATH.io_enq_req_2_bits_wfflags = U_IF_NAME.io_enq_req_2_bits_wfflags; \
        force RTL_PATH.io_enq_req_2_bits_isMove = U_IF_NAME.io_enq_req_2_bits_isMove; \
        force RTL_PATH.io_enq_req_2_bits_isVset = U_IF_NAME.io_enq_req_2_bits_isVset; \
        force RTL_PATH.io_enq_req_2_bits_firstUop = U_IF_NAME.io_enq_req_2_bits_firstUop; \
        force RTL_PATH.io_enq_req_2_bits_lastUop = U_IF_NAME.io_enq_req_2_bits_lastUop; \
        force RTL_PATH.io_enq_req_2_bits_numWB = U_IF_NAME.io_enq_req_2_bits_numWB; \
        force RTL_PATH.io_enq_req_2_bits_commitType = U_IF_NAME.io_enq_req_2_bits_commitType; \
        force RTL_PATH.io_enq_req_2_bits_pdest = U_IF_NAME.io_enq_req_2_bits_pdest; \
        force RTL_PATH.io_enq_req_2_bits_robIdx_flag = U_IF_NAME.io_enq_req_2_bits_robIdx_flag; \
        force RTL_PATH.io_enq_req_2_bits_robIdx_value = U_IF_NAME.io_enq_req_2_bits_robIdx_value; \
        force RTL_PATH.io_enq_req_2_bits_instrSize = U_IF_NAME.io_enq_req_2_bits_instrSize; \
        force RTL_PATH.io_enq_req_2_bits_dirtyFs = U_IF_NAME.io_enq_req_2_bits_dirtyFs; \
        force RTL_PATH.io_enq_req_2_bits_dirtyVs = U_IF_NAME.io_enq_req_2_bits_dirtyVs; \
        force RTL_PATH.io_enq_req_2_bits_traceBlockInPipe_itype = U_IF_NAME.io_enq_req_2_bits_traceBlockInPipe_itype; \
        force RTL_PATH.io_enq_req_2_bits_traceBlockInPipe_iretire = U_IF_NAME.io_enq_req_2_bits_traceBlockInPipe_iretire; \
        force RTL_PATH.io_enq_req_2_bits_traceBlockInPipe_ilastsize = U_IF_NAME.io_enq_req_2_bits_traceBlockInPipe_ilastsize; \
        force RTL_PATH.io_enq_req_2_bits_eliminatedMove = U_IF_NAME.io_enq_req_2_bits_eliminatedMove; \
        force RTL_PATH.io_enq_req_2_bits_snapshot = U_IF_NAME.io_enq_req_2_bits_snapshot; \
        force RTL_PATH.io_enq_req_2_bits_lqIdx_value = U_IF_NAME.io_enq_req_2_bits_lqIdx_value; \
        force RTL_PATH.io_enq_req_2_bits_sqIdx_value = U_IF_NAME.io_enq_req_2_bits_sqIdx_value; \
        force RTL_PATH.io_enq_req_2_bits_singleStep = U_IF_NAME.io_enq_req_2_bits_singleStep; \
        force RTL_PATH.io_enq_req_2_bits_debug_sim_trig = U_IF_NAME.io_enq_req_2_bits_debug_sim_trig; \
        force RTL_PATH.io_enq_req_3_valid = U_IF_NAME.io_enq_req_3_valid; \
        force RTL_PATH.io_enq_req_3_bits_instr = U_IF_NAME.io_enq_req_3_bits_instr; \
        force RTL_PATH.io_enq_req_3_bits_pc = U_IF_NAME.io_enq_req_3_bits_pc; \
        force RTL_PATH.io_enq_req_3_bits_exceptionVec_0 = U_IF_NAME.io_enq_req_3_bits_exceptionVec_0; \
        force RTL_PATH.io_enq_req_3_bits_exceptionVec_1 = U_IF_NAME.io_enq_req_3_bits_exceptionVec_1; \
        force RTL_PATH.io_enq_req_3_bits_exceptionVec_2 = U_IF_NAME.io_enq_req_3_bits_exceptionVec_2; \
        force RTL_PATH.io_enq_req_3_bits_exceptionVec_3 = U_IF_NAME.io_enq_req_3_bits_exceptionVec_3; \
        force RTL_PATH.io_enq_req_3_bits_exceptionVec_12 = U_IF_NAME.io_enq_req_3_bits_exceptionVec_12; \
        force RTL_PATH.io_enq_req_3_bits_exceptionVec_20 = U_IF_NAME.io_enq_req_3_bits_exceptionVec_20; \
        force RTL_PATH.io_enq_req_3_bits_exceptionVec_22 = U_IF_NAME.io_enq_req_3_bits_exceptionVec_22; \
        force RTL_PATH.io_enq_req_3_bits_isFetchMalAddr = U_IF_NAME.io_enq_req_3_bits_isFetchMalAddr; \
        force RTL_PATH.io_enq_req_3_bits_hasException = U_IF_NAME.io_enq_req_3_bits_hasException; \
        force RTL_PATH.io_enq_req_3_bits_trigger = U_IF_NAME.io_enq_req_3_bits_trigger; \
        force RTL_PATH.io_enq_req_3_bits_preDecodeInfo_isRVC = U_IF_NAME.io_enq_req_3_bits_preDecodeInfo_isRVC; \
        force RTL_PATH.io_enq_req_3_bits_crossPageIPFFix = U_IF_NAME.io_enq_req_3_bits_crossPageIPFFix; \
        force RTL_PATH.io_enq_req_3_bits_ftqPtr_flag = U_IF_NAME.io_enq_req_3_bits_ftqPtr_flag; \
        force RTL_PATH.io_enq_req_3_bits_ftqPtr_value = U_IF_NAME.io_enq_req_3_bits_ftqPtr_value; \
        force RTL_PATH.io_enq_req_3_bits_ftqOffset = U_IF_NAME.io_enq_req_3_bits_ftqOffset; \
        force RTL_PATH.io_enq_req_3_bits_ldest = U_IF_NAME.io_enq_req_3_bits_ldest; \
        force RTL_PATH.io_enq_req_3_bits_fuType = U_IF_NAME.io_enq_req_3_bits_fuType; \
        force RTL_PATH.io_enq_req_3_bits_fuOpType = U_IF_NAME.io_enq_req_3_bits_fuOpType; \
        force RTL_PATH.io_enq_req_3_bits_rfWen = U_IF_NAME.io_enq_req_3_bits_rfWen; \
        force RTL_PATH.io_enq_req_3_bits_fpWen = U_IF_NAME.io_enq_req_3_bits_fpWen; \
        force RTL_PATH.io_enq_req_3_bits_vecWen = U_IF_NAME.io_enq_req_3_bits_vecWen; \
        force RTL_PATH.io_enq_req_3_bits_v0Wen = U_IF_NAME.io_enq_req_3_bits_v0Wen; \
        force RTL_PATH.io_enq_req_3_bits_vlWen = U_IF_NAME.io_enq_req_3_bits_vlWen; \
        force RTL_PATH.io_enq_req_3_bits_isXSTrap = U_IF_NAME.io_enq_req_3_bits_isXSTrap; \
        force RTL_PATH.io_enq_req_3_bits_waitForward = U_IF_NAME.io_enq_req_3_bits_waitForward; \
        force RTL_PATH.io_enq_req_3_bits_blockBackward = U_IF_NAME.io_enq_req_3_bits_blockBackward; \
        force RTL_PATH.io_enq_req_3_bits_flushPipe = U_IF_NAME.io_enq_req_3_bits_flushPipe; \
        force RTL_PATH.io_enq_req_3_bits_vpu_vill = U_IF_NAME.io_enq_req_3_bits_vpu_vill; \
        force RTL_PATH.io_enq_req_3_bits_vpu_vma = U_IF_NAME.io_enq_req_3_bits_vpu_vma; \
        force RTL_PATH.io_enq_req_3_bits_vpu_vta = U_IF_NAME.io_enq_req_3_bits_vpu_vta; \
        force RTL_PATH.io_enq_req_3_bits_vpu_vsew = U_IF_NAME.io_enq_req_3_bits_vpu_vsew; \
        force RTL_PATH.io_enq_req_3_bits_vpu_vlmul = U_IF_NAME.io_enq_req_3_bits_vpu_vlmul; \
        force RTL_PATH.io_enq_req_3_bits_vpu_specVill = U_IF_NAME.io_enq_req_3_bits_vpu_specVill; \
        force RTL_PATH.io_enq_req_3_bits_vpu_specVma = U_IF_NAME.io_enq_req_3_bits_vpu_specVma; \
        force RTL_PATH.io_enq_req_3_bits_vpu_specVta = U_IF_NAME.io_enq_req_3_bits_vpu_specVta; \
        force RTL_PATH.io_enq_req_3_bits_vpu_specVsew = U_IF_NAME.io_enq_req_3_bits_vpu_specVsew; \
        force RTL_PATH.io_enq_req_3_bits_vpu_specVlmul = U_IF_NAME.io_enq_req_3_bits_vpu_specVlmul; \
        force RTL_PATH.io_enq_req_3_bits_vlsInstr = U_IF_NAME.io_enq_req_3_bits_vlsInstr; \
        force RTL_PATH.io_enq_req_3_bits_wfflags = U_IF_NAME.io_enq_req_3_bits_wfflags; \
        force RTL_PATH.io_enq_req_3_bits_isMove = U_IF_NAME.io_enq_req_3_bits_isMove; \
        force RTL_PATH.io_enq_req_3_bits_isVset = U_IF_NAME.io_enq_req_3_bits_isVset; \
        force RTL_PATH.io_enq_req_3_bits_firstUop = U_IF_NAME.io_enq_req_3_bits_firstUop; \
        force RTL_PATH.io_enq_req_3_bits_lastUop = U_IF_NAME.io_enq_req_3_bits_lastUop; \
        force RTL_PATH.io_enq_req_3_bits_numWB = U_IF_NAME.io_enq_req_3_bits_numWB; \
        force RTL_PATH.io_enq_req_3_bits_commitType = U_IF_NAME.io_enq_req_3_bits_commitType; \
        force RTL_PATH.io_enq_req_3_bits_pdest = U_IF_NAME.io_enq_req_3_bits_pdest; \
        force RTL_PATH.io_enq_req_3_bits_robIdx_flag = U_IF_NAME.io_enq_req_3_bits_robIdx_flag; \
        force RTL_PATH.io_enq_req_3_bits_robIdx_value = U_IF_NAME.io_enq_req_3_bits_robIdx_value; \
        force RTL_PATH.io_enq_req_3_bits_instrSize = U_IF_NAME.io_enq_req_3_bits_instrSize; \
        force RTL_PATH.io_enq_req_3_bits_dirtyFs = U_IF_NAME.io_enq_req_3_bits_dirtyFs; \
        force RTL_PATH.io_enq_req_3_bits_dirtyVs = U_IF_NAME.io_enq_req_3_bits_dirtyVs; \
        force RTL_PATH.io_enq_req_3_bits_traceBlockInPipe_itype = U_IF_NAME.io_enq_req_3_bits_traceBlockInPipe_itype; \
        force RTL_PATH.io_enq_req_3_bits_traceBlockInPipe_iretire = U_IF_NAME.io_enq_req_3_bits_traceBlockInPipe_iretire; \
        force RTL_PATH.io_enq_req_3_bits_traceBlockInPipe_ilastsize = U_IF_NAME.io_enq_req_3_bits_traceBlockInPipe_ilastsize; \
        force RTL_PATH.io_enq_req_3_bits_eliminatedMove = U_IF_NAME.io_enq_req_3_bits_eliminatedMove; \
        force RTL_PATH.io_enq_req_3_bits_snapshot = U_IF_NAME.io_enq_req_3_bits_snapshot; \
        force RTL_PATH.io_enq_req_3_bits_lqIdx_value = U_IF_NAME.io_enq_req_3_bits_lqIdx_value; \
        force RTL_PATH.io_enq_req_3_bits_sqIdx_value = U_IF_NAME.io_enq_req_3_bits_sqIdx_value; \
        force RTL_PATH.io_enq_req_3_bits_singleStep = U_IF_NAME.io_enq_req_3_bits_singleStep; \
        force RTL_PATH.io_enq_req_3_bits_debug_sim_trig = U_IF_NAME.io_enq_req_3_bits_debug_sim_trig; \
        force RTL_PATH.io_enq_req_4_valid = U_IF_NAME.io_enq_req_4_valid; \
        force RTL_PATH.io_enq_req_4_bits_instr = U_IF_NAME.io_enq_req_4_bits_instr; \
        force RTL_PATH.io_enq_req_4_bits_pc = U_IF_NAME.io_enq_req_4_bits_pc; \
        force RTL_PATH.io_enq_req_4_bits_exceptionVec_0 = U_IF_NAME.io_enq_req_4_bits_exceptionVec_0; \
        force RTL_PATH.io_enq_req_4_bits_exceptionVec_1 = U_IF_NAME.io_enq_req_4_bits_exceptionVec_1; \
        force RTL_PATH.io_enq_req_4_bits_exceptionVec_2 = U_IF_NAME.io_enq_req_4_bits_exceptionVec_2; \
        force RTL_PATH.io_enq_req_4_bits_exceptionVec_3 = U_IF_NAME.io_enq_req_4_bits_exceptionVec_3; \
        force RTL_PATH.io_enq_req_4_bits_exceptionVec_12 = U_IF_NAME.io_enq_req_4_bits_exceptionVec_12; \
        force RTL_PATH.io_enq_req_4_bits_exceptionVec_20 = U_IF_NAME.io_enq_req_4_bits_exceptionVec_20; \
        force RTL_PATH.io_enq_req_4_bits_exceptionVec_22 = U_IF_NAME.io_enq_req_4_bits_exceptionVec_22; \
        force RTL_PATH.io_enq_req_4_bits_isFetchMalAddr = U_IF_NAME.io_enq_req_4_bits_isFetchMalAddr; \
        force RTL_PATH.io_enq_req_4_bits_hasException = U_IF_NAME.io_enq_req_4_bits_hasException; \
        force RTL_PATH.io_enq_req_4_bits_trigger = U_IF_NAME.io_enq_req_4_bits_trigger; \
        force RTL_PATH.io_enq_req_4_bits_preDecodeInfo_isRVC = U_IF_NAME.io_enq_req_4_bits_preDecodeInfo_isRVC; \
        force RTL_PATH.io_enq_req_4_bits_crossPageIPFFix = U_IF_NAME.io_enq_req_4_bits_crossPageIPFFix; \
        force RTL_PATH.io_enq_req_4_bits_ftqPtr_flag = U_IF_NAME.io_enq_req_4_bits_ftqPtr_flag; \
        force RTL_PATH.io_enq_req_4_bits_ftqPtr_value = U_IF_NAME.io_enq_req_4_bits_ftqPtr_value; \
        force RTL_PATH.io_enq_req_4_bits_ftqOffset = U_IF_NAME.io_enq_req_4_bits_ftqOffset; \
        force RTL_PATH.io_enq_req_4_bits_ldest = U_IF_NAME.io_enq_req_4_bits_ldest; \
        force RTL_PATH.io_enq_req_4_bits_fuType = U_IF_NAME.io_enq_req_4_bits_fuType; \
        force RTL_PATH.io_enq_req_4_bits_fuOpType = U_IF_NAME.io_enq_req_4_bits_fuOpType; \
        force RTL_PATH.io_enq_req_4_bits_rfWen = U_IF_NAME.io_enq_req_4_bits_rfWen; \
        force RTL_PATH.io_enq_req_4_bits_fpWen = U_IF_NAME.io_enq_req_4_bits_fpWen; \
        force RTL_PATH.io_enq_req_4_bits_vecWen = U_IF_NAME.io_enq_req_4_bits_vecWen; \
        force RTL_PATH.io_enq_req_4_bits_v0Wen = U_IF_NAME.io_enq_req_4_bits_v0Wen; \
        force RTL_PATH.io_enq_req_4_bits_vlWen = U_IF_NAME.io_enq_req_4_bits_vlWen; \
        force RTL_PATH.io_enq_req_4_bits_isXSTrap = U_IF_NAME.io_enq_req_4_bits_isXSTrap; \
        force RTL_PATH.io_enq_req_4_bits_waitForward = U_IF_NAME.io_enq_req_4_bits_waitForward; \
        force RTL_PATH.io_enq_req_4_bits_blockBackward = U_IF_NAME.io_enq_req_4_bits_blockBackward; \
        force RTL_PATH.io_enq_req_4_bits_flushPipe = U_IF_NAME.io_enq_req_4_bits_flushPipe; \
        force RTL_PATH.io_enq_req_4_bits_vpu_vill = U_IF_NAME.io_enq_req_4_bits_vpu_vill; \
        force RTL_PATH.io_enq_req_4_bits_vpu_vma = U_IF_NAME.io_enq_req_4_bits_vpu_vma; \
        force RTL_PATH.io_enq_req_4_bits_vpu_vta = U_IF_NAME.io_enq_req_4_bits_vpu_vta; \
        force RTL_PATH.io_enq_req_4_bits_vpu_vsew = U_IF_NAME.io_enq_req_4_bits_vpu_vsew; \
        force RTL_PATH.io_enq_req_4_bits_vpu_vlmul = U_IF_NAME.io_enq_req_4_bits_vpu_vlmul; \
        force RTL_PATH.io_enq_req_4_bits_vpu_specVill = U_IF_NAME.io_enq_req_4_bits_vpu_specVill; \
        force RTL_PATH.io_enq_req_4_bits_vpu_specVma = U_IF_NAME.io_enq_req_4_bits_vpu_specVma; \
        force RTL_PATH.io_enq_req_4_bits_vpu_specVta = U_IF_NAME.io_enq_req_4_bits_vpu_specVta; \
        force RTL_PATH.io_enq_req_4_bits_vpu_specVsew = U_IF_NAME.io_enq_req_4_bits_vpu_specVsew; \
        force RTL_PATH.io_enq_req_4_bits_vpu_specVlmul = U_IF_NAME.io_enq_req_4_bits_vpu_specVlmul; \
        force RTL_PATH.io_enq_req_4_bits_vlsInstr = U_IF_NAME.io_enq_req_4_bits_vlsInstr; \
        force RTL_PATH.io_enq_req_4_bits_wfflags = U_IF_NAME.io_enq_req_4_bits_wfflags; \
        force RTL_PATH.io_enq_req_4_bits_isMove = U_IF_NAME.io_enq_req_4_bits_isMove; \
        force RTL_PATH.io_enq_req_4_bits_isVset = U_IF_NAME.io_enq_req_4_bits_isVset; \
        force RTL_PATH.io_enq_req_4_bits_firstUop = U_IF_NAME.io_enq_req_4_bits_firstUop; \
        force RTL_PATH.io_enq_req_4_bits_lastUop = U_IF_NAME.io_enq_req_4_bits_lastUop; \
        force RTL_PATH.io_enq_req_4_bits_numWB = U_IF_NAME.io_enq_req_4_bits_numWB; \
        force RTL_PATH.io_enq_req_4_bits_commitType = U_IF_NAME.io_enq_req_4_bits_commitType; \
        force RTL_PATH.io_enq_req_4_bits_pdest = U_IF_NAME.io_enq_req_4_bits_pdest; \
        force RTL_PATH.io_enq_req_4_bits_robIdx_flag = U_IF_NAME.io_enq_req_4_bits_robIdx_flag; \
        force RTL_PATH.io_enq_req_4_bits_robIdx_value = U_IF_NAME.io_enq_req_4_bits_robIdx_value; \
        force RTL_PATH.io_enq_req_4_bits_instrSize = U_IF_NAME.io_enq_req_4_bits_instrSize; \
        force RTL_PATH.io_enq_req_4_bits_dirtyFs = U_IF_NAME.io_enq_req_4_bits_dirtyFs; \
        force RTL_PATH.io_enq_req_4_bits_dirtyVs = U_IF_NAME.io_enq_req_4_bits_dirtyVs; \
        force RTL_PATH.io_enq_req_4_bits_traceBlockInPipe_itype = U_IF_NAME.io_enq_req_4_bits_traceBlockInPipe_itype; \
        force RTL_PATH.io_enq_req_4_bits_traceBlockInPipe_iretire = U_IF_NAME.io_enq_req_4_bits_traceBlockInPipe_iretire; \
        force RTL_PATH.io_enq_req_4_bits_traceBlockInPipe_ilastsize = U_IF_NAME.io_enq_req_4_bits_traceBlockInPipe_ilastsize; \
        force RTL_PATH.io_enq_req_4_bits_eliminatedMove = U_IF_NAME.io_enq_req_4_bits_eliminatedMove; \
        force RTL_PATH.io_enq_req_4_bits_snapshot = U_IF_NAME.io_enq_req_4_bits_snapshot; \
        force RTL_PATH.io_enq_req_4_bits_lqIdx_value = U_IF_NAME.io_enq_req_4_bits_lqIdx_value; \
        force RTL_PATH.io_enq_req_4_bits_sqIdx_value = U_IF_NAME.io_enq_req_4_bits_sqIdx_value; \
        force RTL_PATH.io_enq_req_4_bits_singleStep = U_IF_NAME.io_enq_req_4_bits_singleStep; \
        force RTL_PATH.io_enq_req_4_bits_debug_sim_trig = U_IF_NAME.io_enq_req_4_bits_debug_sim_trig; \
        force RTL_PATH.io_enq_req_5_valid = U_IF_NAME.io_enq_req_5_valid; \
        force RTL_PATH.io_enq_req_5_bits_instr = U_IF_NAME.io_enq_req_5_bits_instr; \
        force RTL_PATH.io_enq_req_5_bits_pc = U_IF_NAME.io_enq_req_5_bits_pc; \
        force RTL_PATH.io_enq_req_5_bits_exceptionVec_0 = U_IF_NAME.io_enq_req_5_bits_exceptionVec_0; \
        force RTL_PATH.io_enq_req_5_bits_exceptionVec_1 = U_IF_NAME.io_enq_req_5_bits_exceptionVec_1; \
        force RTL_PATH.io_enq_req_5_bits_exceptionVec_2 = U_IF_NAME.io_enq_req_5_bits_exceptionVec_2; \
        force RTL_PATH.io_enq_req_5_bits_exceptionVec_3 = U_IF_NAME.io_enq_req_5_bits_exceptionVec_3; \
        force RTL_PATH.io_enq_req_5_bits_exceptionVec_12 = U_IF_NAME.io_enq_req_5_bits_exceptionVec_12; \
        force RTL_PATH.io_enq_req_5_bits_exceptionVec_20 = U_IF_NAME.io_enq_req_5_bits_exceptionVec_20; \
        force RTL_PATH.io_enq_req_5_bits_exceptionVec_22 = U_IF_NAME.io_enq_req_5_bits_exceptionVec_22; \
        force RTL_PATH.io_enq_req_5_bits_isFetchMalAddr = U_IF_NAME.io_enq_req_5_bits_isFetchMalAddr; \
        force RTL_PATH.io_enq_req_5_bits_hasException = U_IF_NAME.io_enq_req_5_bits_hasException; \
        force RTL_PATH.io_enq_req_5_bits_trigger = U_IF_NAME.io_enq_req_5_bits_trigger; \
        force RTL_PATH.io_enq_req_5_bits_preDecodeInfo_isRVC = U_IF_NAME.io_enq_req_5_bits_preDecodeInfo_isRVC; \
        force RTL_PATH.io_enq_req_5_bits_crossPageIPFFix = U_IF_NAME.io_enq_req_5_bits_crossPageIPFFix; \
        force RTL_PATH.io_enq_req_5_bits_ftqPtr_flag = U_IF_NAME.io_enq_req_5_bits_ftqPtr_flag; \
        force RTL_PATH.io_enq_req_5_bits_ftqPtr_value = U_IF_NAME.io_enq_req_5_bits_ftqPtr_value; \
        force RTL_PATH.io_enq_req_5_bits_ftqOffset = U_IF_NAME.io_enq_req_5_bits_ftqOffset; \
        force RTL_PATH.io_enq_req_5_bits_ldest = U_IF_NAME.io_enq_req_5_bits_ldest; \
        force RTL_PATH.io_enq_req_5_bits_fuType = U_IF_NAME.io_enq_req_5_bits_fuType; \
        force RTL_PATH.io_enq_req_5_bits_fuOpType = U_IF_NAME.io_enq_req_5_bits_fuOpType; \
        force RTL_PATH.io_enq_req_5_bits_rfWen = U_IF_NAME.io_enq_req_5_bits_rfWen; \
        force RTL_PATH.io_enq_req_5_bits_fpWen = U_IF_NAME.io_enq_req_5_bits_fpWen; \
        force RTL_PATH.io_enq_req_5_bits_vecWen = U_IF_NAME.io_enq_req_5_bits_vecWen; \
        force RTL_PATH.io_enq_req_5_bits_v0Wen = U_IF_NAME.io_enq_req_5_bits_v0Wen; \
        force RTL_PATH.io_enq_req_5_bits_vlWen = U_IF_NAME.io_enq_req_5_bits_vlWen; \
        force RTL_PATH.io_enq_req_5_bits_isXSTrap = U_IF_NAME.io_enq_req_5_bits_isXSTrap; \
        force RTL_PATH.io_enq_req_5_bits_waitForward = U_IF_NAME.io_enq_req_5_bits_waitForward; \
        force RTL_PATH.io_enq_req_5_bits_blockBackward = U_IF_NAME.io_enq_req_5_bits_blockBackward; \
        force RTL_PATH.io_enq_req_5_bits_flushPipe = U_IF_NAME.io_enq_req_5_bits_flushPipe; \
        force RTL_PATH.io_enq_req_5_bits_vpu_vill = U_IF_NAME.io_enq_req_5_bits_vpu_vill; \
        force RTL_PATH.io_enq_req_5_bits_vpu_vma = U_IF_NAME.io_enq_req_5_bits_vpu_vma; \
        force RTL_PATH.io_enq_req_5_bits_vpu_vta = U_IF_NAME.io_enq_req_5_bits_vpu_vta; \
        force RTL_PATH.io_enq_req_5_bits_vpu_vsew = U_IF_NAME.io_enq_req_5_bits_vpu_vsew; \
        force RTL_PATH.io_enq_req_5_bits_vpu_vlmul = U_IF_NAME.io_enq_req_5_bits_vpu_vlmul; \
        force RTL_PATH.io_enq_req_5_bits_vpu_specVill = U_IF_NAME.io_enq_req_5_bits_vpu_specVill; \
        force RTL_PATH.io_enq_req_5_bits_vpu_specVma = U_IF_NAME.io_enq_req_5_bits_vpu_specVma; \
        force RTL_PATH.io_enq_req_5_bits_vpu_specVta = U_IF_NAME.io_enq_req_5_bits_vpu_specVta; \
        force RTL_PATH.io_enq_req_5_bits_vpu_specVsew = U_IF_NAME.io_enq_req_5_bits_vpu_specVsew; \
        force RTL_PATH.io_enq_req_5_bits_vpu_specVlmul = U_IF_NAME.io_enq_req_5_bits_vpu_specVlmul; \
        force RTL_PATH.io_enq_req_5_bits_vlsInstr = U_IF_NAME.io_enq_req_5_bits_vlsInstr; \
        force RTL_PATH.io_enq_req_5_bits_wfflags = U_IF_NAME.io_enq_req_5_bits_wfflags; \
        force RTL_PATH.io_enq_req_5_bits_isMove = U_IF_NAME.io_enq_req_5_bits_isMove; \
        force RTL_PATH.io_enq_req_5_bits_isVset = U_IF_NAME.io_enq_req_5_bits_isVset; \
        force RTL_PATH.io_enq_req_5_bits_firstUop = U_IF_NAME.io_enq_req_5_bits_firstUop; \
        force RTL_PATH.io_enq_req_5_bits_lastUop = U_IF_NAME.io_enq_req_5_bits_lastUop; \
        force RTL_PATH.io_enq_req_5_bits_numWB = U_IF_NAME.io_enq_req_5_bits_numWB; \
        force RTL_PATH.io_enq_req_5_bits_commitType = U_IF_NAME.io_enq_req_5_bits_commitType; \
        force RTL_PATH.io_enq_req_5_bits_pdest = U_IF_NAME.io_enq_req_5_bits_pdest; \
        force RTL_PATH.io_enq_req_5_bits_robIdx_flag = U_IF_NAME.io_enq_req_5_bits_robIdx_flag; \
        force RTL_PATH.io_enq_req_5_bits_robIdx_value = U_IF_NAME.io_enq_req_5_bits_robIdx_value; \
        force RTL_PATH.io_enq_req_5_bits_instrSize = U_IF_NAME.io_enq_req_5_bits_instrSize; \
        force RTL_PATH.io_enq_req_5_bits_dirtyFs = U_IF_NAME.io_enq_req_5_bits_dirtyFs; \
        force RTL_PATH.io_enq_req_5_bits_dirtyVs = U_IF_NAME.io_enq_req_5_bits_dirtyVs; \
        force RTL_PATH.io_enq_req_5_bits_traceBlockInPipe_itype = U_IF_NAME.io_enq_req_5_bits_traceBlockInPipe_itype; \
        force RTL_PATH.io_enq_req_5_bits_traceBlockInPipe_iretire = U_IF_NAME.io_enq_req_5_bits_traceBlockInPipe_iretire; \
        force RTL_PATH.io_enq_req_5_bits_traceBlockInPipe_ilastsize = U_IF_NAME.io_enq_req_5_bits_traceBlockInPipe_ilastsize; \
        force RTL_PATH.io_enq_req_5_bits_eliminatedMove = U_IF_NAME.io_enq_req_5_bits_eliminatedMove; \
        force RTL_PATH.io_enq_req_5_bits_snapshot = U_IF_NAME.io_enq_req_5_bits_snapshot; \
        force RTL_PATH.io_enq_req_5_bits_lqIdx_value = U_IF_NAME.io_enq_req_5_bits_lqIdx_value; \
        force RTL_PATH.io_enq_req_5_bits_sqIdx_value = U_IF_NAME.io_enq_req_5_bits_sqIdx_value; \
        force RTL_PATH.io_enq_req_5_bits_singleStep = U_IF_NAME.io_enq_req_5_bits_singleStep; \
        force RTL_PATH.io_enq_req_5_bits_debug_sim_trig = U_IF_NAME.io_enq_req_5_bits_debug_sim_trig; \
    end \
    `else \
    initial begin \
        force U_IF_NAME.clock = RTL_PATH.clock; \
        force U_IF_NAME.reset = RTL_PATH.reset; \
        force U_IF_NAME.io_hartId = RTL_PATH.io_hartId; \
        force U_IF_NAME.io_enq_req_0_valid = RTL_PATH.io_enq_req_0_valid; \
        force U_IF_NAME.io_enq_req_0_bits_instr = RTL_PATH.io_enq_req_0_bits_instr; \
        force U_IF_NAME.io_enq_req_0_bits_pc = RTL_PATH.io_enq_req_0_bits_pc; \
        force U_IF_NAME.io_enq_req_0_bits_exceptionVec_0 = RTL_PATH.io_enq_req_0_bits_exceptionVec_0; \
        force U_IF_NAME.io_enq_req_0_bits_exceptionVec_1 = RTL_PATH.io_enq_req_0_bits_exceptionVec_1; \
        force U_IF_NAME.io_enq_req_0_bits_exceptionVec_2 = RTL_PATH.io_enq_req_0_bits_exceptionVec_2; \
        force U_IF_NAME.io_enq_req_0_bits_exceptionVec_3 = RTL_PATH.io_enq_req_0_bits_exceptionVec_3; \
        force U_IF_NAME.io_enq_req_0_bits_exceptionVec_12 = RTL_PATH.io_enq_req_0_bits_exceptionVec_12; \
        force U_IF_NAME.io_enq_req_0_bits_exceptionVec_20 = RTL_PATH.io_enq_req_0_bits_exceptionVec_20; \
        force U_IF_NAME.io_enq_req_0_bits_exceptionVec_22 = RTL_PATH.io_enq_req_0_bits_exceptionVec_22; \
        force U_IF_NAME.io_enq_req_0_bits_isFetchMalAddr = RTL_PATH.io_enq_req_0_bits_isFetchMalAddr; \
        force U_IF_NAME.io_enq_req_0_bits_hasException = RTL_PATH.io_enq_req_0_bits_hasException; \
        force U_IF_NAME.io_enq_req_0_bits_trigger = RTL_PATH.io_enq_req_0_bits_trigger; \
        force U_IF_NAME.io_enq_req_0_bits_preDecodeInfo_isRVC = RTL_PATH.io_enq_req_0_bits_preDecodeInfo_isRVC; \
        force U_IF_NAME.io_enq_req_0_bits_crossPageIPFFix = RTL_PATH.io_enq_req_0_bits_crossPageIPFFix; \
        force U_IF_NAME.io_enq_req_0_bits_ftqPtr_flag = RTL_PATH.io_enq_req_0_bits_ftqPtr_flag; \
        force U_IF_NAME.io_enq_req_0_bits_ftqPtr_value = RTL_PATH.io_enq_req_0_bits_ftqPtr_value; \
        force U_IF_NAME.io_enq_req_0_bits_ftqOffset = RTL_PATH.io_enq_req_0_bits_ftqOffset; \
        force U_IF_NAME.io_enq_req_0_bits_ldest = RTL_PATH.io_enq_req_0_bits_ldest; \
        force U_IF_NAME.io_enq_req_0_bits_fuType = RTL_PATH.io_enq_req_0_bits_fuType; \
        force U_IF_NAME.io_enq_req_0_bits_fuOpType = RTL_PATH.io_enq_req_0_bits_fuOpType; \
        force U_IF_NAME.io_enq_req_0_bits_rfWen = RTL_PATH.io_enq_req_0_bits_rfWen; \
        force U_IF_NAME.io_enq_req_0_bits_fpWen = RTL_PATH.io_enq_req_0_bits_fpWen; \
        force U_IF_NAME.io_enq_req_0_bits_vecWen = RTL_PATH.io_enq_req_0_bits_vecWen; \
        force U_IF_NAME.io_enq_req_0_bits_v0Wen = RTL_PATH.io_enq_req_0_bits_v0Wen; \
        force U_IF_NAME.io_enq_req_0_bits_vlWen = RTL_PATH.io_enq_req_0_bits_vlWen; \
        force U_IF_NAME.io_enq_req_0_bits_isXSTrap = RTL_PATH.io_enq_req_0_bits_isXSTrap; \
        force U_IF_NAME.io_enq_req_0_bits_waitForward = RTL_PATH.io_enq_req_0_bits_waitForward; \
        force U_IF_NAME.io_enq_req_0_bits_blockBackward = RTL_PATH.io_enq_req_0_bits_blockBackward; \
        force U_IF_NAME.io_enq_req_0_bits_flushPipe = RTL_PATH.io_enq_req_0_bits_flushPipe; \
        force U_IF_NAME.io_enq_req_0_bits_vpu_vill = RTL_PATH.io_enq_req_0_bits_vpu_vill; \
        force U_IF_NAME.io_enq_req_0_bits_vpu_vma = RTL_PATH.io_enq_req_0_bits_vpu_vma; \
        force U_IF_NAME.io_enq_req_0_bits_vpu_vta = RTL_PATH.io_enq_req_0_bits_vpu_vta; \
        force U_IF_NAME.io_enq_req_0_bits_vpu_vsew = RTL_PATH.io_enq_req_0_bits_vpu_vsew; \
        force U_IF_NAME.io_enq_req_0_bits_vpu_vlmul = RTL_PATH.io_enq_req_0_bits_vpu_vlmul; \
        force U_IF_NAME.io_enq_req_0_bits_vpu_specVill = RTL_PATH.io_enq_req_0_bits_vpu_specVill; \
        force U_IF_NAME.io_enq_req_0_bits_vpu_specVma = RTL_PATH.io_enq_req_0_bits_vpu_specVma; \
        force U_IF_NAME.io_enq_req_0_bits_vpu_specVta = RTL_PATH.io_enq_req_0_bits_vpu_specVta; \
        force U_IF_NAME.io_enq_req_0_bits_vpu_specVsew = RTL_PATH.io_enq_req_0_bits_vpu_specVsew; \
        force U_IF_NAME.io_enq_req_0_bits_vpu_specVlmul = RTL_PATH.io_enq_req_0_bits_vpu_specVlmul; \
        force U_IF_NAME.io_enq_req_0_bits_vlsInstr = RTL_PATH.io_enq_req_0_bits_vlsInstr; \
        force U_IF_NAME.io_enq_req_0_bits_wfflags = RTL_PATH.io_enq_req_0_bits_wfflags; \
        force U_IF_NAME.io_enq_req_0_bits_isMove = RTL_PATH.io_enq_req_0_bits_isMove; \
        force U_IF_NAME.io_enq_req_0_bits_isVset = RTL_PATH.io_enq_req_0_bits_isVset; \
        force U_IF_NAME.io_enq_req_0_bits_firstUop = RTL_PATH.io_enq_req_0_bits_firstUop; \
        force U_IF_NAME.io_enq_req_0_bits_lastUop = RTL_PATH.io_enq_req_0_bits_lastUop; \
        force U_IF_NAME.io_enq_req_0_bits_numWB = RTL_PATH.io_enq_req_0_bits_numWB; \
        force U_IF_NAME.io_enq_req_0_bits_commitType = RTL_PATH.io_enq_req_0_bits_commitType; \
        force U_IF_NAME.io_enq_req_0_bits_pdest = RTL_PATH.io_enq_req_0_bits_pdest; \
        force U_IF_NAME.io_enq_req_0_bits_robIdx_flag = RTL_PATH.io_enq_req_0_bits_robIdx_flag; \
        force U_IF_NAME.io_enq_req_0_bits_robIdx_value = RTL_PATH.io_enq_req_0_bits_robIdx_value; \
        force U_IF_NAME.io_enq_req_0_bits_instrSize = RTL_PATH.io_enq_req_0_bits_instrSize; \
        force U_IF_NAME.io_enq_req_0_bits_dirtyFs = RTL_PATH.io_enq_req_0_bits_dirtyFs; \
        force U_IF_NAME.io_enq_req_0_bits_dirtyVs = RTL_PATH.io_enq_req_0_bits_dirtyVs; \
        force U_IF_NAME.io_enq_req_0_bits_traceBlockInPipe_itype = RTL_PATH.io_enq_req_0_bits_traceBlockInPipe_itype; \
        force U_IF_NAME.io_enq_req_0_bits_traceBlockInPipe_iretire = RTL_PATH.io_enq_req_0_bits_traceBlockInPipe_iretire; \
        force U_IF_NAME.io_enq_req_0_bits_traceBlockInPipe_ilastsize = RTL_PATH.io_enq_req_0_bits_traceBlockInPipe_ilastsize; \
        force U_IF_NAME.io_enq_req_0_bits_eliminatedMove = RTL_PATH.io_enq_req_0_bits_eliminatedMove; \
        force U_IF_NAME.io_enq_req_0_bits_snapshot = RTL_PATH.io_enq_req_0_bits_snapshot; \
        force U_IF_NAME.io_enq_req_0_bits_lqIdx_value = RTL_PATH.io_enq_req_0_bits_lqIdx_value; \
        force U_IF_NAME.io_enq_req_0_bits_sqIdx_value = RTL_PATH.io_enq_req_0_bits_sqIdx_value; \
        force U_IF_NAME.io_enq_req_0_bits_singleStep = RTL_PATH.io_enq_req_0_bits_singleStep; \
        force U_IF_NAME.io_enq_req_0_bits_debug_sim_trig = RTL_PATH.io_enq_req_0_bits_debug_sim_trig; \
        force U_IF_NAME.io_enq_req_1_valid = RTL_PATH.io_enq_req_1_valid; \
        force U_IF_NAME.io_enq_req_1_bits_instr = RTL_PATH.io_enq_req_1_bits_instr; \
        force U_IF_NAME.io_enq_req_1_bits_pc = RTL_PATH.io_enq_req_1_bits_pc; \
        force U_IF_NAME.io_enq_req_1_bits_exceptionVec_0 = RTL_PATH.io_enq_req_1_bits_exceptionVec_0; \
        force U_IF_NAME.io_enq_req_1_bits_exceptionVec_1 = RTL_PATH.io_enq_req_1_bits_exceptionVec_1; \
        force U_IF_NAME.io_enq_req_1_bits_exceptionVec_2 = RTL_PATH.io_enq_req_1_bits_exceptionVec_2; \
        force U_IF_NAME.io_enq_req_1_bits_exceptionVec_3 = RTL_PATH.io_enq_req_1_bits_exceptionVec_3; \
        force U_IF_NAME.io_enq_req_1_bits_exceptionVec_12 = RTL_PATH.io_enq_req_1_bits_exceptionVec_12; \
        force U_IF_NAME.io_enq_req_1_bits_exceptionVec_20 = RTL_PATH.io_enq_req_1_bits_exceptionVec_20; \
        force U_IF_NAME.io_enq_req_1_bits_exceptionVec_22 = RTL_PATH.io_enq_req_1_bits_exceptionVec_22; \
        force U_IF_NAME.io_enq_req_1_bits_isFetchMalAddr = RTL_PATH.io_enq_req_1_bits_isFetchMalAddr; \
        force U_IF_NAME.io_enq_req_1_bits_hasException = RTL_PATH.io_enq_req_1_bits_hasException; \
        force U_IF_NAME.io_enq_req_1_bits_trigger = RTL_PATH.io_enq_req_1_bits_trigger; \
        force U_IF_NAME.io_enq_req_1_bits_preDecodeInfo_isRVC = RTL_PATH.io_enq_req_1_bits_preDecodeInfo_isRVC; \
        force U_IF_NAME.io_enq_req_1_bits_crossPageIPFFix = RTL_PATH.io_enq_req_1_bits_crossPageIPFFix; \
        force U_IF_NAME.io_enq_req_1_bits_ftqPtr_flag = RTL_PATH.io_enq_req_1_bits_ftqPtr_flag; \
        force U_IF_NAME.io_enq_req_1_bits_ftqPtr_value = RTL_PATH.io_enq_req_1_bits_ftqPtr_value; \
        force U_IF_NAME.io_enq_req_1_bits_ftqOffset = RTL_PATH.io_enq_req_1_bits_ftqOffset; \
        force U_IF_NAME.io_enq_req_1_bits_ldest = RTL_PATH.io_enq_req_1_bits_ldest; \
        force U_IF_NAME.io_enq_req_1_bits_fuType = RTL_PATH.io_enq_req_1_bits_fuType; \
        force U_IF_NAME.io_enq_req_1_bits_fuOpType = RTL_PATH.io_enq_req_1_bits_fuOpType; \
        force U_IF_NAME.io_enq_req_1_bits_rfWen = RTL_PATH.io_enq_req_1_bits_rfWen; \
        force U_IF_NAME.io_enq_req_1_bits_fpWen = RTL_PATH.io_enq_req_1_bits_fpWen; \
        force U_IF_NAME.io_enq_req_1_bits_vecWen = RTL_PATH.io_enq_req_1_bits_vecWen; \
        force U_IF_NAME.io_enq_req_1_bits_v0Wen = RTL_PATH.io_enq_req_1_bits_v0Wen; \
        force U_IF_NAME.io_enq_req_1_bits_vlWen = RTL_PATH.io_enq_req_1_bits_vlWen; \
        force U_IF_NAME.io_enq_req_1_bits_isXSTrap = RTL_PATH.io_enq_req_1_bits_isXSTrap; \
        force U_IF_NAME.io_enq_req_1_bits_waitForward = RTL_PATH.io_enq_req_1_bits_waitForward; \
        force U_IF_NAME.io_enq_req_1_bits_blockBackward = RTL_PATH.io_enq_req_1_bits_blockBackward; \
        force U_IF_NAME.io_enq_req_1_bits_flushPipe = RTL_PATH.io_enq_req_1_bits_flushPipe; \
        force U_IF_NAME.io_enq_req_1_bits_vpu_vill = RTL_PATH.io_enq_req_1_bits_vpu_vill; \
        force U_IF_NAME.io_enq_req_1_bits_vpu_vma = RTL_PATH.io_enq_req_1_bits_vpu_vma; \
        force U_IF_NAME.io_enq_req_1_bits_vpu_vta = RTL_PATH.io_enq_req_1_bits_vpu_vta; \
        force U_IF_NAME.io_enq_req_1_bits_vpu_vsew = RTL_PATH.io_enq_req_1_bits_vpu_vsew; \
        force U_IF_NAME.io_enq_req_1_bits_vpu_vlmul = RTL_PATH.io_enq_req_1_bits_vpu_vlmul; \
        force U_IF_NAME.io_enq_req_1_bits_vpu_specVill = RTL_PATH.io_enq_req_1_bits_vpu_specVill; \
        force U_IF_NAME.io_enq_req_1_bits_vpu_specVma = RTL_PATH.io_enq_req_1_bits_vpu_specVma; \
        force U_IF_NAME.io_enq_req_1_bits_vpu_specVta = RTL_PATH.io_enq_req_1_bits_vpu_specVta; \
        force U_IF_NAME.io_enq_req_1_bits_vpu_specVsew = RTL_PATH.io_enq_req_1_bits_vpu_specVsew; \
        force U_IF_NAME.io_enq_req_1_bits_vpu_specVlmul = RTL_PATH.io_enq_req_1_bits_vpu_specVlmul; \
        force U_IF_NAME.io_enq_req_1_bits_vlsInstr = RTL_PATH.io_enq_req_1_bits_vlsInstr; \
        force U_IF_NAME.io_enq_req_1_bits_wfflags = RTL_PATH.io_enq_req_1_bits_wfflags; \
        force U_IF_NAME.io_enq_req_1_bits_isMove = RTL_PATH.io_enq_req_1_bits_isMove; \
        force U_IF_NAME.io_enq_req_1_bits_isVset = RTL_PATH.io_enq_req_1_bits_isVset; \
        force U_IF_NAME.io_enq_req_1_bits_firstUop = RTL_PATH.io_enq_req_1_bits_firstUop; \
        force U_IF_NAME.io_enq_req_1_bits_lastUop = RTL_PATH.io_enq_req_1_bits_lastUop; \
        force U_IF_NAME.io_enq_req_1_bits_numWB = RTL_PATH.io_enq_req_1_bits_numWB; \
        force U_IF_NAME.io_enq_req_1_bits_commitType = RTL_PATH.io_enq_req_1_bits_commitType; \
        force U_IF_NAME.io_enq_req_1_bits_pdest = RTL_PATH.io_enq_req_1_bits_pdest; \
        force U_IF_NAME.io_enq_req_1_bits_robIdx_flag = RTL_PATH.io_enq_req_1_bits_robIdx_flag; \
        force U_IF_NAME.io_enq_req_1_bits_robIdx_value = RTL_PATH.io_enq_req_1_bits_robIdx_value; \
        force U_IF_NAME.io_enq_req_1_bits_instrSize = RTL_PATH.io_enq_req_1_bits_instrSize; \
        force U_IF_NAME.io_enq_req_1_bits_dirtyFs = RTL_PATH.io_enq_req_1_bits_dirtyFs; \
        force U_IF_NAME.io_enq_req_1_bits_dirtyVs = RTL_PATH.io_enq_req_1_bits_dirtyVs; \
        force U_IF_NAME.io_enq_req_1_bits_traceBlockInPipe_itype = RTL_PATH.io_enq_req_1_bits_traceBlockInPipe_itype; \
        force U_IF_NAME.io_enq_req_1_bits_traceBlockInPipe_iretire = RTL_PATH.io_enq_req_1_bits_traceBlockInPipe_iretire; \
        force U_IF_NAME.io_enq_req_1_bits_traceBlockInPipe_ilastsize = RTL_PATH.io_enq_req_1_bits_traceBlockInPipe_ilastsize; \
        force U_IF_NAME.io_enq_req_1_bits_eliminatedMove = RTL_PATH.io_enq_req_1_bits_eliminatedMove; \
        force U_IF_NAME.io_enq_req_1_bits_snapshot = RTL_PATH.io_enq_req_1_bits_snapshot; \
        force U_IF_NAME.io_enq_req_1_bits_lqIdx_value = RTL_PATH.io_enq_req_1_bits_lqIdx_value; \
        force U_IF_NAME.io_enq_req_1_bits_sqIdx_value = RTL_PATH.io_enq_req_1_bits_sqIdx_value; \
        force U_IF_NAME.io_enq_req_1_bits_singleStep = RTL_PATH.io_enq_req_1_bits_singleStep; \
        force U_IF_NAME.io_enq_req_1_bits_debug_sim_trig = RTL_PATH.io_enq_req_1_bits_debug_sim_trig; \
        force U_IF_NAME.io_enq_req_2_valid = RTL_PATH.io_enq_req_2_valid; \
        force U_IF_NAME.io_enq_req_2_bits_instr = RTL_PATH.io_enq_req_2_bits_instr; \
        force U_IF_NAME.io_enq_req_2_bits_pc = RTL_PATH.io_enq_req_2_bits_pc; \
        force U_IF_NAME.io_enq_req_2_bits_exceptionVec_0 = RTL_PATH.io_enq_req_2_bits_exceptionVec_0; \
        force U_IF_NAME.io_enq_req_2_bits_exceptionVec_1 = RTL_PATH.io_enq_req_2_bits_exceptionVec_1; \
        force U_IF_NAME.io_enq_req_2_bits_exceptionVec_2 = RTL_PATH.io_enq_req_2_bits_exceptionVec_2; \
        force U_IF_NAME.io_enq_req_2_bits_exceptionVec_3 = RTL_PATH.io_enq_req_2_bits_exceptionVec_3; \
        force U_IF_NAME.io_enq_req_2_bits_exceptionVec_12 = RTL_PATH.io_enq_req_2_bits_exceptionVec_12; \
        force U_IF_NAME.io_enq_req_2_bits_exceptionVec_20 = RTL_PATH.io_enq_req_2_bits_exceptionVec_20; \
        force U_IF_NAME.io_enq_req_2_bits_exceptionVec_22 = RTL_PATH.io_enq_req_2_bits_exceptionVec_22; \
        force U_IF_NAME.io_enq_req_2_bits_isFetchMalAddr = RTL_PATH.io_enq_req_2_bits_isFetchMalAddr; \
        force U_IF_NAME.io_enq_req_2_bits_hasException = RTL_PATH.io_enq_req_2_bits_hasException; \
        force U_IF_NAME.io_enq_req_2_bits_trigger = RTL_PATH.io_enq_req_2_bits_trigger; \
        force U_IF_NAME.io_enq_req_2_bits_preDecodeInfo_isRVC = RTL_PATH.io_enq_req_2_bits_preDecodeInfo_isRVC; \
        force U_IF_NAME.io_enq_req_2_bits_crossPageIPFFix = RTL_PATH.io_enq_req_2_bits_crossPageIPFFix; \
        force U_IF_NAME.io_enq_req_2_bits_ftqPtr_flag = RTL_PATH.io_enq_req_2_bits_ftqPtr_flag; \
        force U_IF_NAME.io_enq_req_2_bits_ftqPtr_value = RTL_PATH.io_enq_req_2_bits_ftqPtr_value; \
        force U_IF_NAME.io_enq_req_2_bits_ftqOffset = RTL_PATH.io_enq_req_2_bits_ftqOffset; \
        force U_IF_NAME.io_enq_req_2_bits_ldest = RTL_PATH.io_enq_req_2_bits_ldest; \
        force U_IF_NAME.io_enq_req_2_bits_fuType = RTL_PATH.io_enq_req_2_bits_fuType; \
        force U_IF_NAME.io_enq_req_2_bits_fuOpType = RTL_PATH.io_enq_req_2_bits_fuOpType; \
        force U_IF_NAME.io_enq_req_2_bits_rfWen = RTL_PATH.io_enq_req_2_bits_rfWen; \
        force U_IF_NAME.io_enq_req_2_bits_fpWen = RTL_PATH.io_enq_req_2_bits_fpWen; \
        force U_IF_NAME.io_enq_req_2_bits_vecWen = RTL_PATH.io_enq_req_2_bits_vecWen; \
        force U_IF_NAME.io_enq_req_2_bits_v0Wen = RTL_PATH.io_enq_req_2_bits_v0Wen; \
        force U_IF_NAME.io_enq_req_2_bits_vlWen = RTL_PATH.io_enq_req_2_bits_vlWen; \
        force U_IF_NAME.io_enq_req_2_bits_isXSTrap = RTL_PATH.io_enq_req_2_bits_isXSTrap; \
        force U_IF_NAME.io_enq_req_2_bits_waitForward = RTL_PATH.io_enq_req_2_bits_waitForward; \
        force U_IF_NAME.io_enq_req_2_bits_blockBackward = RTL_PATH.io_enq_req_2_bits_blockBackward; \
        force U_IF_NAME.io_enq_req_2_bits_flushPipe = RTL_PATH.io_enq_req_2_bits_flushPipe; \
        force U_IF_NAME.io_enq_req_2_bits_vpu_vill = RTL_PATH.io_enq_req_2_bits_vpu_vill; \
        force U_IF_NAME.io_enq_req_2_bits_vpu_vma = RTL_PATH.io_enq_req_2_bits_vpu_vma; \
        force U_IF_NAME.io_enq_req_2_bits_vpu_vta = RTL_PATH.io_enq_req_2_bits_vpu_vta; \
        force U_IF_NAME.io_enq_req_2_bits_vpu_vsew = RTL_PATH.io_enq_req_2_bits_vpu_vsew; \
        force U_IF_NAME.io_enq_req_2_bits_vpu_vlmul = RTL_PATH.io_enq_req_2_bits_vpu_vlmul; \
        force U_IF_NAME.io_enq_req_2_bits_vpu_specVill = RTL_PATH.io_enq_req_2_bits_vpu_specVill; \
        force U_IF_NAME.io_enq_req_2_bits_vpu_specVma = RTL_PATH.io_enq_req_2_bits_vpu_specVma; \
        force U_IF_NAME.io_enq_req_2_bits_vpu_specVta = RTL_PATH.io_enq_req_2_bits_vpu_specVta; \
        force U_IF_NAME.io_enq_req_2_bits_vpu_specVsew = RTL_PATH.io_enq_req_2_bits_vpu_specVsew; \
        force U_IF_NAME.io_enq_req_2_bits_vpu_specVlmul = RTL_PATH.io_enq_req_2_bits_vpu_specVlmul; \
        force U_IF_NAME.io_enq_req_2_bits_vlsInstr = RTL_PATH.io_enq_req_2_bits_vlsInstr; \
        force U_IF_NAME.io_enq_req_2_bits_wfflags = RTL_PATH.io_enq_req_2_bits_wfflags; \
        force U_IF_NAME.io_enq_req_2_bits_isMove = RTL_PATH.io_enq_req_2_bits_isMove; \
        force U_IF_NAME.io_enq_req_2_bits_isVset = RTL_PATH.io_enq_req_2_bits_isVset; \
        force U_IF_NAME.io_enq_req_2_bits_firstUop = RTL_PATH.io_enq_req_2_bits_firstUop; \
        force U_IF_NAME.io_enq_req_2_bits_lastUop = RTL_PATH.io_enq_req_2_bits_lastUop; \
        force U_IF_NAME.io_enq_req_2_bits_numWB = RTL_PATH.io_enq_req_2_bits_numWB; \
        force U_IF_NAME.io_enq_req_2_bits_commitType = RTL_PATH.io_enq_req_2_bits_commitType; \
        force U_IF_NAME.io_enq_req_2_bits_pdest = RTL_PATH.io_enq_req_2_bits_pdest; \
        force U_IF_NAME.io_enq_req_2_bits_robIdx_flag = RTL_PATH.io_enq_req_2_bits_robIdx_flag; \
        force U_IF_NAME.io_enq_req_2_bits_robIdx_value = RTL_PATH.io_enq_req_2_bits_robIdx_value; \
        force U_IF_NAME.io_enq_req_2_bits_instrSize = RTL_PATH.io_enq_req_2_bits_instrSize; \
        force U_IF_NAME.io_enq_req_2_bits_dirtyFs = RTL_PATH.io_enq_req_2_bits_dirtyFs; \
        force U_IF_NAME.io_enq_req_2_bits_dirtyVs = RTL_PATH.io_enq_req_2_bits_dirtyVs; \
        force U_IF_NAME.io_enq_req_2_bits_traceBlockInPipe_itype = RTL_PATH.io_enq_req_2_bits_traceBlockInPipe_itype; \
        force U_IF_NAME.io_enq_req_2_bits_traceBlockInPipe_iretire = RTL_PATH.io_enq_req_2_bits_traceBlockInPipe_iretire; \
        force U_IF_NAME.io_enq_req_2_bits_traceBlockInPipe_ilastsize = RTL_PATH.io_enq_req_2_bits_traceBlockInPipe_ilastsize; \
        force U_IF_NAME.io_enq_req_2_bits_eliminatedMove = RTL_PATH.io_enq_req_2_bits_eliminatedMove; \
        force U_IF_NAME.io_enq_req_2_bits_snapshot = RTL_PATH.io_enq_req_2_bits_snapshot; \
        force U_IF_NAME.io_enq_req_2_bits_lqIdx_value = RTL_PATH.io_enq_req_2_bits_lqIdx_value; \
        force U_IF_NAME.io_enq_req_2_bits_sqIdx_value = RTL_PATH.io_enq_req_2_bits_sqIdx_value; \
        force U_IF_NAME.io_enq_req_2_bits_singleStep = RTL_PATH.io_enq_req_2_bits_singleStep; \
        force U_IF_NAME.io_enq_req_2_bits_debug_sim_trig = RTL_PATH.io_enq_req_2_bits_debug_sim_trig; \
        force U_IF_NAME.io_enq_req_3_valid = RTL_PATH.io_enq_req_3_valid; \
        force U_IF_NAME.io_enq_req_3_bits_instr = RTL_PATH.io_enq_req_3_bits_instr; \
        force U_IF_NAME.io_enq_req_3_bits_pc = RTL_PATH.io_enq_req_3_bits_pc; \
        force U_IF_NAME.io_enq_req_3_bits_exceptionVec_0 = RTL_PATH.io_enq_req_3_bits_exceptionVec_0; \
        force U_IF_NAME.io_enq_req_3_bits_exceptionVec_1 = RTL_PATH.io_enq_req_3_bits_exceptionVec_1; \
        force U_IF_NAME.io_enq_req_3_bits_exceptionVec_2 = RTL_PATH.io_enq_req_3_bits_exceptionVec_2; \
        force U_IF_NAME.io_enq_req_3_bits_exceptionVec_3 = RTL_PATH.io_enq_req_3_bits_exceptionVec_3; \
        force U_IF_NAME.io_enq_req_3_bits_exceptionVec_12 = RTL_PATH.io_enq_req_3_bits_exceptionVec_12; \
        force U_IF_NAME.io_enq_req_3_bits_exceptionVec_20 = RTL_PATH.io_enq_req_3_bits_exceptionVec_20; \
        force U_IF_NAME.io_enq_req_3_bits_exceptionVec_22 = RTL_PATH.io_enq_req_3_bits_exceptionVec_22; \
        force U_IF_NAME.io_enq_req_3_bits_isFetchMalAddr = RTL_PATH.io_enq_req_3_bits_isFetchMalAddr; \
        force U_IF_NAME.io_enq_req_3_bits_hasException = RTL_PATH.io_enq_req_3_bits_hasException; \
        force U_IF_NAME.io_enq_req_3_bits_trigger = RTL_PATH.io_enq_req_3_bits_trigger; \
        force U_IF_NAME.io_enq_req_3_bits_preDecodeInfo_isRVC = RTL_PATH.io_enq_req_3_bits_preDecodeInfo_isRVC; \
        force U_IF_NAME.io_enq_req_3_bits_crossPageIPFFix = RTL_PATH.io_enq_req_3_bits_crossPageIPFFix; \
        force U_IF_NAME.io_enq_req_3_bits_ftqPtr_flag = RTL_PATH.io_enq_req_3_bits_ftqPtr_flag; \
        force U_IF_NAME.io_enq_req_3_bits_ftqPtr_value = RTL_PATH.io_enq_req_3_bits_ftqPtr_value; \
        force U_IF_NAME.io_enq_req_3_bits_ftqOffset = RTL_PATH.io_enq_req_3_bits_ftqOffset; \
        force U_IF_NAME.io_enq_req_3_bits_ldest = RTL_PATH.io_enq_req_3_bits_ldest; \
        force U_IF_NAME.io_enq_req_3_bits_fuType = RTL_PATH.io_enq_req_3_bits_fuType; \
        force U_IF_NAME.io_enq_req_3_bits_fuOpType = RTL_PATH.io_enq_req_3_bits_fuOpType; \
        force U_IF_NAME.io_enq_req_3_bits_rfWen = RTL_PATH.io_enq_req_3_bits_rfWen; \
        force U_IF_NAME.io_enq_req_3_bits_fpWen = RTL_PATH.io_enq_req_3_bits_fpWen; \
        force U_IF_NAME.io_enq_req_3_bits_vecWen = RTL_PATH.io_enq_req_3_bits_vecWen; \
        force U_IF_NAME.io_enq_req_3_bits_v0Wen = RTL_PATH.io_enq_req_3_bits_v0Wen; \
        force U_IF_NAME.io_enq_req_3_bits_vlWen = RTL_PATH.io_enq_req_3_bits_vlWen; \
        force U_IF_NAME.io_enq_req_3_bits_isXSTrap = RTL_PATH.io_enq_req_3_bits_isXSTrap; \
        force U_IF_NAME.io_enq_req_3_bits_waitForward = RTL_PATH.io_enq_req_3_bits_waitForward; \
        force U_IF_NAME.io_enq_req_3_bits_blockBackward = RTL_PATH.io_enq_req_3_bits_blockBackward; \
        force U_IF_NAME.io_enq_req_3_bits_flushPipe = RTL_PATH.io_enq_req_3_bits_flushPipe; \
        force U_IF_NAME.io_enq_req_3_bits_vpu_vill = RTL_PATH.io_enq_req_3_bits_vpu_vill; \
        force U_IF_NAME.io_enq_req_3_bits_vpu_vma = RTL_PATH.io_enq_req_3_bits_vpu_vma; \
        force U_IF_NAME.io_enq_req_3_bits_vpu_vta = RTL_PATH.io_enq_req_3_bits_vpu_vta; \
        force U_IF_NAME.io_enq_req_3_bits_vpu_vsew = RTL_PATH.io_enq_req_3_bits_vpu_vsew; \
        force U_IF_NAME.io_enq_req_3_bits_vpu_vlmul = RTL_PATH.io_enq_req_3_bits_vpu_vlmul; \
        force U_IF_NAME.io_enq_req_3_bits_vpu_specVill = RTL_PATH.io_enq_req_3_bits_vpu_specVill; \
        force U_IF_NAME.io_enq_req_3_bits_vpu_specVma = RTL_PATH.io_enq_req_3_bits_vpu_specVma; \
        force U_IF_NAME.io_enq_req_3_bits_vpu_specVta = RTL_PATH.io_enq_req_3_bits_vpu_specVta; \
        force U_IF_NAME.io_enq_req_3_bits_vpu_specVsew = RTL_PATH.io_enq_req_3_bits_vpu_specVsew; \
        force U_IF_NAME.io_enq_req_3_bits_vpu_specVlmul = RTL_PATH.io_enq_req_3_bits_vpu_specVlmul; \
        force U_IF_NAME.io_enq_req_3_bits_vlsInstr = RTL_PATH.io_enq_req_3_bits_vlsInstr; \
        force U_IF_NAME.io_enq_req_3_bits_wfflags = RTL_PATH.io_enq_req_3_bits_wfflags; \
        force U_IF_NAME.io_enq_req_3_bits_isMove = RTL_PATH.io_enq_req_3_bits_isMove; \
        force U_IF_NAME.io_enq_req_3_bits_isVset = RTL_PATH.io_enq_req_3_bits_isVset; \
        force U_IF_NAME.io_enq_req_3_bits_firstUop = RTL_PATH.io_enq_req_3_bits_firstUop; \
        force U_IF_NAME.io_enq_req_3_bits_lastUop = RTL_PATH.io_enq_req_3_bits_lastUop; \
        force U_IF_NAME.io_enq_req_3_bits_numWB = RTL_PATH.io_enq_req_3_bits_numWB; \
        force U_IF_NAME.io_enq_req_3_bits_commitType = RTL_PATH.io_enq_req_3_bits_commitType; \
        force U_IF_NAME.io_enq_req_3_bits_pdest = RTL_PATH.io_enq_req_3_bits_pdest; \
        force U_IF_NAME.io_enq_req_3_bits_robIdx_flag = RTL_PATH.io_enq_req_3_bits_robIdx_flag; \
        force U_IF_NAME.io_enq_req_3_bits_robIdx_value = RTL_PATH.io_enq_req_3_bits_robIdx_value; \
        force U_IF_NAME.io_enq_req_3_bits_instrSize = RTL_PATH.io_enq_req_3_bits_instrSize; \
        force U_IF_NAME.io_enq_req_3_bits_dirtyFs = RTL_PATH.io_enq_req_3_bits_dirtyFs; \
        force U_IF_NAME.io_enq_req_3_bits_dirtyVs = RTL_PATH.io_enq_req_3_bits_dirtyVs; \
        force U_IF_NAME.io_enq_req_3_bits_traceBlockInPipe_itype = RTL_PATH.io_enq_req_3_bits_traceBlockInPipe_itype; \
        force U_IF_NAME.io_enq_req_3_bits_traceBlockInPipe_iretire = RTL_PATH.io_enq_req_3_bits_traceBlockInPipe_iretire; \
        force U_IF_NAME.io_enq_req_3_bits_traceBlockInPipe_ilastsize = RTL_PATH.io_enq_req_3_bits_traceBlockInPipe_ilastsize; \
        force U_IF_NAME.io_enq_req_3_bits_eliminatedMove = RTL_PATH.io_enq_req_3_bits_eliminatedMove; \
        force U_IF_NAME.io_enq_req_3_bits_snapshot = RTL_PATH.io_enq_req_3_bits_snapshot; \
        force U_IF_NAME.io_enq_req_3_bits_lqIdx_value = RTL_PATH.io_enq_req_3_bits_lqIdx_value; \
        force U_IF_NAME.io_enq_req_3_bits_sqIdx_value = RTL_PATH.io_enq_req_3_bits_sqIdx_value; \
        force U_IF_NAME.io_enq_req_3_bits_singleStep = RTL_PATH.io_enq_req_3_bits_singleStep; \
        force U_IF_NAME.io_enq_req_3_bits_debug_sim_trig = RTL_PATH.io_enq_req_3_bits_debug_sim_trig; \
        force U_IF_NAME.io_enq_req_4_valid = RTL_PATH.io_enq_req_4_valid; \
        force U_IF_NAME.io_enq_req_4_bits_instr = RTL_PATH.io_enq_req_4_bits_instr; \
        force U_IF_NAME.io_enq_req_4_bits_pc = RTL_PATH.io_enq_req_4_bits_pc; \
        force U_IF_NAME.io_enq_req_4_bits_exceptionVec_0 = RTL_PATH.io_enq_req_4_bits_exceptionVec_0; \
        force U_IF_NAME.io_enq_req_4_bits_exceptionVec_1 = RTL_PATH.io_enq_req_4_bits_exceptionVec_1; \
        force U_IF_NAME.io_enq_req_4_bits_exceptionVec_2 = RTL_PATH.io_enq_req_4_bits_exceptionVec_2; \
        force U_IF_NAME.io_enq_req_4_bits_exceptionVec_3 = RTL_PATH.io_enq_req_4_bits_exceptionVec_3; \
        force U_IF_NAME.io_enq_req_4_bits_exceptionVec_12 = RTL_PATH.io_enq_req_4_bits_exceptionVec_12; \
        force U_IF_NAME.io_enq_req_4_bits_exceptionVec_20 = RTL_PATH.io_enq_req_4_bits_exceptionVec_20; \
        force U_IF_NAME.io_enq_req_4_bits_exceptionVec_22 = RTL_PATH.io_enq_req_4_bits_exceptionVec_22; \
        force U_IF_NAME.io_enq_req_4_bits_isFetchMalAddr = RTL_PATH.io_enq_req_4_bits_isFetchMalAddr; \
        force U_IF_NAME.io_enq_req_4_bits_hasException = RTL_PATH.io_enq_req_4_bits_hasException; \
        force U_IF_NAME.io_enq_req_4_bits_trigger = RTL_PATH.io_enq_req_4_bits_trigger; \
        force U_IF_NAME.io_enq_req_4_bits_preDecodeInfo_isRVC = RTL_PATH.io_enq_req_4_bits_preDecodeInfo_isRVC; \
        force U_IF_NAME.io_enq_req_4_bits_crossPageIPFFix = RTL_PATH.io_enq_req_4_bits_crossPageIPFFix; \
        force U_IF_NAME.io_enq_req_4_bits_ftqPtr_flag = RTL_PATH.io_enq_req_4_bits_ftqPtr_flag; \
        force U_IF_NAME.io_enq_req_4_bits_ftqPtr_value = RTL_PATH.io_enq_req_4_bits_ftqPtr_value; \
        force U_IF_NAME.io_enq_req_4_bits_ftqOffset = RTL_PATH.io_enq_req_4_bits_ftqOffset; \
        force U_IF_NAME.io_enq_req_4_bits_ldest = RTL_PATH.io_enq_req_4_bits_ldest; \
        force U_IF_NAME.io_enq_req_4_bits_fuType = RTL_PATH.io_enq_req_4_bits_fuType; \
        force U_IF_NAME.io_enq_req_4_bits_fuOpType = RTL_PATH.io_enq_req_4_bits_fuOpType; \
        force U_IF_NAME.io_enq_req_4_bits_rfWen = RTL_PATH.io_enq_req_4_bits_rfWen; \
        force U_IF_NAME.io_enq_req_4_bits_fpWen = RTL_PATH.io_enq_req_4_bits_fpWen; \
        force U_IF_NAME.io_enq_req_4_bits_vecWen = RTL_PATH.io_enq_req_4_bits_vecWen; \
        force U_IF_NAME.io_enq_req_4_bits_v0Wen = RTL_PATH.io_enq_req_4_bits_v0Wen; \
        force U_IF_NAME.io_enq_req_4_bits_vlWen = RTL_PATH.io_enq_req_4_bits_vlWen; \
        force U_IF_NAME.io_enq_req_4_bits_isXSTrap = RTL_PATH.io_enq_req_4_bits_isXSTrap; \
        force U_IF_NAME.io_enq_req_4_bits_waitForward = RTL_PATH.io_enq_req_4_bits_waitForward; \
        force U_IF_NAME.io_enq_req_4_bits_blockBackward = RTL_PATH.io_enq_req_4_bits_blockBackward; \
        force U_IF_NAME.io_enq_req_4_bits_flushPipe = RTL_PATH.io_enq_req_4_bits_flushPipe; \
        force U_IF_NAME.io_enq_req_4_bits_vpu_vill = RTL_PATH.io_enq_req_4_bits_vpu_vill; \
        force U_IF_NAME.io_enq_req_4_bits_vpu_vma = RTL_PATH.io_enq_req_4_bits_vpu_vma; \
        force U_IF_NAME.io_enq_req_4_bits_vpu_vta = RTL_PATH.io_enq_req_4_bits_vpu_vta; \
        force U_IF_NAME.io_enq_req_4_bits_vpu_vsew = RTL_PATH.io_enq_req_4_bits_vpu_vsew; \
        force U_IF_NAME.io_enq_req_4_bits_vpu_vlmul = RTL_PATH.io_enq_req_4_bits_vpu_vlmul; \
        force U_IF_NAME.io_enq_req_4_bits_vpu_specVill = RTL_PATH.io_enq_req_4_bits_vpu_specVill; \
        force U_IF_NAME.io_enq_req_4_bits_vpu_specVma = RTL_PATH.io_enq_req_4_bits_vpu_specVma; \
        force U_IF_NAME.io_enq_req_4_bits_vpu_specVta = RTL_PATH.io_enq_req_4_bits_vpu_specVta; \
        force U_IF_NAME.io_enq_req_4_bits_vpu_specVsew = RTL_PATH.io_enq_req_4_bits_vpu_specVsew; \
        force U_IF_NAME.io_enq_req_4_bits_vpu_specVlmul = RTL_PATH.io_enq_req_4_bits_vpu_specVlmul; \
        force U_IF_NAME.io_enq_req_4_bits_vlsInstr = RTL_PATH.io_enq_req_4_bits_vlsInstr; \
        force U_IF_NAME.io_enq_req_4_bits_wfflags = RTL_PATH.io_enq_req_4_bits_wfflags; \
        force U_IF_NAME.io_enq_req_4_bits_isMove = RTL_PATH.io_enq_req_4_bits_isMove; \
        force U_IF_NAME.io_enq_req_4_bits_isVset = RTL_PATH.io_enq_req_4_bits_isVset; \
        force U_IF_NAME.io_enq_req_4_bits_firstUop = RTL_PATH.io_enq_req_4_bits_firstUop; \
        force U_IF_NAME.io_enq_req_4_bits_lastUop = RTL_PATH.io_enq_req_4_bits_lastUop; \
        force U_IF_NAME.io_enq_req_4_bits_numWB = RTL_PATH.io_enq_req_4_bits_numWB; \
        force U_IF_NAME.io_enq_req_4_bits_commitType = RTL_PATH.io_enq_req_4_bits_commitType; \
        force U_IF_NAME.io_enq_req_4_bits_pdest = RTL_PATH.io_enq_req_4_bits_pdest; \
        force U_IF_NAME.io_enq_req_4_bits_robIdx_flag = RTL_PATH.io_enq_req_4_bits_robIdx_flag; \
        force U_IF_NAME.io_enq_req_4_bits_robIdx_value = RTL_PATH.io_enq_req_4_bits_robIdx_value; \
        force U_IF_NAME.io_enq_req_4_bits_instrSize = RTL_PATH.io_enq_req_4_bits_instrSize; \
        force U_IF_NAME.io_enq_req_4_bits_dirtyFs = RTL_PATH.io_enq_req_4_bits_dirtyFs; \
        force U_IF_NAME.io_enq_req_4_bits_dirtyVs = RTL_PATH.io_enq_req_4_bits_dirtyVs; \
        force U_IF_NAME.io_enq_req_4_bits_traceBlockInPipe_itype = RTL_PATH.io_enq_req_4_bits_traceBlockInPipe_itype; \
        force U_IF_NAME.io_enq_req_4_bits_traceBlockInPipe_iretire = RTL_PATH.io_enq_req_4_bits_traceBlockInPipe_iretire; \
        force U_IF_NAME.io_enq_req_4_bits_traceBlockInPipe_ilastsize = RTL_PATH.io_enq_req_4_bits_traceBlockInPipe_ilastsize; \
        force U_IF_NAME.io_enq_req_4_bits_eliminatedMove = RTL_PATH.io_enq_req_4_bits_eliminatedMove; \
        force U_IF_NAME.io_enq_req_4_bits_snapshot = RTL_PATH.io_enq_req_4_bits_snapshot; \
        force U_IF_NAME.io_enq_req_4_bits_lqIdx_value = RTL_PATH.io_enq_req_4_bits_lqIdx_value; \
        force U_IF_NAME.io_enq_req_4_bits_sqIdx_value = RTL_PATH.io_enq_req_4_bits_sqIdx_value; \
        force U_IF_NAME.io_enq_req_4_bits_singleStep = RTL_PATH.io_enq_req_4_bits_singleStep; \
        force U_IF_NAME.io_enq_req_4_bits_debug_sim_trig = RTL_PATH.io_enq_req_4_bits_debug_sim_trig; \
        force U_IF_NAME.io_enq_req_5_valid = RTL_PATH.io_enq_req_5_valid; \
        force U_IF_NAME.io_enq_req_5_bits_instr = RTL_PATH.io_enq_req_5_bits_instr; \
        force U_IF_NAME.io_enq_req_5_bits_pc = RTL_PATH.io_enq_req_5_bits_pc; \
        force U_IF_NAME.io_enq_req_5_bits_exceptionVec_0 = RTL_PATH.io_enq_req_5_bits_exceptionVec_0; \
        force U_IF_NAME.io_enq_req_5_bits_exceptionVec_1 = RTL_PATH.io_enq_req_5_bits_exceptionVec_1; \
        force U_IF_NAME.io_enq_req_5_bits_exceptionVec_2 = RTL_PATH.io_enq_req_5_bits_exceptionVec_2; \
        force U_IF_NAME.io_enq_req_5_bits_exceptionVec_3 = RTL_PATH.io_enq_req_5_bits_exceptionVec_3; \
        force U_IF_NAME.io_enq_req_5_bits_exceptionVec_12 = RTL_PATH.io_enq_req_5_bits_exceptionVec_12; \
        force U_IF_NAME.io_enq_req_5_bits_exceptionVec_20 = RTL_PATH.io_enq_req_5_bits_exceptionVec_20; \
        force U_IF_NAME.io_enq_req_5_bits_exceptionVec_22 = RTL_PATH.io_enq_req_5_bits_exceptionVec_22; \
        force U_IF_NAME.io_enq_req_5_bits_isFetchMalAddr = RTL_PATH.io_enq_req_5_bits_isFetchMalAddr; \
        force U_IF_NAME.io_enq_req_5_bits_hasException = RTL_PATH.io_enq_req_5_bits_hasException; \
        force U_IF_NAME.io_enq_req_5_bits_trigger = RTL_PATH.io_enq_req_5_bits_trigger; \
        force U_IF_NAME.io_enq_req_5_bits_preDecodeInfo_isRVC = RTL_PATH.io_enq_req_5_bits_preDecodeInfo_isRVC; \
        force U_IF_NAME.io_enq_req_5_bits_crossPageIPFFix = RTL_PATH.io_enq_req_5_bits_crossPageIPFFix; \
        force U_IF_NAME.io_enq_req_5_bits_ftqPtr_flag = RTL_PATH.io_enq_req_5_bits_ftqPtr_flag; \
        force U_IF_NAME.io_enq_req_5_bits_ftqPtr_value = RTL_PATH.io_enq_req_5_bits_ftqPtr_value; \
        force U_IF_NAME.io_enq_req_5_bits_ftqOffset = RTL_PATH.io_enq_req_5_bits_ftqOffset; \
        force U_IF_NAME.io_enq_req_5_bits_ldest = RTL_PATH.io_enq_req_5_bits_ldest; \
        force U_IF_NAME.io_enq_req_5_bits_fuType = RTL_PATH.io_enq_req_5_bits_fuType; \
        force U_IF_NAME.io_enq_req_5_bits_fuOpType = RTL_PATH.io_enq_req_5_bits_fuOpType; \
        force U_IF_NAME.io_enq_req_5_bits_rfWen = RTL_PATH.io_enq_req_5_bits_rfWen; \
        force U_IF_NAME.io_enq_req_5_bits_fpWen = RTL_PATH.io_enq_req_5_bits_fpWen; \
        force U_IF_NAME.io_enq_req_5_bits_vecWen = RTL_PATH.io_enq_req_5_bits_vecWen; \
        force U_IF_NAME.io_enq_req_5_bits_v0Wen = RTL_PATH.io_enq_req_5_bits_v0Wen; \
        force U_IF_NAME.io_enq_req_5_bits_vlWen = RTL_PATH.io_enq_req_5_bits_vlWen; \
        force U_IF_NAME.io_enq_req_5_bits_isXSTrap = RTL_PATH.io_enq_req_5_bits_isXSTrap; \
        force U_IF_NAME.io_enq_req_5_bits_waitForward = RTL_PATH.io_enq_req_5_bits_waitForward; \
        force U_IF_NAME.io_enq_req_5_bits_blockBackward = RTL_PATH.io_enq_req_5_bits_blockBackward; \
        force U_IF_NAME.io_enq_req_5_bits_flushPipe = RTL_PATH.io_enq_req_5_bits_flushPipe; \
        force U_IF_NAME.io_enq_req_5_bits_vpu_vill = RTL_PATH.io_enq_req_5_bits_vpu_vill; \
        force U_IF_NAME.io_enq_req_5_bits_vpu_vma = RTL_PATH.io_enq_req_5_bits_vpu_vma; \
        force U_IF_NAME.io_enq_req_5_bits_vpu_vta = RTL_PATH.io_enq_req_5_bits_vpu_vta; \
        force U_IF_NAME.io_enq_req_5_bits_vpu_vsew = RTL_PATH.io_enq_req_5_bits_vpu_vsew; \
        force U_IF_NAME.io_enq_req_5_bits_vpu_vlmul = RTL_PATH.io_enq_req_5_bits_vpu_vlmul; \
        force U_IF_NAME.io_enq_req_5_bits_vpu_specVill = RTL_PATH.io_enq_req_5_bits_vpu_specVill; \
        force U_IF_NAME.io_enq_req_5_bits_vpu_specVma = RTL_PATH.io_enq_req_5_bits_vpu_specVma; \
        force U_IF_NAME.io_enq_req_5_bits_vpu_specVta = RTL_PATH.io_enq_req_5_bits_vpu_specVta; \
        force U_IF_NAME.io_enq_req_5_bits_vpu_specVsew = RTL_PATH.io_enq_req_5_bits_vpu_specVsew; \
        force U_IF_NAME.io_enq_req_5_bits_vpu_specVlmul = RTL_PATH.io_enq_req_5_bits_vpu_specVlmul; \
        force U_IF_NAME.io_enq_req_5_bits_vlsInstr = RTL_PATH.io_enq_req_5_bits_vlsInstr; \
        force U_IF_NAME.io_enq_req_5_bits_wfflags = RTL_PATH.io_enq_req_5_bits_wfflags; \
        force U_IF_NAME.io_enq_req_5_bits_isMove = RTL_PATH.io_enq_req_5_bits_isMove; \
        force U_IF_NAME.io_enq_req_5_bits_isVset = RTL_PATH.io_enq_req_5_bits_isVset; \
        force U_IF_NAME.io_enq_req_5_bits_firstUop = RTL_PATH.io_enq_req_5_bits_firstUop; \
        force U_IF_NAME.io_enq_req_5_bits_lastUop = RTL_PATH.io_enq_req_5_bits_lastUop; \
        force U_IF_NAME.io_enq_req_5_bits_numWB = RTL_PATH.io_enq_req_5_bits_numWB; \
        force U_IF_NAME.io_enq_req_5_bits_commitType = RTL_PATH.io_enq_req_5_bits_commitType; \
        force U_IF_NAME.io_enq_req_5_bits_pdest = RTL_PATH.io_enq_req_5_bits_pdest; \
        force U_IF_NAME.io_enq_req_5_bits_robIdx_flag = RTL_PATH.io_enq_req_5_bits_robIdx_flag; \
        force U_IF_NAME.io_enq_req_5_bits_robIdx_value = RTL_PATH.io_enq_req_5_bits_robIdx_value; \
        force U_IF_NAME.io_enq_req_5_bits_instrSize = RTL_PATH.io_enq_req_5_bits_instrSize; \
        force U_IF_NAME.io_enq_req_5_bits_dirtyFs = RTL_PATH.io_enq_req_5_bits_dirtyFs; \
        force U_IF_NAME.io_enq_req_5_bits_dirtyVs = RTL_PATH.io_enq_req_5_bits_dirtyVs; \
        force U_IF_NAME.io_enq_req_5_bits_traceBlockInPipe_itype = RTL_PATH.io_enq_req_5_bits_traceBlockInPipe_itype; \
        force U_IF_NAME.io_enq_req_5_bits_traceBlockInPipe_iretire = RTL_PATH.io_enq_req_5_bits_traceBlockInPipe_iretire; \
        force U_IF_NAME.io_enq_req_5_bits_traceBlockInPipe_ilastsize = RTL_PATH.io_enq_req_5_bits_traceBlockInPipe_ilastsize; \
        force U_IF_NAME.io_enq_req_5_bits_eliminatedMove = RTL_PATH.io_enq_req_5_bits_eliminatedMove; \
        force U_IF_NAME.io_enq_req_5_bits_snapshot = RTL_PATH.io_enq_req_5_bits_snapshot; \
        force U_IF_NAME.io_enq_req_5_bits_lqIdx_value = RTL_PATH.io_enq_req_5_bits_lqIdx_value; \
        force U_IF_NAME.io_enq_req_5_bits_sqIdx_value = RTL_PATH.io_enq_req_5_bits_sqIdx_value; \
        force U_IF_NAME.io_enq_req_5_bits_singleStep = RTL_PATH.io_enq_req_5_bits_singleStep; \
        force U_IF_NAME.io_enq_req_5_bits_debug_sim_trig = RTL_PATH.io_enq_req_5_bits_debug_sim_trig; \
    end \
    `endif

`endif

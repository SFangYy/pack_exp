//=========================================================
//File name    : rename_in_agent_interface.sv
//Author       : nanyunhao
//Module name  : rename_in_agent_interface
//Discribution : rename_in_agent_interface : signal interface
//Date         : 2026-01-22
//=========================================================
`ifndef RENAME_IN_AGENT_INTERFACE__SV
`define RENAME_IN_AGENT_INTERFACE__SV

`ifndef DEF_SETUP_TIME
    `define DEF_SETUP_TIME 1
`endif
`ifndef DEF_HOLD_TIME
    `define DEF_HOLD_TIME 1
`endif

interface rename_in_agent_interface  (input bit clk,input bit rst_n);

    logic         clock                ;
    logic         reset                ;
    logic [5:0]   io_hartId            ;
    logic         io_enq_req_0_valid   ;
    logic [31:0]  io_enq_req_0_bits_instr;
    logic [49:0]  io_enq_req_0_bits_pc ;
    logic         io_enq_req_0_bits_exceptionVec_0;
    logic         io_enq_req_0_bits_exceptionVec_1;
    logic         io_enq_req_0_bits_exceptionVec_2;
    logic         io_enq_req_0_bits_exceptionVec_3;
    logic         io_enq_req_0_bits_exceptionVec_12;
    logic         io_enq_req_0_bits_exceptionVec_20;
    logic         io_enq_req_0_bits_exceptionVec_22;
    logic         io_enq_req_0_bits_isFetchMalAddr;
    logic         io_enq_req_0_bits_hasException;
    logic [3:0]   io_enq_req_0_bits_trigger;
    logic         io_enq_req_0_bits_preDecodeInfo_isRVC;
    logic         io_enq_req_0_bits_crossPageIPFFix;
    logic         io_enq_req_0_bits_ftqPtr_flag;
    logic [5:0]   io_enq_req_0_bits_ftqPtr_value;
    logic [3:0]   io_enq_req_0_bits_ftqOffset;
    logic [5:0]   io_enq_req_0_bits_ldest;
    logic [34:0]  io_enq_req_0_bits_fuType;
    logic [8:0]   io_enq_req_0_bits_fuOpType;
    logic         io_enq_req_0_bits_rfWen;
    logic         io_enq_req_0_bits_fpWen;
    logic         io_enq_req_0_bits_vecWen;
    logic         io_enq_req_0_bits_v0Wen;
    logic         io_enq_req_0_bits_vlWen;
    logic         io_enq_req_0_bits_isXSTrap;
    logic         io_enq_req_0_bits_waitForward;
    logic         io_enq_req_0_bits_blockBackward;
    logic         io_enq_req_0_bits_flushPipe;
    logic         io_enq_req_0_bits_vpu_vill;
    logic         io_enq_req_0_bits_vpu_vma;
    logic         io_enq_req_0_bits_vpu_vta;
    logic [1:0]   io_enq_req_0_bits_vpu_vsew;
    logic [2:0]   io_enq_req_0_bits_vpu_vlmul;
    logic         io_enq_req_0_bits_vpu_specVill;
    logic         io_enq_req_0_bits_vpu_specVma;
    logic         io_enq_req_0_bits_vpu_specVta;
    logic [1:0]   io_enq_req_0_bits_vpu_specVsew;
    logic [2:0]   io_enq_req_0_bits_vpu_specVlmul;
    logic         io_enq_req_0_bits_vlsInstr;
    logic         io_enq_req_0_bits_wfflags;
    logic         io_enq_req_0_bits_isMove;
    logic         io_enq_req_0_bits_isVset;
    logic         io_enq_req_0_bits_firstUop;
    logic         io_enq_req_0_bits_lastUop;
    logic [6:0]   io_enq_req_0_bits_numWB;
    logic [2:0]   io_enq_req_0_bits_commitType;
    logic [7:0]   io_enq_req_0_bits_pdest;
    logic         io_enq_req_0_bits_robIdx_flag;
    logic [7:0]   io_enq_req_0_bits_robIdx_value;
    logic [2:0]   io_enq_req_0_bits_instrSize;
    logic         io_enq_req_0_bits_dirtyFs;
    logic         io_enq_req_0_bits_dirtyVs;
    logic [3:0]   io_enq_req_0_bits_traceBlockInPipe_itype;
    logic [3:0]   io_enq_req_0_bits_traceBlockInPipe_iretire;
    logic         io_enq_req_0_bits_traceBlockInPipe_ilastsize;
    logic         io_enq_req_0_bits_eliminatedMove;
    logic         io_enq_req_0_bits_snapshot;
    logic [6:0]   io_enq_req_0_bits_lqIdx_value;
    logic [5:0]   io_enq_req_0_bits_sqIdx_value;
    logic         io_enq_req_0_bits_singleStep;
    logic         io_enq_req_0_bits_debug_sim_trig;
    logic         io_enq_req_1_valid   ;
    logic [31:0]  io_enq_req_1_bits_instr;
    logic [49:0]  io_enq_req_1_bits_pc ;
    logic         io_enq_req_1_bits_exceptionVec_0;
    logic         io_enq_req_1_bits_exceptionVec_1;
    logic         io_enq_req_1_bits_exceptionVec_2;
    logic         io_enq_req_1_bits_exceptionVec_3;
    logic         io_enq_req_1_bits_exceptionVec_12;
    logic         io_enq_req_1_bits_exceptionVec_20;
    logic         io_enq_req_1_bits_exceptionVec_22;
    logic         io_enq_req_1_bits_isFetchMalAddr;
    logic         io_enq_req_1_bits_hasException;
    logic [3:0]   io_enq_req_1_bits_trigger;
    logic         io_enq_req_1_bits_preDecodeInfo_isRVC;
    logic         io_enq_req_1_bits_crossPageIPFFix;
    logic         io_enq_req_1_bits_ftqPtr_flag;
    logic [5:0]   io_enq_req_1_bits_ftqPtr_value;
    logic [3:0]   io_enq_req_1_bits_ftqOffset;
    logic [5:0]   io_enq_req_1_bits_ldest;
    logic [34:0]  io_enq_req_1_bits_fuType;
    logic [8:0]   io_enq_req_1_bits_fuOpType;
    logic         io_enq_req_1_bits_rfWen;
    logic         io_enq_req_1_bits_fpWen;
    logic         io_enq_req_1_bits_vecWen;
    logic         io_enq_req_1_bits_v0Wen;
    logic         io_enq_req_1_bits_vlWen;
    logic         io_enq_req_1_bits_isXSTrap;
    logic         io_enq_req_1_bits_waitForward;
    logic         io_enq_req_1_bits_blockBackward;
    logic         io_enq_req_1_bits_flushPipe;
    logic         io_enq_req_1_bits_vpu_vill;
    logic         io_enq_req_1_bits_vpu_vma;
    logic         io_enq_req_1_bits_vpu_vta;
    logic [1:0]   io_enq_req_1_bits_vpu_vsew;
    logic [2:0]   io_enq_req_1_bits_vpu_vlmul;
    logic         io_enq_req_1_bits_vpu_specVill;
    logic         io_enq_req_1_bits_vpu_specVma;
    logic         io_enq_req_1_bits_vpu_specVta;
    logic [1:0]   io_enq_req_1_bits_vpu_specVsew;
    logic [2:0]   io_enq_req_1_bits_vpu_specVlmul;
    logic         io_enq_req_1_bits_vlsInstr;
    logic         io_enq_req_1_bits_wfflags;
    logic         io_enq_req_1_bits_isMove;
    logic         io_enq_req_1_bits_isVset;
    logic         io_enq_req_1_bits_firstUop;
    logic         io_enq_req_1_bits_lastUop;
    logic [6:0]   io_enq_req_1_bits_numWB;
    logic [2:0]   io_enq_req_1_bits_commitType;
    logic [7:0]   io_enq_req_1_bits_pdest;
    logic         io_enq_req_1_bits_robIdx_flag;
    logic [7:0]   io_enq_req_1_bits_robIdx_value;
    logic [2:0]   io_enq_req_1_bits_instrSize;
    logic         io_enq_req_1_bits_dirtyFs;
    logic         io_enq_req_1_bits_dirtyVs;
    logic [3:0]   io_enq_req_1_bits_traceBlockInPipe_itype;
    logic [3:0]   io_enq_req_1_bits_traceBlockInPipe_iretire;
    logic         io_enq_req_1_bits_traceBlockInPipe_ilastsize;
    logic         io_enq_req_1_bits_eliminatedMove;
    logic         io_enq_req_1_bits_snapshot;
    logic [6:0]   io_enq_req_1_bits_lqIdx_value;
    logic [5:0]   io_enq_req_1_bits_sqIdx_value;
    logic         io_enq_req_1_bits_singleStep;
    logic         io_enq_req_1_bits_debug_sim_trig;
    logic         io_enq_req_2_valid   ;
    logic [31:0]  io_enq_req_2_bits_instr;
    logic [49:0]  io_enq_req_2_bits_pc ;
    logic         io_enq_req_2_bits_exceptionVec_0;
    logic         io_enq_req_2_bits_exceptionVec_1;
    logic         io_enq_req_2_bits_exceptionVec_2;
    logic         io_enq_req_2_bits_exceptionVec_3;
    logic         io_enq_req_2_bits_exceptionVec_12;
    logic         io_enq_req_2_bits_exceptionVec_20;
    logic         io_enq_req_2_bits_exceptionVec_22;
    logic         io_enq_req_2_bits_isFetchMalAddr;
    logic         io_enq_req_2_bits_hasException;
    logic [3:0]   io_enq_req_2_bits_trigger;
    logic         io_enq_req_2_bits_preDecodeInfo_isRVC;
    logic         io_enq_req_2_bits_crossPageIPFFix;
    logic         io_enq_req_2_bits_ftqPtr_flag;
    logic [5:0]   io_enq_req_2_bits_ftqPtr_value;
    logic [3:0]   io_enq_req_2_bits_ftqOffset;
    logic [5:0]   io_enq_req_2_bits_ldest;
    logic [34:0]  io_enq_req_2_bits_fuType;
    logic [8:0]   io_enq_req_2_bits_fuOpType;
    logic         io_enq_req_2_bits_rfWen;
    logic         io_enq_req_2_bits_fpWen;
    logic         io_enq_req_2_bits_vecWen;
    logic         io_enq_req_2_bits_v0Wen;
    logic         io_enq_req_2_bits_vlWen;
    logic         io_enq_req_2_bits_isXSTrap;
    logic         io_enq_req_2_bits_waitForward;
    logic         io_enq_req_2_bits_blockBackward;
    logic         io_enq_req_2_bits_flushPipe;
    logic         io_enq_req_2_bits_vpu_vill;
    logic         io_enq_req_2_bits_vpu_vma;
    logic         io_enq_req_2_bits_vpu_vta;
    logic [1:0]   io_enq_req_2_bits_vpu_vsew;
    logic [2:0]   io_enq_req_2_bits_vpu_vlmul;
    logic         io_enq_req_2_bits_vpu_specVill;
    logic         io_enq_req_2_bits_vpu_specVma;
    logic         io_enq_req_2_bits_vpu_specVta;
    logic [1:0]   io_enq_req_2_bits_vpu_specVsew;
    logic [2:0]   io_enq_req_2_bits_vpu_specVlmul;
    logic         io_enq_req_2_bits_vlsInstr;
    logic         io_enq_req_2_bits_wfflags;
    logic         io_enq_req_2_bits_isMove;
    logic         io_enq_req_2_bits_isVset;
    logic         io_enq_req_2_bits_firstUop;
    logic         io_enq_req_2_bits_lastUop;
    logic [6:0]   io_enq_req_2_bits_numWB;
    logic [2:0]   io_enq_req_2_bits_commitType;
    logic [7:0]   io_enq_req_2_bits_pdest;
    logic         io_enq_req_2_bits_robIdx_flag;
    logic [7:0]   io_enq_req_2_bits_robIdx_value;
    logic [2:0]   io_enq_req_2_bits_instrSize;
    logic         io_enq_req_2_bits_dirtyFs;
    logic         io_enq_req_2_bits_dirtyVs;
    logic [3:0]   io_enq_req_2_bits_traceBlockInPipe_itype;
    logic [3:0]   io_enq_req_2_bits_traceBlockInPipe_iretire;
    logic         io_enq_req_2_bits_traceBlockInPipe_ilastsize;
    logic         io_enq_req_2_bits_eliminatedMove;
    logic         io_enq_req_2_bits_snapshot;
    logic [6:0]   io_enq_req_2_bits_lqIdx_value;
    logic [5:0]   io_enq_req_2_bits_sqIdx_value;
    logic         io_enq_req_2_bits_singleStep;
    logic         io_enq_req_2_bits_debug_sim_trig;
    logic         io_enq_req_3_valid   ;
    logic [31:0]  io_enq_req_3_bits_instr;
    logic [49:0]  io_enq_req_3_bits_pc ;
    logic         io_enq_req_3_bits_exceptionVec_0;
    logic         io_enq_req_3_bits_exceptionVec_1;
    logic         io_enq_req_3_bits_exceptionVec_2;
    logic         io_enq_req_3_bits_exceptionVec_3;
    logic         io_enq_req_3_bits_exceptionVec_12;
    logic         io_enq_req_3_bits_exceptionVec_20;
    logic         io_enq_req_3_bits_exceptionVec_22;
    logic         io_enq_req_3_bits_isFetchMalAddr;
    logic         io_enq_req_3_bits_hasException;
    logic [3:0]   io_enq_req_3_bits_trigger;
    logic         io_enq_req_3_bits_preDecodeInfo_isRVC;
    logic         io_enq_req_3_bits_crossPageIPFFix;
    logic         io_enq_req_3_bits_ftqPtr_flag;
    logic [5:0]   io_enq_req_3_bits_ftqPtr_value;
    logic [3:0]   io_enq_req_3_bits_ftqOffset;
    logic [5:0]   io_enq_req_3_bits_ldest;
    logic [34:0]  io_enq_req_3_bits_fuType;
    logic [8:0]   io_enq_req_3_bits_fuOpType;
    logic         io_enq_req_3_bits_rfWen;
    logic         io_enq_req_3_bits_fpWen;
    logic         io_enq_req_3_bits_vecWen;
    logic         io_enq_req_3_bits_v0Wen;
    logic         io_enq_req_3_bits_vlWen;
    logic         io_enq_req_3_bits_isXSTrap;
    logic         io_enq_req_3_bits_waitForward;
    logic         io_enq_req_3_bits_blockBackward;
    logic         io_enq_req_3_bits_flushPipe;
    logic         io_enq_req_3_bits_vpu_vill;
    logic         io_enq_req_3_bits_vpu_vma;
    logic         io_enq_req_3_bits_vpu_vta;
    logic [1:0]   io_enq_req_3_bits_vpu_vsew;
    logic [2:0]   io_enq_req_3_bits_vpu_vlmul;
    logic         io_enq_req_3_bits_vpu_specVill;
    logic         io_enq_req_3_bits_vpu_specVma;
    logic         io_enq_req_3_bits_vpu_specVta;
    logic [1:0]   io_enq_req_3_bits_vpu_specVsew;
    logic [2:0]   io_enq_req_3_bits_vpu_specVlmul;
    logic         io_enq_req_3_bits_vlsInstr;
    logic         io_enq_req_3_bits_wfflags;
    logic         io_enq_req_3_bits_isMove;
    logic         io_enq_req_3_bits_isVset;
    logic         io_enq_req_3_bits_firstUop;
    logic         io_enq_req_3_bits_lastUop;
    logic [6:0]   io_enq_req_3_bits_numWB;
    logic [2:0]   io_enq_req_3_bits_commitType;
    logic [7:0]   io_enq_req_3_bits_pdest;
    logic         io_enq_req_3_bits_robIdx_flag;
    logic [7:0]   io_enq_req_3_bits_robIdx_value;
    logic [2:0]   io_enq_req_3_bits_instrSize;
    logic         io_enq_req_3_bits_dirtyFs;
    logic         io_enq_req_3_bits_dirtyVs;
    logic [3:0]   io_enq_req_3_bits_traceBlockInPipe_itype;
    logic [3:0]   io_enq_req_3_bits_traceBlockInPipe_iretire;
    logic         io_enq_req_3_bits_traceBlockInPipe_ilastsize;
    logic         io_enq_req_3_bits_eliminatedMove;
    logic         io_enq_req_3_bits_snapshot;
    logic [6:0]   io_enq_req_3_bits_lqIdx_value;
    logic [5:0]   io_enq_req_3_bits_sqIdx_value;
    logic         io_enq_req_3_bits_singleStep;
    logic         io_enq_req_3_bits_debug_sim_trig;
    logic         io_enq_req_4_valid   ;
    logic [31:0]  io_enq_req_4_bits_instr;
    logic [49:0]  io_enq_req_4_bits_pc ;
    logic         io_enq_req_4_bits_exceptionVec_0;
    logic         io_enq_req_4_bits_exceptionVec_1;
    logic         io_enq_req_4_bits_exceptionVec_2;
    logic         io_enq_req_4_bits_exceptionVec_3;
    logic         io_enq_req_4_bits_exceptionVec_12;
    logic         io_enq_req_4_bits_exceptionVec_20;
    logic         io_enq_req_4_bits_exceptionVec_22;
    logic         io_enq_req_4_bits_isFetchMalAddr;
    logic         io_enq_req_4_bits_hasException;
    logic [3:0]   io_enq_req_4_bits_trigger;
    logic         io_enq_req_4_bits_preDecodeInfo_isRVC;
    logic         io_enq_req_4_bits_crossPageIPFFix;
    logic         io_enq_req_4_bits_ftqPtr_flag;
    logic [5:0]   io_enq_req_4_bits_ftqPtr_value;
    logic [3:0]   io_enq_req_4_bits_ftqOffset;
    logic [5:0]   io_enq_req_4_bits_ldest;
    logic [34:0]  io_enq_req_4_bits_fuType;
    logic [8:0]   io_enq_req_4_bits_fuOpType;
    logic         io_enq_req_4_bits_rfWen;
    logic         io_enq_req_4_bits_fpWen;
    logic         io_enq_req_4_bits_vecWen;
    logic         io_enq_req_4_bits_v0Wen;
    logic         io_enq_req_4_bits_vlWen;
    logic         io_enq_req_4_bits_isXSTrap;
    logic         io_enq_req_4_bits_waitForward;
    logic         io_enq_req_4_bits_blockBackward;
    logic         io_enq_req_4_bits_flushPipe;
    logic         io_enq_req_4_bits_vpu_vill;
    logic         io_enq_req_4_bits_vpu_vma;
    logic         io_enq_req_4_bits_vpu_vta;
    logic [1:0]   io_enq_req_4_bits_vpu_vsew;
    logic [2:0]   io_enq_req_4_bits_vpu_vlmul;
    logic         io_enq_req_4_bits_vpu_specVill;
    logic         io_enq_req_4_bits_vpu_specVma;
    logic         io_enq_req_4_bits_vpu_specVta;
    logic [1:0]   io_enq_req_4_bits_vpu_specVsew;
    logic [2:0]   io_enq_req_4_bits_vpu_specVlmul;
    logic         io_enq_req_4_bits_vlsInstr;
    logic         io_enq_req_4_bits_wfflags;
    logic         io_enq_req_4_bits_isMove;
    logic         io_enq_req_4_bits_isVset;
    logic         io_enq_req_4_bits_firstUop;
    logic         io_enq_req_4_bits_lastUop;
    logic [6:0]   io_enq_req_4_bits_numWB;
    logic [2:0]   io_enq_req_4_bits_commitType;
    logic [7:0]   io_enq_req_4_bits_pdest;
    logic         io_enq_req_4_bits_robIdx_flag;
    logic [7:0]   io_enq_req_4_bits_robIdx_value;
    logic [2:0]   io_enq_req_4_bits_instrSize;
    logic         io_enq_req_4_bits_dirtyFs;
    logic         io_enq_req_4_bits_dirtyVs;
    logic [3:0]   io_enq_req_4_bits_traceBlockInPipe_itype;
    logic [3:0]   io_enq_req_4_bits_traceBlockInPipe_iretire;
    logic         io_enq_req_4_bits_traceBlockInPipe_ilastsize;
    logic         io_enq_req_4_bits_eliminatedMove;
    logic         io_enq_req_4_bits_snapshot;
    logic [6:0]   io_enq_req_4_bits_lqIdx_value;
    logic [5:0]   io_enq_req_4_bits_sqIdx_value;
    logic         io_enq_req_4_bits_singleStep;
    logic         io_enq_req_4_bits_debug_sim_trig;
    logic         io_enq_req_5_valid   ;
    logic [31:0]  io_enq_req_5_bits_instr;
    logic [49:0]  io_enq_req_5_bits_pc ;
    logic         io_enq_req_5_bits_exceptionVec_0;
    logic         io_enq_req_5_bits_exceptionVec_1;
    logic         io_enq_req_5_bits_exceptionVec_2;
    logic         io_enq_req_5_bits_exceptionVec_3;
    logic         io_enq_req_5_bits_exceptionVec_12;
    logic         io_enq_req_5_bits_exceptionVec_20;
    logic         io_enq_req_5_bits_exceptionVec_22;
    logic         io_enq_req_5_bits_isFetchMalAddr;
    logic         io_enq_req_5_bits_hasException;
    logic [3:0]   io_enq_req_5_bits_trigger;
    logic         io_enq_req_5_bits_preDecodeInfo_isRVC;
    logic         io_enq_req_5_bits_crossPageIPFFix;
    logic         io_enq_req_5_bits_ftqPtr_flag;
    logic [5:0]   io_enq_req_5_bits_ftqPtr_value;
    logic [3:0]   io_enq_req_5_bits_ftqOffset;
    logic [5:0]   io_enq_req_5_bits_ldest;
    logic [34:0]  io_enq_req_5_bits_fuType;
    logic [8:0]   io_enq_req_5_bits_fuOpType;
    logic         io_enq_req_5_bits_rfWen;
    logic         io_enq_req_5_bits_fpWen;
    logic         io_enq_req_5_bits_vecWen;
    logic         io_enq_req_5_bits_v0Wen;
    logic         io_enq_req_5_bits_vlWen;
    logic         io_enq_req_5_bits_isXSTrap;
    logic         io_enq_req_5_bits_waitForward;
    logic         io_enq_req_5_bits_blockBackward;
    logic         io_enq_req_5_bits_flushPipe;
    logic         io_enq_req_5_bits_vpu_vill;
    logic         io_enq_req_5_bits_vpu_vma;
    logic         io_enq_req_5_bits_vpu_vta;
    logic [1:0]   io_enq_req_5_bits_vpu_vsew;
    logic [2:0]   io_enq_req_5_bits_vpu_vlmul;
    logic         io_enq_req_5_bits_vpu_specVill;
    logic         io_enq_req_5_bits_vpu_specVma;
    logic         io_enq_req_5_bits_vpu_specVta;
    logic [1:0]   io_enq_req_5_bits_vpu_specVsew;
    logic [2:0]   io_enq_req_5_bits_vpu_specVlmul;
    logic         io_enq_req_5_bits_vlsInstr;
    logic         io_enq_req_5_bits_wfflags;
    logic         io_enq_req_5_bits_isMove;
    logic         io_enq_req_5_bits_isVset;
    logic         io_enq_req_5_bits_firstUop;
    logic         io_enq_req_5_bits_lastUop;
    logic [6:0]   io_enq_req_5_bits_numWB;
    logic [2:0]   io_enq_req_5_bits_commitType;
    logic [7:0]   io_enq_req_5_bits_pdest;
    logic         io_enq_req_5_bits_robIdx_flag;
    logic [7:0]   io_enq_req_5_bits_robIdx_value;
    logic [2:0]   io_enq_req_5_bits_instrSize;
    logic         io_enq_req_5_bits_dirtyFs;
    logic         io_enq_req_5_bits_dirtyVs;
    logic [3:0]   io_enq_req_5_bits_traceBlockInPipe_itype;
    logic [3:0]   io_enq_req_5_bits_traceBlockInPipe_iretire;
    logic         io_enq_req_5_bits_traceBlockInPipe_ilastsize;
    logic         io_enq_req_5_bits_eliminatedMove;
    logic         io_enq_req_5_bits_snapshot;
    logic [6:0]   io_enq_req_5_bits_lqIdx_value;
    logic [5:0]   io_enq_req_5_bits_sqIdx_value;
    logic         io_enq_req_5_bits_singleStep;
    logic         io_enq_req_5_bits_debug_sim_trig;

    clocking drv_cb @(posedge clk);
        `ifdef INTERFACE_ADD_DELAY
            default input #`DEF_SETUP_TIME output #`DEF_HOLD_TIME;
        `endif
        output clock;
        output reset;
        output io_hartId;
        output io_enq_req_0_valid;
        output io_enq_req_0_bits_instr;
        output io_enq_req_0_bits_pc;
        output io_enq_req_0_bits_exceptionVec_0;
        output io_enq_req_0_bits_exceptionVec_1;
        output io_enq_req_0_bits_exceptionVec_2;
        output io_enq_req_0_bits_exceptionVec_3;
        output io_enq_req_0_bits_exceptionVec_12;
        output io_enq_req_0_bits_exceptionVec_20;
        output io_enq_req_0_bits_exceptionVec_22;
        output io_enq_req_0_bits_isFetchMalAddr;
        output io_enq_req_0_bits_hasException;
        output io_enq_req_0_bits_trigger;
        output io_enq_req_0_bits_preDecodeInfo_isRVC;
        output io_enq_req_0_bits_crossPageIPFFix;
        output io_enq_req_0_bits_ftqPtr_flag;
        output io_enq_req_0_bits_ftqPtr_value;
        output io_enq_req_0_bits_ftqOffset;
        output io_enq_req_0_bits_ldest;
        output io_enq_req_0_bits_fuType;
        output io_enq_req_0_bits_fuOpType;
        output io_enq_req_0_bits_rfWen;
        output io_enq_req_0_bits_fpWen;
        output io_enq_req_0_bits_vecWen;
        output io_enq_req_0_bits_v0Wen;
        output io_enq_req_0_bits_vlWen;
        output io_enq_req_0_bits_isXSTrap;
        output io_enq_req_0_bits_waitForward;
        output io_enq_req_0_bits_blockBackward;
        output io_enq_req_0_bits_flushPipe;
        output io_enq_req_0_bits_vpu_vill;
        output io_enq_req_0_bits_vpu_vma;
        output io_enq_req_0_bits_vpu_vta;
        output io_enq_req_0_bits_vpu_vsew;
        output io_enq_req_0_bits_vpu_vlmul;
        output io_enq_req_0_bits_vpu_specVill;
        output io_enq_req_0_bits_vpu_specVma;
        output io_enq_req_0_bits_vpu_specVta;
        output io_enq_req_0_bits_vpu_specVsew;
        output io_enq_req_0_bits_vpu_specVlmul;
        output io_enq_req_0_bits_vlsInstr;
        output io_enq_req_0_bits_wfflags;
        output io_enq_req_0_bits_isMove;
        output io_enq_req_0_bits_isVset;
        output io_enq_req_0_bits_firstUop;
        output io_enq_req_0_bits_lastUop;
        output io_enq_req_0_bits_numWB;
        output io_enq_req_0_bits_commitType;
        output io_enq_req_0_bits_pdest;
        output io_enq_req_0_bits_robIdx_flag;
        output io_enq_req_0_bits_robIdx_value;
        output io_enq_req_0_bits_instrSize;
        output io_enq_req_0_bits_dirtyFs;
        output io_enq_req_0_bits_dirtyVs;
        output io_enq_req_0_bits_traceBlockInPipe_itype;
        output io_enq_req_0_bits_traceBlockInPipe_iretire;
        output io_enq_req_0_bits_traceBlockInPipe_ilastsize;
        output io_enq_req_0_bits_eliminatedMove;
        output io_enq_req_0_bits_snapshot;
        output io_enq_req_0_bits_lqIdx_value;
        output io_enq_req_0_bits_sqIdx_value;
        output io_enq_req_0_bits_singleStep;
        output io_enq_req_0_bits_debug_sim_trig;
        output io_enq_req_1_valid;
        output io_enq_req_1_bits_instr;
        output io_enq_req_1_bits_pc;
        output io_enq_req_1_bits_exceptionVec_0;
        output io_enq_req_1_bits_exceptionVec_1;
        output io_enq_req_1_bits_exceptionVec_2;
        output io_enq_req_1_bits_exceptionVec_3;
        output io_enq_req_1_bits_exceptionVec_12;
        output io_enq_req_1_bits_exceptionVec_20;
        output io_enq_req_1_bits_exceptionVec_22;
        output io_enq_req_1_bits_isFetchMalAddr;
        output io_enq_req_1_bits_hasException;
        output io_enq_req_1_bits_trigger;
        output io_enq_req_1_bits_preDecodeInfo_isRVC;
        output io_enq_req_1_bits_crossPageIPFFix;
        output io_enq_req_1_bits_ftqPtr_flag;
        output io_enq_req_1_bits_ftqPtr_value;
        output io_enq_req_1_bits_ftqOffset;
        output io_enq_req_1_bits_ldest;
        output io_enq_req_1_bits_fuType;
        output io_enq_req_1_bits_fuOpType;
        output io_enq_req_1_bits_rfWen;
        output io_enq_req_1_bits_fpWen;
        output io_enq_req_1_bits_vecWen;
        output io_enq_req_1_bits_v0Wen;
        output io_enq_req_1_bits_vlWen;
        output io_enq_req_1_bits_isXSTrap;
        output io_enq_req_1_bits_waitForward;
        output io_enq_req_1_bits_blockBackward;
        output io_enq_req_1_bits_flushPipe;
        output io_enq_req_1_bits_vpu_vill;
        output io_enq_req_1_bits_vpu_vma;
        output io_enq_req_1_bits_vpu_vta;
        output io_enq_req_1_bits_vpu_vsew;
        output io_enq_req_1_bits_vpu_vlmul;
        output io_enq_req_1_bits_vpu_specVill;
        output io_enq_req_1_bits_vpu_specVma;
        output io_enq_req_1_bits_vpu_specVta;
        output io_enq_req_1_bits_vpu_specVsew;
        output io_enq_req_1_bits_vpu_specVlmul;
        output io_enq_req_1_bits_vlsInstr;
        output io_enq_req_1_bits_wfflags;
        output io_enq_req_1_bits_isMove;
        output io_enq_req_1_bits_isVset;
        output io_enq_req_1_bits_firstUop;
        output io_enq_req_1_bits_lastUop;
        output io_enq_req_1_bits_numWB;
        output io_enq_req_1_bits_commitType;
        output io_enq_req_1_bits_pdest;
        output io_enq_req_1_bits_robIdx_flag;
        output io_enq_req_1_bits_robIdx_value;
        output io_enq_req_1_bits_instrSize;
        output io_enq_req_1_bits_dirtyFs;
        output io_enq_req_1_bits_dirtyVs;
        output io_enq_req_1_bits_traceBlockInPipe_itype;
        output io_enq_req_1_bits_traceBlockInPipe_iretire;
        output io_enq_req_1_bits_traceBlockInPipe_ilastsize;
        output io_enq_req_1_bits_eliminatedMove;
        output io_enq_req_1_bits_snapshot;
        output io_enq_req_1_bits_lqIdx_value;
        output io_enq_req_1_bits_sqIdx_value;
        output io_enq_req_1_bits_singleStep;
        output io_enq_req_1_bits_debug_sim_trig;
        output io_enq_req_2_valid;
        output io_enq_req_2_bits_instr;
        output io_enq_req_2_bits_pc;
        output io_enq_req_2_bits_exceptionVec_0;
        output io_enq_req_2_bits_exceptionVec_1;
        output io_enq_req_2_bits_exceptionVec_2;
        output io_enq_req_2_bits_exceptionVec_3;
        output io_enq_req_2_bits_exceptionVec_12;
        output io_enq_req_2_bits_exceptionVec_20;
        output io_enq_req_2_bits_exceptionVec_22;
        output io_enq_req_2_bits_isFetchMalAddr;
        output io_enq_req_2_bits_hasException;
        output io_enq_req_2_bits_trigger;
        output io_enq_req_2_bits_preDecodeInfo_isRVC;
        output io_enq_req_2_bits_crossPageIPFFix;
        output io_enq_req_2_bits_ftqPtr_flag;
        output io_enq_req_2_bits_ftqPtr_value;
        output io_enq_req_2_bits_ftqOffset;
        output io_enq_req_2_bits_ldest;
        output io_enq_req_2_bits_fuType;
        output io_enq_req_2_bits_fuOpType;
        output io_enq_req_2_bits_rfWen;
        output io_enq_req_2_bits_fpWen;
        output io_enq_req_2_bits_vecWen;
        output io_enq_req_2_bits_v0Wen;
        output io_enq_req_2_bits_vlWen;
        output io_enq_req_2_bits_isXSTrap;
        output io_enq_req_2_bits_waitForward;
        output io_enq_req_2_bits_blockBackward;
        output io_enq_req_2_bits_flushPipe;
        output io_enq_req_2_bits_vpu_vill;
        output io_enq_req_2_bits_vpu_vma;
        output io_enq_req_2_bits_vpu_vta;
        output io_enq_req_2_bits_vpu_vsew;
        output io_enq_req_2_bits_vpu_vlmul;
        output io_enq_req_2_bits_vpu_specVill;
        output io_enq_req_2_bits_vpu_specVma;
        output io_enq_req_2_bits_vpu_specVta;
        output io_enq_req_2_bits_vpu_specVsew;
        output io_enq_req_2_bits_vpu_specVlmul;
        output io_enq_req_2_bits_vlsInstr;
        output io_enq_req_2_bits_wfflags;
        output io_enq_req_2_bits_isMove;
        output io_enq_req_2_bits_isVset;
        output io_enq_req_2_bits_firstUop;
        output io_enq_req_2_bits_lastUop;
        output io_enq_req_2_bits_numWB;
        output io_enq_req_2_bits_commitType;
        output io_enq_req_2_bits_pdest;
        output io_enq_req_2_bits_robIdx_flag;
        output io_enq_req_2_bits_robIdx_value;
        output io_enq_req_2_bits_instrSize;
        output io_enq_req_2_bits_dirtyFs;
        output io_enq_req_2_bits_dirtyVs;
        output io_enq_req_2_bits_traceBlockInPipe_itype;
        output io_enq_req_2_bits_traceBlockInPipe_iretire;
        output io_enq_req_2_bits_traceBlockInPipe_ilastsize;
        output io_enq_req_2_bits_eliminatedMove;
        output io_enq_req_2_bits_snapshot;
        output io_enq_req_2_bits_lqIdx_value;
        output io_enq_req_2_bits_sqIdx_value;
        output io_enq_req_2_bits_singleStep;
        output io_enq_req_2_bits_debug_sim_trig;
        output io_enq_req_3_valid;
        output io_enq_req_3_bits_instr;
        output io_enq_req_3_bits_pc;
        output io_enq_req_3_bits_exceptionVec_0;
        output io_enq_req_3_bits_exceptionVec_1;
        output io_enq_req_3_bits_exceptionVec_2;
        output io_enq_req_3_bits_exceptionVec_3;
        output io_enq_req_3_bits_exceptionVec_12;
        output io_enq_req_3_bits_exceptionVec_20;
        output io_enq_req_3_bits_exceptionVec_22;
        output io_enq_req_3_bits_isFetchMalAddr;
        output io_enq_req_3_bits_hasException;
        output io_enq_req_3_bits_trigger;
        output io_enq_req_3_bits_preDecodeInfo_isRVC;
        output io_enq_req_3_bits_crossPageIPFFix;
        output io_enq_req_3_bits_ftqPtr_flag;
        output io_enq_req_3_bits_ftqPtr_value;
        output io_enq_req_3_bits_ftqOffset;
        output io_enq_req_3_bits_ldest;
        output io_enq_req_3_bits_fuType;
        output io_enq_req_3_bits_fuOpType;
        output io_enq_req_3_bits_rfWen;
        output io_enq_req_3_bits_fpWen;
        output io_enq_req_3_bits_vecWen;
        output io_enq_req_3_bits_v0Wen;
        output io_enq_req_3_bits_vlWen;
        output io_enq_req_3_bits_isXSTrap;
        output io_enq_req_3_bits_waitForward;
        output io_enq_req_3_bits_blockBackward;
        output io_enq_req_3_bits_flushPipe;
        output io_enq_req_3_bits_vpu_vill;
        output io_enq_req_3_bits_vpu_vma;
        output io_enq_req_3_bits_vpu_vta;
        output io_enq_req_3_bits_vpu_vsew;
        output io_enq_req_3_bits_vpu_vlmul;
        output io_enq_req_3_bits_vpu_specVill;
        output io_enq_req_3_bits_vpu_specVma;
        output io_enq_req_3_bits_vpu_specVta;
        output io_enq_req_3_bits_vpu_specVsew;
        output io_enq_req_3_bits_vpu_specVlmul;
        output io_enq_req_3_bits_vlsInstr;
        output io_enq_req_3_bits_wfflags;
        output io_enq_req_3_bits_isMove;
        output io_enq_req_3_bits_isVset;
        output io_enq_req_3_bits_firstUop;
        output io_enq_req_3_bits_lastUop;
        output io_enq_req_3_bits_numWB;
        output io_enq_req_3_bits_commitType;
        output io_enq_req_3_bits_pdest;
        output io_enq_req_3_bits_robIdx_flag;
        output io_enq_req_3_bits_robIdx_value;
        output io_enq_req_3_bits_instrSize;
        output io_enq_req_3_bits_dirtyFs;
        output io_enq_req_3_bits_dirtyVs;
        output io_enq_req_3_bits_traceBlockInPipe_itype;
        output io_enq_req_3_bits_traceBlockInPipe_iretire;
        output io_enq_req_3_bits_traceBlockInPipe_ilastsize;
        output io_enq_req_3_bits_eliminatedMove;
        output io_enq_req_3_bits_snapshot;
        output io_enq_req_3_bits_lqIdx_value;
        output io_enq_req_3_bits_sqIdx_value;
        output io_enq_req_3_bits_singleStep;
        output io_enq_req_3_bits_debug_sim_trig;
        output io_enq_req_4_valid;
        output io_enq_req_4_bits_instr;
        output io_enq_req_4_bits_pc;
        output io_enq_req_4_bits_exceptionVec_0;
        output io_enq_req_4_bits_exceptionVec_1;
        output io_enq_req_4_bits_exceptionVec_2;
        output io_enq_req_4_bits_exceptionVec_3;
        output io_enq_req_4_bits_exceptionVec_12;
        output io_enq_req_4_bits_exceptionVec_20;
        output io_enq_req_4_bits_exceptionVec_22;
        output io_enq_req_4_bits_isFetchMalAddr;
        output io_enq_req_4_bits_hasException;
        output io_enq_req_4_bits_trigger;
        output io_enq_req_4_bits_preDecodeInfo_isRVC;
        output io_enq_req_4_bits_crossPageIPFFix;
        output io_enq_req_4_bits_ftqPtr_flag;
        output io_enq_req_4_bits_ftqPtr_value;
        output io_enq_req_4_bits_ftqOffset;
        output io_enq_req_4_bits_ldest;
        output io_enq_req_4_bits_fuType;
        output io_enq_req_4_bits_fuOpType;
        output io_enq_req_4_bits_rfWen;
        output io_enq_req_4_bits_fpWen;
        output io_enq_req_4_bits_vecWen;
        output io_enq_req_4_bits_v0Wen;
        output io_enq_req_4_bits_vlWen;
        output io_enq_req_4_bits_isXSTrap;
        output io_enq_req_4_bits_waitForward;
        output io_enq_req_4_bits_blockBackward;
        output io_enq_req_4_bits_flushPipe;
        output io_enq_req_4_bits_vpu_vill;
        output io_enq_req_4_bits_vpu_vma;
        output io_enq_req_4_bits_vpu_vta;
        output io_enq_req_4_bits_vpu_vsew;
        output io_enq_req_4_bits_vpu_vlmul;
        output io_enq_req_4_bits_vpu_specVill;
        output io_enq_req_4_bits_vpu_specVma;
        output io_enq_req_4_bits_vpu_specVta;
        output io_enq_req_4_bits_vpu_specVsew;
        output io_enq_req_4_bits_vpu_specVlmul;
        output io_enq_req_4_bits_vlsInstr;
        output io_enq_req_4_bits_wfflags;
        output io_enq_req_4_bits_isMove;
        output io_enq_req_4_bits_isVset;
        output io_enq_req_4_bits_firstUop;
        output io_enq_req_4_bits_lastUop;
        output io_enq_req_4_bits_numWB;
        output io_enq_req_4_bits_commitType;
        output io_enq_req_4_bits_pdest;
        output io_enq_req_4_bits_robIdx_flag;
        output io_enq_req_4_bits_robIdx_value;
        output io_enq_req_4_bits_instrSize;
        output io_enq_req_4_bits_dirtyFs;
        output io_enq_req_4_bits_dirtyVs;
        output io_enq_req_4_bits_traceBlockInPipe_itype;
        output io_enq_req_4_bits_traceBlockInPipe_iretire;
        output io_enq_req_4_bits_traceBlockInPipe_ilastsize;
        output io_enq_req_4_bits_eliminatedMove;
        output io_enq_req_4_bits_snapshot;
        output io_enq_req_4_bits_lqIdx_value;
        output io_enq_req_4_bits_sqIdx_value;
        output io_enq_req_4_bits_singleStep;
        output io_enq_req_4_bits_debug_sim_trig;
        output io_enq_req_5_valid;
        output io_enq_req_5_bits_instr;
        output io_enq_req_5_bits_pc;
        output io_enq_req_5_bits_exceptionVec_0;
        output io_enq_req_5_bits_exceptionVec_1;
        output io_enq_req_5_bits_exceptionVec_2;
        output io_enq_req_5_bits_exceptionVec_3;
        output io_enq_req_5_bits_exceptionVec_12;
        output io_enq_req_5_bits_exceptionVec_20;
        output io_enq_req_5_bits_exceptionVec_22;
        output io_enq_req_5_bits_isFetchMalAddr;
        output io_enq_req_5_bits_hasException;
        output io_enq_req_5_bits_trigger;
        output io_enq_req_5_bits_preDecodeInfo_isRVC;
        output io_enq_req_5_bits_crossPageIPFFix;
        output io_enq_req_5_bits_ftqPtr_flag;
        output io_enq_req_5_bits_ftqPtr_value;
        output io_enq_req_5_bits_ftqOffset;
        output io_enq_req_5_bits_ldest;
        output io_enq_req_5_bits_fuType;
        output io_enq_req_5_bits_fuOpType;
        output io_enq_req_5_bits_rfWen;
        output io_enq_req_5_bits_fpWen;
        output io_enq_req_5_bits_vecWen;
        output io_enq_req_5_bits_v0Wen;
        output io_enq_req_5_bits_vlWen;
        output io_enq_req_5_bits_isXSTrap;
        output io_enq_req_5_bits_waitForward;
        output io_enq_req_5_bits_blockBackward;
        output io_enq_req_5_bits_flushPipe;
        output io_enq_req_5_bits_vpu_vill;
        output io_enq_req_5_bits_vpu_vma;
        output io_enq_req_5_bits_vpu_vta;
        output io_enq_req_5_bits_vpu_vsew;
        output io_enq_req_5_bits_vpu_vlmul;
        output io_enq_req_5_bits_vpu_specVill;
        output io_enq_req_5_bits_vpu_specVma;
        output io_enq_req_5_bits_vpu_specVta;
        output io_enq_req_5_bits_vpu_specVsew;
        output io_enq_req_5_bits_vpu_specVlmul;
        output io_enq_req_5_bits_vlsInstr;
        output io_enq_req_5_bits_wfflags;
        output io_enq_req_5_bits_isMove;
        output io_enq_req_5_bits_isVset;
        output io_enq_req_5_bits_firstUop;
        output io_enq_req_5_bits_lastUop;
        output io_enq_req_5_bits_numWB;
        output io_enq_req_5_bits_commitType;
        output io_enq_req_5_bits_pdest;
        output io_enq_req_5_bits_robIdx_flag;
        output io_enq_req_5_bits_robIdx_value;
        output io_enq_req_5_bits_instrSize;
        output io_enq_req_5_bits_dirtyFs;
        output io_enq_req_5_bits_dirtyVs;
        output io_enq_req_5_bits_traceBlockInPipe_itype;
        output io_enq_req_5_bits_traceBlockInPipe_iretire;
        output io_enq_req_5_bits_traceBlockInPipe_ilastsize;
        output io_enq_req_5_bits_eliminatedMove;
        output io_enq_req_5_bits_snapshot;
        output io_enq_req_5_bits_lqIdx_value;
        output io_enq_req_5_bits_sqIdx_value;
        output io_enq_req_5_bits_singleStep;
        output io_enq_req_5_bits_debug_sim_trig;

    endclocking:drv_cb

    clocking mon_cb @(posedge clk);
        `ifdef INTERFACE_ADD_DELAY
            default input #`DEF_SETUP_TIME output #`DEF_HOLD_TIME;
        `endif
        input  clock;
        input  reset;
        input  io_hartId;
        input  io_enq_req_0_valid;
        input  io_enq_req_0_bits_instr;
        input  io_enq_req_0_bits_pc;
        input  io_enq_req_0_bits_exceptionVec_0;
        input  io_enq_req_0_bits_exceptionVec_1;
        input  io_enq_req_0_bits_exceptionVec_2;
        input  io_enq_req_0_bits_exceptionVec_3;
        input  io_enq_req_0_bits_exceptionVec_12;
        input  io_enq_req_0_bits_exceptionVec_20;
        input  io_enq_req_0_bits_exceptionVec_22;
        input  io_enq_req_0_bits_isFetchMalAddr;
        input  io_enq_req_0_bits_hasException;
        input  io_enq_req_0_bits_trigger;
        input  io_enq_req_0_bits_preDecodeInfo_isRVC;
        input  io_enq_req_0_bits_crossPageIPFFix;
        input  io_enq_req_0_bits_ftqPtr_flag;
        input  io_enq_req_0_bits_ftqPtr_value;
        input  io_enq_req_0_bits_ftqOffset;
        input  io_enq_req_0_bits_ldest;
        input  io_enq_req_0_bits_fuType;
        input  io_enq_req_0_bits_fuOpType;
        input  io_enq_req_0_bits_rfWen;
        input  io_enq_req_0_bits_fpWen;
        input  io_enq_req_0_bits_vecWen;
        input  io_enq_req_0_bits_v0Wen;
        input  io_enq_req_0_bits_vlWen;
        input  io_enq_req_0_bits_isXSTrap;
        input  io_enq_req_0_bits_waitForward;
        input  io_enq_req_0_bits_blockBackward;
        input  io_enq_req_0_bits_flushPipe;
        input  io_enq_req_0_bits_vpu_vill;
        input  io_enq_req_0_bits_vpu_vma;
        input  io_enq_req_0_bits_vpu_vta;
        input  io_enq_req_0_bits_vpu_vsew;
        input  io_enq_req_0_bits_vpu_vlmul;
        input  io_enq_req_0_bits_vpu_specVill;
        input  io_enq_req_0_bits_vpu_specVma;
        input  io_enq_req_0_bits_vpu_specVta;
        input  io_enq_req_0_bits_vpu_specVsew;
        input  io_enq_req_0_bits_vpu_specVlmul;
        input  io_enq_req_0_bits_vlsInstr;
        input  io_enq_req_0_bits_wfflags;
        input  io_enq_req_0_bits_isMove;
        input  io_enq_req_0_bits_isVset;
        input  io_enq_req_0_bits_firstUop;
        input  io_enq_req_0_bits_lastUop;
        input  io_enq_req_0_bits_numWB;
        input  io_enq_req_0_bits_commitType;
        input  io_enq_req_0_bits_pdest;
        input  io_enq_req_0_bits_robIdx_flag;
        input  io_enq_req_0_bits_robIdx_value;
        input  io_enq_req_0_bits_instrSize;
        input  io_enq_req_0_bits_dirtyFs;
        input  io_enq_req_0_bits_dirtyVs;
        input  io_enq_req_0_bits_traceBlockInPipe_itype;
        input  io_enq_req_0_bits_traceBlockInPipe_iretire;
        input  io_enq_req_0_bits_traceBlockInPipe_ilastsize;
        input  io_enq_req_0_bits_eliminatedMove;
        input  io_enq_req_0_bits_snapshot;
        input  io_enq_req_0_bits_lqIdx_value;
        input  io_enq_req_0_bits_sqIdx_value;
        input  io_enq_req_0_bits_singleStep;
        input  io_enq_req_0_bits_debug_sim_trig;
        input  io_enq_req_1_valid;
        input  io_enq_req_1_bits_instr;
        input  io_enq_req_1_bits_pc;
        input  io_enq_req_1_bits_exceptionVec_0;
        input  io_enq_req_1_bits_exceptionVec_1;
        input  io_enq_req_1_bits_exceptionVec_2;
        input  io_enq_req_1_bits_exceptionVec_3;
        input  io_enq_req_1_bits_exceptionVec_12;
        input  io_enq_req_1_bits_exceptionVec_20;
        input  io_enq_req_1_bits_exceptionVec_22;
        input  io_enq_req_1_bits_isFetchMalAddr;
        input  io_enq_req_1_bits_hasException;
        input  io_enq_req_1_bits_trigger;
        input  io_enq_req_1_bits_preDecodeInfo_isRVC;
        input  io_enq_req_1_bits_crossPageIPFFix;
        input  io_enq_req_1_bits_ftqPtr_flag;
        input  io_enq_req_1_bits_ftqPtr_value;
        input  io_enq_req_1_bits_ftqOffset;
        input  io_enq_req_1_bits_ldest;
        input  io_enq_req_1_bits_fuType;
        input  io_enq_req_1_bits_fuOpType;
        input  io_enq_req_1_bits_rfWen;
        input  io_enq_req_1_bits_fpWen;
        input  io_enq_req_1_bits_vecWen;
        input  io_enq_req_1_bits_v0Wen;
        input  io_enq_req_1_bits_vlWen;
        input  io_enq_req_1_bits_isXSTrap;
        input  io_enq_req_1_bits_waitForward;
        input  io_enq_req_1_bits_blockBackward;
        input  io_enq_req_1_bits_flushPipe;
        input  io_enq_req_1_bits_vpu_vill;
        input  io_enq_req_1_bits_vpu_vma;
        input  io_enq_req_1_bits_vpu_vta;
        input  io_enq_req_1_bits_vpu_vsew;
        input  io_enq_req_1_bits_vpu_vlmul;
        input  io_enq_req_1_bits_vpu_specVill;
        input  io_enq_req_1_bits_vpu_specVma;
        input  io_enq_req_1_bits_vpu_specVta;
        input  io_enq_req_1_bits_vpu_specVsew;
        input  io_enq_req_1_bits_vpu_specVlmul;
        input  io_enq_req_1_bits_vlsInstr;
        input  io_enq_req_1_bits_wfflags;
        input  io_enq_req_1_bits_isMove;
        input  io_enq_req_1_bits_isVset;
        input  io_enq_req_1_bits_firstUop;
        input  io_enq_req_1_bits_lastUop;
        input  io_enq_req_1_bits_numWB;
        input  io_enq_req_1_bits_commitType;
        input  io_enq_req_1_bits_pdest;
        input  io_enq_req_1_bits_robIdx_flag;
        input  io_enq_req_1_bits_robIdx_value;
        input  io_enq_req_1_bits_instrSize;
        input  io_enq_req_1_bits_dirtyFs;
        input  io_enq_req_1_bits_dirtyVs;
        input  io_enq_req_1_bits_traceBlockInPipe_itype;
        input  io_enq_req_1_bits_traceBlockInPipe_iretire;
        input  io_enq_req_1_bits_traceBlockInPipe_ilastsize;
        input  io_enq_req_1_bits_eliminatedMove;
        input  io_enq_req_1_bits_snapshot;
        input  io_enq_req_1_bits_lqIdx_value;
        input  io_enq_req_1_bits_sqIdx_value;
        input  io_enq_req_1_bits_singleStep;
        input  io_enq_req_1_bits_debug_sim_trig;
        input  io_enq_req_2_valid;
        input  io_enq_req_2_bits_instr;
        input  io_enq_req_2_bits_pc;
        input  io_enq_req_2_bits_exceptionVec_0;
        input  io_enq_req_2_bits_exceptionVec_1;
        input  io_enq_req_2_bits_exceptionVec_2;
        input  io_enq_req_2_bits_exceptionVec_3;
        input  io_enq_req_2_bits_exceptionVec_12;
        input  io_enq_req_2_bits_exceptionVec_20;
        input  io_enq_req_2_bits_exceptionVec_22;
        input  io_enq_req_2_bits_isFetchMalAddr;
        input  io_enq_req_2_bits_hasException;
        input  io_enq_req_2_bits_trigger;
        input  io_enq_req_2_bits_preDecodeInfo_isRVC;
        input  io_enq_req_2_bits_crossPageIPFFix;
        input  io_enq_req_2_bits_ftqPtr_flag;
        input  io_enq_req_2_bits_ftqPtr_value;
        input  io_enq_req_2_bits_ftqOffset;
        input  io_enq_req_2_bits_ldest;
        input  io_enq_req_2_bits_fuType;
        input  io_enq_req_2_bits_fuOpType;
        input  io_enq_req_2_bits_rfWen;
        input  io_enq_req_2_bits_fpWen;
        input  io_enq_req_2_bits_vecWen;
        input  io_enq_req_2_bits_v0Wen;
        input  io_enq_req_2_bits_vlWen;
        input  io_enq_req_2_bits_isXSTrap;
        input  io_enq_req_2_bits_waitForward;
        input  io_enq_req_2_bits_blockBackward;
        input  io_enq_req_2_bits_flushPipe;
        input  io_enq_req_2_bits_vpu_vill;
        input  io_enq_req_2_bits_vpu_vma;
        input  io_enq_req_2_bits_vpu_vta;
        input  io_enq_req_2_bits_vpu_vsew;
        input  io_enq_req_2_bits_vpu_vlmul;
        input  io_enq_req_2_bits_vpu_specVill;
        input  io_enq_req_2_bits_vpu_specVma;
        input  io_enq_req_2_bits_vpu_specVta;
        input  io_enq_req_2_bits_vpu_specVsew;
        input  io_enq_req_2_bits_vpu_specVlmul;
        input  io_enq_req_2_bits_vlsInstr;
        input  io_enq_req_2_bits_wfflags;
        input  io_enq_req_2_bits_isMove;
        input  io_enq_req_2_bits_isVset;
        input  io_enq_req_2_bits_firstUop;
        input  io_enq_req_2_bits_lastUop;
        input  io_enq_req_2_bits_numWB;
        input  io_enq_req_2_bits_commitType;
        input  io_enq_req_2_bits_pdest;
        input  io_enq_req_2_bits_robIdx_flag;
        input  io_enq_req_2_bits_robIdx_value;
        input  io_enq_req_2_bits_instrSize;
        input  io_enq_req_2_bits_dirtyFs;
        input  io_enq_req_2_bits_dirtyVs;
        input  io_enq_req_2_bits_traceBlockInPipe_itype;
        input  io_enq_req_2_bits_traceBlockInPipe_iretire;
        input  io_enq_req_2_bits_traceBlockInPipe_ilastsize;
        input  io_enq_req_2_bits_eliminatedMove;
        input  io_enq_req_2_bits_snapshot;
        input  io_enq_req_2_bits_lqIdx_value;
        input  io_enq_req_2_bits_sqIdx_value;
        input  io_enq_req_2_bits_singleStep;
        input  io_enq_req_2_bits_debug_sim_trig;
        input  io_enq_req_3_valid;
        input  io_enq_req_3_bits_instr;
        input  io_enq_req_3_bits_pc;
        input  io_enq_req_3_bits_exceptionVec_0;
        input  io_enq_req_3_bits_exceptionVec_1;
        input  io_enq_req_3_bits_exceptionVec_2;
        input  io_enq_req_3_bits_exceptionVec_3;
        input  io_enq_req_3_bits_exceptionVec_12;
        input  io_enq_req_3_bits_exceptionVec_20;
        input  io_enq_req_3_bits_exceptionVec_22;
        input  io_enq_req_3_bits_isFetchMalAddr;
        input  io_enq_req_3_bits_hasException;
        input  io_enq_req_3_bits_trigger;
        input  io_enq_req_3_bits_preDecodeInfo_isRVC;
        input  io_enq_req_3_bits_crossPageIPFFix;
        input  io_enq_req_3_bits_ftqPtr_flag;
        input  io_enq_req_3_bits_ftqPtr_value;
        input  io_enq_req_3_bits_ftqOffset;
        input  io_enq_req_3_bits_ldest;
        input  io_enq_req_3_bits_fuType;
        input  io_enq_req_3_bits_fuOpType;
        input  io_enq_req_3_bits_rfWen;
        input  io_enq_req_3_bits_fpWen;
        input  io_enq_req_3_bits_vecWen;
        input  io_enq_req_3_bits_v0Wen;
        input  io_enq_req_3_bits_vlWen;
        input  io_enq_req_3_bits_isXSTrap;
        input  io_enq_req_3_bits_waitForward;
        input  io_enq_req_3_bits_blockBackward;
        input  io_enq_req_3_bits_flushPipe;
        input  io_enq_req_3_bits_vpu_vill;
        input  io_enq_req_3_bits_vpu_vma;
        input  io_enq_req_3_bits_vpu_vta;
        input  io_enq_req_3_bits_vpu_vsew;
        input  io_enq_req_3_bits_vpu_vlmul;
        input  io_enq_req_3_bits_vpu_specVill;
        input  io_enq_req_3_bits_vpu_specVma;
        input  io_enq_req_3_bits_vpu_specVta;
        input  io_enq_req_3_bits_vpu_specVsew;
        input  io_enq_req_3_bits_vpu_specVlmul;
        input  io_enq_req_3_bits_vlsInstr;
        input  io_enq_req_3_bits_wfflags;
        input  io_enq_req_3_bits_isMove;
        input  io_enq_req_3_bits_isVset;
        input  io_enq_req_3_bits_firstUop;
        input  io_enq_req_3_bits_lastUop;
        input  io_enq_req_3_bits_numWB;
        input  io_enq_req_3_bits_commitType;
        input  io_enq_req_3_bits_pdest;
        input  io_enq_req_3_bits_robIdx_flag;
        input  io_enq_req_3_bits_robIdx_value;
        input  io_enq_req_3_bits_instrSize;
        input  io_enq_req_3_bits_dirtyFs;
        input  io_enq_req_3_bits_dirtyVs;
        input  io_enq_req_3_bits_traceBlockInPipe_itype;
        input  io_enq_req_3_bits_traceBlockInPipe_iretire;
        input  io_enq_req_3_bits_traceBlockInPipe_ilastsize;
        input  io_enq_req_3_bits_eliminatedMove;
        input  io_enq_req_3_bits_snapshot;
        input  io_enq_req_3_bits_lqIdx_value;
        input  io_enq_req_3_bits_sqIdx_value;
        input  io_enq_req_3_bits_singleStep;
        input  io_enq_req_3_bits_debug_sim_trig;
        input  io_enq_req_4_valid;
        input  io_enq_req_4_bits_instr;
        input  io_enq_req_4_bits_pc;
        input  io_enq_req_4_bits_exceptionVec_0;
        input  io_enq_req_4_bits_exceptionVec_1;
        input  io_enq_req_4_bits_exceptionVec_2;
        input  io_enq_req_4_bits_exceptionVec_3;
        input  io_enq_req_4_bits_exceptionVec_12;
        input  io_enq_req_4_bits_exceptionVec_20;
        input  io_enq_req_4_bits_exceptionVec_22;
        input  io_enq_req_4_bits_isFetchMalAddr;
        input  io_enq_req_4_bits_hasException;
        input  io_enq_req_4_bits_trigger;
        input  io_enq_req_4_bits_preDecodeInfo_isRVC;
        input  io_enq_req_4_bits_crossPageIPFFix;
        input  io_enq_req_4_bits_ftqPtr_flag;
        input  io_enq_req_4_bits_ftqPtr_value;
        input  io_enq_req_4_bits_ftqOffset;
        input  io_enq_req_4_bits_ldest;
        input  io_enq_req_4_bits_fuType;
        input  io_enq_req_4_bits_fuOpType;
        input  io_enq_req_4_bits_rfWen;
        input  io_enq_req_4_bits_fpWen;
        input  io_enq_req_4_bits_vecWen;
        input  io_enq_req_4_bits_v0Wen;
        input  io_enq_req_4_bits_vlWen;
        input  io_enq_req_4_bits_isXSTrap;
        input  io_enq_req_4_bits_waitForward;
        input  io_enq_req_4_bits_blockBackward;
        input  io_enq_req_4_bits_flushPipe;
        input  io_enq_req_4_bits_vpu_vill;
        input  io_enq_req_4_bits_vpu_vma;
        input  io_enq_req_4_bits_vpu_vta;
        input  io_enq_req_4_bits_vpu_vsew;
        input  io_enq_req_4_bits_vpu_vlmul;
        input  io_enq_req_4_bits_vpu_specVill;
        input  io_enq_req_4_bits_vpu_specVma;
        input  io_enq_req_4_bits_vpu_specVta;
        input  io_enq_req_4_bits_vpu_specVsew;
        input  io_enq_req_4_bits_vpu_specVlmul;
        input  io_enq_req_4_bits_vlsInstr;
        input  io_enq_req_4_bits_wfflags;
        input  io_enq_req_4_bits_isMove;
        input  io_enq_req_4_bits_isVset;
        input  io_enq_req_4_bits_firstUop;
        input  io_enq_req_4_bits_lastUop;
        input  io_enq_req_4_bits_numWB;
        input  io_enq_req_4_bits_commitType;
        input  io_enq_req_4_bits_pdest;
        input  io_enq_req_4_bits_robIdx_flag;
        input  io_enq_req_4_bits_robIdx_value;
        input  io_enq_req_4_bits_instrSize;
        input  io_enq_req_4_bits_dirtyFs;
        input  io_enq_req_4_bits_dirtyVs;
        input  io_enq_req_4_bits_traceBlockInPipe_itype;
        input  io_enq_req_4_bits_traceBlockInPipe_iretire;
        input  io_enq_req_4_bits_traceBlockInPipe_ilastsize;
        input  io_enq_req_4_bits_eliminatedMove;
        input  io_enq_req_4_bits_snapshot;
        input  io_enq_req_4_bits_lqIdx_value;
        input  io_enq_req_4_bits_sqIdx_value;
        input  io_enq_req_4_bits_singleStep;
        input  io_enq_req_4_bits_debug_sim_trig;
        input  io_enq_req_5_valid;
        input  io_enq_req_5_bits_instr;
        input  io_enq_req_5_bits_pc;
        input  io_enq_req_5_bits_exceptionVec_0;
        input  io_enq_req_5_bits_exceptionVec_1;
        input  io_enq_req_5_bits_exceptionVec_2;
        input  io_enq_req_5_bits_exceptionVec_3;
        input  io_enq_req_5_bits_exceptionVec_12;
        input  io_enq_req_5_bits_exceptionVec_20;
        input  io_enq_req_5_bits_exceptionVec_22;
        input  io_enq_req_5_bits_isFetchMalAddr;
        input  io_enq_req_5_bits_hasException;
        input  io_enq_req_5_bits_trigger;
        input  io_enq_req_5_bits_preDecodeInfo_isRVC;
        input  io_enq_req_5_bits_crossPageIPFFix;
        input  io_enq_req_5_bits_ftqPtr_flag;
        input  io_enq_req_5_bits_ftqPtr_value;
        input  io_enq_req_5_bits_ftqOffset;
        input  io_enq_req_5_bits_ldest;
        input  io_enq_req_5_bits_fuType;
        input  io_enq_req_5_bits_fuOpType;
        input  io_enq_req_5_bits_rfWen;
        input  io_enq_req_5_bits_fpWen;
        input  io_enq_req_5_bits_vecWen;
        input  io_enq_req_5_bits_v0Wen;
        input  io_enq_req_5_bits_vlWen;
        input  io_enq_req_5_bits_isXSTrap;
        input  io_enq_req_5_bits_waitForward;
        input  io_enq_req_5_bits_blockBackward;
        input  io_enq_req_5_bits_flushPipe;
        input  io_enq_req_5_bits_vpu_vill;
        input  io_enq_req_5_bits_vpu_vma;
        input  io_enq_req_5_bits_vpu_vta;
        input  io_enq_req_5_bits_vpu_vsew;
        input  io_enq_req_5_bits_vpu_vlmul;
        input  io_enq_req_5_bits_vpu_specVill;
        input  io_enq_req_5_bits_vpu_specVma;
        input  io_enq_req_5_bits_vpu_specVta;
        input  io_enq_req_5_bits_vpu_specVsew;
        input  io_enq_req_5_bits_vpu_specVlmul;
        input  io_enq_req_5_bits_vlsInstr;
        input  io_enq_req_5_bits_wfflags;
        input  io_enq_req_5_bits_isMove;
        input  io_enq_req_5_bits_isVset;
        input  io_enq_req_5_bits_firstUop;
        input  io_enq_req_5_bits_lastUop;
        input  io_enq_req_5_bits_numWB;
        input  io_enq_req_5_bits_commitType;
        input  io_enq_req_5_bits_pdest;
        input  io_enq_req_5_bits_robIdx_flag;
        input  io_enq_req_5_bits_robIdx_value;
        input  io_enq_req_5_bits_instrSize;
        input  io_enq_req_5_bits_dirtyFs;
        input  io_enq_req_5_bits_dirtyVs;
        input  io_enq_req_5_bits_traceBlockInPipe_itype;
        input  io_enq_req_5_bits_traceBlockInPipe_iretire;
        input  io_enq_req_5_bits_traceBlockInPipe_ilastsize;
        input  io_enq_req_5_bits_eliminatedMove;
        input  io_enq_req_5_bits_snapshot;
        input  io_enq_req_5_bits_lqIdx_value;
        input  io_enq_req_5_bits_sqIdx_value;
        input  io_enq_req_5_bits_singleStep;
        input  io_enq_req_5_bits_debug_sim_trig;

    endclocking:mon_cb

    modport drv_mp (clocking drv_cb);
    modport mon_mp (clocking mon_cb);

endinterface:rename_in_agent_interface

`endif


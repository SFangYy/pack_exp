`ifndef SV_MAIN__SV
`define SV_MAIN__SV

module sv_main;
    // Instantiate top_tb module
    top_tb u_top_tb();
endmodule

`endif
//==============================================================================
// Transaction: CSR_in_agent_xaction
//==============================================================================

import uvm_pkg::*;
import uvmc_pkg::*;
import utils_pkg::*;
import CSR_in_agent_pkg::*;

`include "uvm_macros.svh"

class CSR_in_agent_xaction_xmonitor extends uvm_monitor;
    `uvm_component_utils(CSR_in_agent_xaction_xmonitor)

    uvm_tlm_b_initiator_socket #() out;
    byte unsigned m_transport_data[];
    uvm_tlm_gp m_transport_msg;
    uvm_tlm_time m_delay;
    uvm_active_passive_enum m_exist_xmonitor;
    CSR_in_agent_xaction m_tr;

    function new(string name, uvm_component parent=null);
        super.new(name,parent);
        if(!uvm_config_db#(uvm_active_passive_enum)::get(this,"","CSR_in_agent_xaction_exist_xmonitor",m_exist_xmonitor))
            m_exist_xmonitor = UVM_ACTIVE; // Default to active if not configured
        out = new("out",this);
        m_transport_msg = new;
        m_transport_data = new[58];
        m_delay = new("delay", TIME_UNIT);
    endfunction

    virtual task run_phase(uvm_phase phase);
        // Monitor typically doesn't need an active run_phase unless actively sampling
        // Remove forever loop to prevent simulation hang
        // Users can override this method if active monitoring is needed 
    endtask

    virtual task sequence_send(CSR_in_agent_xaction tr);
        // Optimized serialization using pre-allocated array and utility functions
        
        `PICKER_PACK_BYTE(tr.io_csr_intrBitSet, 0);
        
        
        `PICKER_PACK_BYTE(tr.io_csr_wfiEvent, 1);
        
        
        `PICKER_PACK_BYTE(tr.io_csr_criticalErrorState, 2);
        
        
        `PICKER_PACK_BYTE(tr.io_snpt_snptDeq, 3);
        
        
        `PICKER_PACK_BYTE(tr.io_snpt_useSnpt, 4);
        
        
        `PICKER_PACK_BYTE(tr.io_snpt_snptSelect, 5);
        
        
        `PICKER_PACK_BYTE(tr.io_snpt_flushVec_0, 6);
        
        
        `PICKER_PACK_BYTE(tr.io_snpt_flushVec_1, 7);
        
        
        `PICKER_PACK_BYTE(tr.io_snpt_flushVec_2, 8);
        
        
        `PICKER_PACK_BYTE(tr.io_snpt_flushVec_3, 9);
        
        
        `PICKER_PACK_BYTE(tr.io_wfi_safeFromMem, 10);
        
        
        `PICKER_PACK_BYTE(tr.io_wfi_safeFromFrontend, 11);
        
        
        `PICKER_PACK_BYTE(tr.io_wfi_enable, 12);
        
        
        `PICKER_PACK_BYTE(tr.io_fromVecExcpMod_busy, 13);
        
        
        `PICKER_PACK_STREAM(tr.io_readGPAMemData_gpaddr, 14, 56);
        
        
        `PICKER_PACK_BYTE(tr.io_readGPAMemData_isForVSnonLeafPTE, 21);
        
        
        `PICKER_PACK_BYTE(tr.io_vstartIsZero, 22);
        
        
        `PICKER_PACK_BYTE(tr.io_debugEnqLsq_canAccept, 23);
        
        
        `PICKER_PACK_BYTE(tr.io_debugEnqLsq_needAlloc_0, 24);
        
        
        `PICKER_PACK_BYTE(tr.io_debugEnqLsq_needAlloc_1, 25);
        
        
        `PICKER_PACK_BYTE(tr.io_debugEnqLsq_needAlloc_2, 26);
        
        
        `PICKER_PACK_BYTE(tr.io_debugEnqLsq_needAlloc_3, 27);
        
        
        `PICKER_PACK_BYTE(tr.io_debugEnqLsq_needAlloc_4, 28);
        
        
        `PICKER_PACK_BYTE(tr.io_debugEnqLsq_needAlloc_5, 29);
        
        
        `PICKER_PACK_BYTE(tr.io_debugEnqLsq_req_0_valid, 30);
        
        
        `PICKER_PACK_BYTE(tr.io_debugEnqLsq_req_0_bits_robIdx_value, 31);
        
        
        `PICKER_PACK_BYTE(tr.io_debugEnqLsq_req_0_bits_lqIdx_value, 32);
        
        
        `PICKER_PACK_BYTE(tr.io_debugEnqLsq_req_1_valid, 33);
        
        
        `PICKER_PACK_BYTE(tr.io_debugEnqLsq_req_1_bits_robIdx_value, 34);
        
        
        `PICKER_PACK_BYTE(tr.io_debugEnqLsq_req_1_bits_lqIdx_value, 35);
        
        
        `PICKER_PACK_BYTE(tr.io_debugEnqLsq_req_2_valid, 36);
        
        
        `PICKER_PACK_BYTE(tr.io_debugEnqLsq_req_2_bits_robIdx_value, 37);
        
        
        `PICKER_PACK_BYTE(tr.io_debugEnqLsq_req_2_bits_lqIdx_value, 38);
        
        
        `PICKER_PACK_BYTE(tr.io_debugEnqLsq_req_3_valid, 39);
        
        
        `PICKER_PACK_BYTE(tr.io_debugEnqLsq_req_3_bits_robIdx_value, 40);
        
        
        `PICKER_PACK_BYTE(tr.io_debugEnqLsq_req_3_bits_lqIdx_value, 41);
        
        
        `PICKER_PACK_BYTE(tr.io_debugEnqLsq_req_4_valid, 42);
        
        
        `PICKER_PACK_BYTE(tr.io_debugEnqLsq_req_4_bits_robIdx_value, 43);
        
        
        `PICKER_PACK_BYTE(tr.io_debugEnqLsq_req_4_bits_lqIdx_value, 44);
        
        
        `PICKER_PACK_BYTE(tr.io_debugEnqLsq_req_5_valid, 45);
        
        
        `PICKER_PACK_BYTE(tr.io_debugEnqLsq_req_5_bits_robIdx_value, 46);
        
        
        `PICKER_PACK_BYTE(tr.io_debugEnqLsq_req_5_bits_lqIdx_value, 47);
        
        
        `PICKER_PACK_BYTE(tr.io_debugInstrAddrTransType_bare, 48);
        
        
        `PICKER_PACK_BYTE(tr.io_debugInstrAddrTransType_sv39, 49);
        
        
        `PICKER_PACK_BYTE(tr.io_debugInstrAddrTransType_sv39x4, 50);
        
        
        `PICKER_PACK_BYTE(tr.io_debugInstrAddrTransType_sv48, 51);
        
        
        `PICKER_PACK_BYTE(tr.io_debugInstrAddrTransType_sv48x4, 52);
        
        
        `PICKER_PACK_BYTE(tr.io_storeDebugInfo_0_robidx_value, 53);
        
        
        `PICKER_PACK_BYTE(tr.io_storeDebugInfo_1_robidx_value, 54);
        
        
        `PICKER_PACK_BYTE(tr.compare, 55);
        
        
        `PICKER_PACK_BYTE(tr.CSR_in_agent_xaction, 56);
        
        
        `PICKER_PACK_BYTE(tr.super_result, 57);
        
        m_transport_msg.set_data_length(58);
        m_transport_msg.set_data(m_transport_data);
        m_delay.set_abstime(0, TRANSPORT_DELAY);
        out.b_transport(m_transport_msg, m_delay);
    endtask

endclass
    
class CSR_in_agent_xaction_xdriver extends uvm_driver;
    `uvm_component_utils(CSR_in_agent_xaction_xdriver)

    uvm_tlm_gp m_transport_msg;
    uvm_tlm_time m_delay;
    byte unsigned m_transport_data[];
    uvm_tlm_b_target_socket #(CSR_in_agent_xaction_xdriver) in;
    CSR_in_agent_xaction m_tr;

    function new(string name, uvm_component parent=null);
        super.new(name,parent);
        in = new("in",this);
        m_transport_msg = new("transport_msg");
        m_tr = new("tr");
        m_delay = new("delay", TIME_UNIT);
    endfunction

    virtual task b_transport(uvm_tlm_gp t, uvm_tlm_time delay);
        t.get_data(m_transport_data);
        // Deserialize using optimized utility functions
        m_tr.io_csr_intrBitSet = m_transport_data[0];
        m_tr.io_csr_wfiEvent = m_transport_data[1];
        m_tr.io_csr_criticalErrorState = m_transport_data[2];
        m_tr.io_snpt_snptDeq = m_transport_data[3];
        m_tr.io_snpt_useSnpt = m_transport_data[4];
        m_tr.io_snpt_snptSelect = m_transport_data[5];
        m_tr.io_snpt_flushVec_0 = m_transport_data[6];
        m_tr.io_snpt_flushVec_1 = m_transport_data[7];
        m_tr.io_snpt_flushVec_2 = m_transport_data[8];
        m_tr.io_snpt_flushVec_3 = m_transport_data[9];
        m_tr.io_wfi_safeFromMem = m_transport_data[10];
        m_tr.io_wfi_safeFromFrontend = m_transport_data[11];
        m_tr.io_wfi_enable = m_transport_data[12];
        m_tr.io_fromVecExcpMod_busy = m_transport_data[13];
        
        `PICKER_UNPACK_STREAM(m_tr.io_readGPAMemData_gpaddr, 14, 56);
        
        m_tr.io_readGPAMemData_isForVSnonLeafPTE = m_transport_data[21];
        m_tr.io_vstartIsZero = m_transport_data[22];
        m_tr.io_debugEnqLsq_canAccept = m_transport_data[23];
        m_tr.io_debugEnqLsq_needAlloc_0 = m_transport_data[24];
        m_tr.io_debugEnqLsq_needAlloc_1 = m_transport_data[25];
        m_tr.io_debugEnqLsq_needAlloc_2 = m_transport_data[26];
        m_tr.io_debugEnqLsq_needAlloc_3 = m_transport_data[27];
        m_tr.io_debugEnqLsq_needAlloc_4 = m_transport_data[28];
        m_tr.io_debugEnqLsq_needAlloc_5 = m_transport_data[29];
        m_tr.io_debugEnqLsq_req_0_valid = m_transport_data[30];
        m_tr.io_debugEnqLsq_req_0_bits_robIdx_value = m_transport_data[31];
        m_tr.io_debugEnqLsq_req_0_bits_lqIdx_value = m_transport_data[32];
        m_tr.io_debugEnqLsq_req_1_valid = m_transport_data[33];
        m_tr.io_debugEnqLsq_req_1_bits_robIdx_value = m_transport_data[34];
        m_tr.io_debugEnqLsq_req_1_bits_lqIdx_value = m_transport_data[35];
        m_tr.io_debugEnqLsq_req_2_valid = m_transport_data[36];
        m_tr.io_debugEnqLsq_req_2_bits_robIdx_value = m_transport_data[37];
        m_tr.io_debugEnqLsq_req_2_bits_lqIdx_value = m_transport_data[38];
        m_tr.io_debugEnqLsq_req_3_valid = m_transport_data[39];
        m_tr.io_debugEnqLsq_req_3_bits_robIdx_value = m_transport_data[40];
        m_tr.io_debugEnqLsq_req_3_bits_lqIdx_value = m_transport_data[41];
        m_tr.io_debugEnqLsq_req_4_valid = m_transport_data[42];
        m_tr.io_debugEnqLsq_req_4_bits_robIdx_value = m_transport_data[43];
        m_tr.io_debugEnqLsq_req_4_bits_lqIdx_value = m_transport_data[44];
        m_tr.io_debugEnqLsq_req_5_valid = m_transport_data[45];
        m_tr.io_debugEnqLsq_req_5_bits_robIdx_value = m_transport_data[46];
        m_tr.io_debugEnqLsq_req_5_bits_lqIdx_value = m_transport_data[47];
        m_tr.io_debugInstrAddrTransType_bare = m_transport_data[48];
        m_tr.io_debugInstrAddrTransType_sv39 = m_transport_data[49];
        m_tr.io_debugInstrAddrTransType_sv39x4 = m_transport_data[50];
        m_tr.io_debugInstrAddrTransType_sv48 = m_transport_data[51];
        m_tr.io_debugInstrAddrTransType_sv48x4 = m_transport_data[52];
        m_tr.io_storeDebugInfo_0_robidx_value = m_transport_data[53];
        m_tr.io_storeDebugInfo_1_robidx_value = m_transport_data[54];
        m_tr.compare = m_transport_data[55];
        m_tr.CSR_in_agent_xaction = m_transport_data[56];
        m_tr.super_result = m_transport_data[57];
        delay.reset();
        sequence_receive(m_tr);
    endtask

    virtual task sequence_receive(CSR_in_agent_xaction tr);
    endtask
endclass

class CSR_in_agent_xaction_xagent_config extends uvm_object;
    // UVM standard configuration using is_active
    uvm_active_passive_enum is_active = UVM_ACTIVE;  // UVM_ACTIVE: monitor+driver, UVM_PASSIVE: monitor only
    string channel_name;    // TLM channel name for both monitor and driver

    `uvm_object_utils_begin(CSR_in_agent_xaction_xagent_config)
        `uvm_field_enum(uvm_active_passive_enum, is_active, UVM_DEFAULT)
        `uvm_field_string(channel_name, UVM_DEFAULT)
    `uvm_object_utils_end

    function new(string name = "CSR_in_agent_xaction_xagent_config");
        super.new(name);
        this.channel_name = "CSR_in_agent_xaction";
    endfunction
endclass

class CSR_in_agent_xaction_xagent extends uvm_agent;
    `uvm_component_utils(CSR_in_agent_xaction_xagent)

    CSR_in_agent_xaction_xagent_config cfg;
    CSR_in_agent_xaction_xmonitor CSR_in_agent_xaction_xmon;
    CSR_in_agent_xaction_xdriver CSR_in_agent_xaction_xdrv;

    function new(string name, uvm_component parent = null);
        super.new(name,parent);
        if (!uvm_config_db#(CSR_in_agent_xaction_xagent_config)::get(this, "", "CSR_in_agent_xaction_xagent_config", cfg))
            `uvm_fatal("CFGERR", "Could not get xagent_config")

        // Set is_active for monitor (always exists, just needs to know mode for potential internal logic)
        uvm_config_db#(uvm_active_passive_enum)::set(this, "*", "CSR_in_agent_xaction_exist_xmonitor", cfg.is_active);
    endfunction

    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        // Monitor always created (both ACTIVE and PASSIVE modes have monitors)
        CSR_in_agent_xaction_xmon = CSR_in_agent_xaction_xmonitor::type_id::create($sformatf("%s_sub", cfg.channel_name), this);

        // Driver only created in ACTIVE mode
        if(cfg.is_active == UVM_ACTIVE) begin
            CSR_in_agent_xaction_xdrv = CSR_in_agent_xaction_xdriver::type_id::create($sformatf("%s.pub", cfg.channel_name), this);
        end
    endfunction

    // Standard UVM connect_phase for TLM connections
    function void connect_phase(uvm_phase phase);
        super.connect_phase(phase);

        // Monitor TLM connection (always present)
        uvmc_tlm #()::connect(CSR_in_agent_xaction_xmon.out, $sformatf("%s.sub", cfg.channel_name));

        // Driver TLM connection (only in ACTIVE mode)
        if(cfg.is_active == UVM_ACTIVE) begin
            uvmc_tlm #()::connect(CSR_in_agent_xaction_xdrv.in, $sformatf("%s.pub", cfg.channel_name));
        end
    endfunction

endclass


//=========================================================
//File name    : Rob_output_agent_interface.sv
//Author       : nanyunhao
//Module name  : Rob_output_agent_interface
//Discribution : Rob_output_agent_interface : signal interface
//Date         : 2026-01-22
//=========================================================
`ifndef ROB_OUTPUT_AGENT_INTERFACE__SV
`define ROB_OUTPUT_AGENT_INTERFACE__SV

`ifndef DEF_SETUP_TIME
    `define DEF_SETUP_TIME 1
`endif
`ifndef DEF_HOLD_TIME
    `define DEF_HOLD_TIME 1
`endif

interface Rob_output_agent_interface  (input bit clk,input bit rst_n);

    logic         io_enq_canAccept     ;
    logic         io_enq_canAcceptForDispatch;
    logic         io_enq_isEmpty       ;
    logic         io_flushOut_valid    ;
    logic         io_flushOut_bits_isRVC;
    logic         io_flushOut_bits_robIdx_flag;
    logic [7:0]   io_flushOut_bits_robIdx_value;
    logic         io_flushOut_bits_ftqIdx_flag;
    logic [5:0]   io_flushOut_bits_ftqIdx_value;
    logic [3:0]   io_flushOut_bits_ftqOffset;
    logic         io_flushOut_bits_level;
    logic         io_exception_valid   ;
    logic [31:0]  io_exception_bits_instr;
    logic [2:0]   io_exception_bits_commitType;
    logic         io_exception_bits_exceptionVec_0;
    logic         io_exception_bits_exceptionVec_1;
    logic         io_exception_bits_exceptionVec_2;
    logic         io_exception_bits_exceptionVec_3;
    logic         io_exception_bits_exceptionVec_4;
    logic         io_exception_bits_exceptionVec_5;
    logic         io_exception_bits_exceptionVec_6;
    logic         io_exception_bits_exceptionVec_7;
    logic         io_exception_bits_exceptionVec_8;
    logic         io_exception_bits_exceptionVec_9;
    logic         io_exception_bits_exceptionVec_10;
    logic         io_exception_bits_exceptionVec_11;
    logic         io_exception_bits_exceptionVec_12;
    logic         io_exception_bits_exceptionVec_13;
    logic         io_exception_bits_exceptionVec_14;
    logic         io_exception_bits_exceptionVec_15;
    logic         io_exception_bits_exceptionVec_16;
    logic         io_exception_bits_exceptionVec_17;
    logic         io_exception_bits_exceptionVec_18;
    logic         io_exception_bits_exceptionVec_19;
    logic         io_exception_bits_exceptionVec_20;
    logic         io_exception_bits_exceptionVec_21;
    logic         io_exception_bits_exceptionVec_22;
    logic         io_exception_bits_exceptionVec_23;
    logic         io_exception_bits_isPcBkpt;
    logic         io_exception_bits_isFetchMalAddr;
    logic [63:0]  io_exception_bits_gpaddr;
    logic         io_exception_bits_singleStep;
    logic         io_exception_bits_crossPageIPFFix;
    logic         io_exception_bits_isInterrupt;
    logic         io_exception_bits_isHls;
    logic [3:0]   io_exception_bits_trigger;
    logic         io_exception_bits_isForVSnonLeafPTE;
    logic         io_commits_isCommit  ;
    logic         io_commits_commitValid_0;
    logic         io_commits_commitValid_1;
    logic         io_commits_commitValid_2;
    logic         io_commits_commitValid_3;
    logic         io_commits_commitValid_4;
    logic         io_commits_commitValid_5;
    logic         io_commits_commitValid_6;
    logic         io_commits_commitValid_7;
    logic         io_commits_isWalk    ;
    logic         io_commits_walkValid_0;
    logic         io_commits_walkValid_1;
    logic         io_commits_walkValid_2;
    logic         io_commits_walkValid_3;
    logic         io_commits_walkValid_4;
    logic         io_commits_walkValid_5;
    logic         io_commits_walkValid_6;
    logic         io_commits_walkValid_7;
    logic         io_commits_info_0_walk_v;
    logic         io_commits_info_0_commit_v;
    logic         io_commits_info_0_commit_w;
    logic [6:0]   io_commits_info_0_realDestSize;
    logic         io_commits_info_0_interrupt_safe;
    logic         io_commits_info_0_wflags;
    logic [4:0]   io_commits_info_0_fflags;
    logic         io_commits_info_0_vxsat;
    logic         io_commits_info_0_isRVC;
    logic         io_commits_info_0_isVset;
    logic         io_commits_info_0_isHls;
    logic         io_commits_info_0_isVls;
    logic         io_commits_info_0_vls;
    logic         io_commits_info_0_mmio;
    logic [2:0]   io_commits_info_0_commitType;
    logic         io_commits_info_0_ftqIdx_flag;
    logic [5:0]   io_commits_info_0_ftqIdx_value;
    logic [3:0]   io_commits_info_0_ftqOffset;
    logic [2:0]   io_commits_info_0_instrSize;
    logic         io_commits_info_0_fpWen;
    logic         io_commits_info_0_rfWen;
    logic         io_commits_info_0_needFlush;
    logic [3:0]   io_commits_info_0_traceBlockInPipe_itype;
    logic [3:0]   io_commits_info_0_traceBlockInPipe_iretire;
    logic         io_commits_info_0_traceBlockInPipe_ilastsize;
    logic [49:0]  io_commits_info_0_debug_pc;
    logic [31:0]  io_commits_info_0_debug_instr;
    logic [5:0]   io_commits_info_0_debug_ldest;
    logic [7:0]   io_commits_info_0_debug_pdest;
    logic [7:0]   io_commits_info_0_debug_otherPdest_0;
    logic [7:0]   io_commits_info_0_debug_otherPdest_1;
    logic [7:0]   io_commits_info_0_debug_otherPdest_2;
    logic [7:0]   io_commits_info_0_debug_otherPdest_3;
    logic [7:0]   io_commits_info_0_debug_otherPdest_4;
    logic [7:0]   io_commits_info_0_debug_otherPdest_5;
    logic [7:0]   io_commits_info_0_debug_otherPdest_6;
    logic [34:0]  io_commits_info_0_debug_fuType;
    logic         io_commits_info_0_dirtyFs;
    logic         io_commits_info_0_dirtyVs;
    logic         io_commits_info_1_walk_v;
    logic         io_commits_info_1_commit_v;
    logic         io_commits_info_1_commit_w;
    logic [6:0]   io_commits_info_1_realDestSize;
    logic         io_commits_info_1_interrupt_safe;
    logic         io_commits_info_1_wflags;
    logic [4:0]   io_commits_info_1_fflags;
    logic         io_commits_info_1_vxsat;
    logic         io_commits_info_1_isRVC;
    logic         io_commits_info_1_isVset;
    logic         io_commits_info_1_isHls;
    logic         io_commits_info_1_isVls;
    logic         io_commits_info_1_vls;
    logic         io_commits_info_1_mmio;
    logic [2:0]   io_commits_info_1_commitType;
    logic         io_commits_info_1_ftqIdx_flag;
    logic [5:0]   io_commits_info_1_ftqIdx_value;
    logic [3:0]   io_commits_info_1_ftqOffset;
    logic [2:0]   io_commits_info_1_instrSize;
    logic         io_commits_info_1_fpWen;
    logic         io_commits_info_1_rfWen;
    logic         io_commits_info_1_needFlush;
    logic [3:0]   io_commits_info_1_traceBlockInPipe_itype;
    logic [3:0]   io_commits_info_1_traceBlockInPipe_iretire;
    logic         io_commits_info_1_traceBlockInPipe_ilastsize;
    logic [49:0]  io_commits_info_1_debug_pc;
    logic [31:0]  io_commits_info_1_debug_instr;
    logic [5:0]   io_commits_info_1_debug_ldest;
    logic [7:0]   io_commits_info_1_debug_pdest;
    logic [7:0]   io_commits_info_1_debug_otherPdest_0;
    logic [7:0]   io_commits_info_1_debug_otherPdest_1;
    logic [7:0]   io_commits_info_1_debug_otherPdest_2;
    logic [7:0]   io_commits_info_1_debug_otherPdest_3;
    logic [7:0]   io_commits_info_1_debug_otherPdest_4;
    logic [7:0]   io_commits_info_1_debug_otherPdest_5;
    logic [7:0]   io_commits_info_1_debug_otherPdest_6;
    logic [34:0]  io_commits_info_1_debug_fuType;
    logic         io_commits_info_1_dirtyFs;
    logic         io_commits_info_1_dirtyVs;
    logic         io_commits_info_2_walk_v;
    logic         io_commits_info_2_commit_v;
    logic         io_commits_info_2_commit_w;
    logic [6:0]   io_commits_info_2_realDestSize;
    logic         io_commits_info_2_interrupt_safe;
    logic         io_commits_info_2_wflags;
    logic [4:0]   io_commits_info_2_fflags;
    logic         io_commits_info_2_vxsat;
    logic         io_commits_info_2_isRVC;
    logic         io_commits_info_2_isVset;
    logic         io_commits_info_2_isHls;
    logic         io_commits_info_2_isVls;
    logic         io_commits_info_2_vls;
    logic         io_commits_info_2_mmio;
    logic [2:0]   io_commits_info_2_commitType;
    logic         io_commits_info_2_ftqIdx_flag;
    logic [5:0]   io_commits_info_2_ftqIdx_value;
    logic [3:0]   io_commits_info_2_ftqOffset;
    logic [2:0]   io_commits_info_2_instrSize;
    logic         io_commits_info_2_fpWen;
    logic         io_commits_info_2_rfWen;
    logic         io_commits_info_2_needFlush;
    logic [3:0]   io_commits_info_2_traceBlockInPipe_itype;
    logic [3:0]   io_commits_info_2_traceBlockInPipe_iretire;
    logic         io_commits_info_2_traceBlockInPipe_ilastsize;
    logic [49:0]  io_commits_info_2_debug_pc;
    logic [31:0]  io_commits_info_2_debug_instr;
    logic [5:0]   io_commits_info_2_debug_ldest;
    logic [7:0]   io_commits_info_2_debug_pdest;
    logic [7:0]   io_commits_info_2_debug_otherPdest_0;
    logic [7:0]   io_commits_info_2_debug_otherPdest_1;
    logic [7:0]   io_commits_info_2_debug_otherPdest_2;
    logic [7:0]   io_commits_info_2_debug_otherPdest_3;
    logic [7:0]   io_commits_info_2_debug_otherPdest_4;
    logic [7:0]   io_commits_info_2_debug_otherPdest_5;
    logic [7:0]   io_commits_info_2_debug_otherPdest_6;
    logic [34:0]  io_commits_info_2_debug_fuType;
    logic         io_commits_info_2_dirtyFs;
    logic         io_commits_info_2_dirtyVs;
    logic         io_commits_info_3_walk_v;
    logic         io_commits_info_3_commit_v;
    logic         io_commits_info_3_commit_w;
    logic [6:0]   io_commits_info_3_realDestSize;
    logic         io_commits_info_3_interrupt_safe;
    logic         io_commits_info_3_wflags;
    logic [4:0]   io_commits_info_3_fflags;
    logic         io_commits_info_3_vxsat;
    logic         io_commits_info_3_isRVC;
    logic         io_commits_info_3_isVset;
    logic         io_commits_info_3_isHls;
    logic         io_commits_info_3_isVls;
    logic         io_commits_info_3_vls;
    logic         io_commits_info_3_mmio;
    logic [2:0]   io_commits_info_3_commitType;
    logic         io_commits_info_3_ftqIdx_flag;
    logic [5:0]   io_commits_info_3_ftqIdx_value;
    logic [3:0]   io_commits_info_3_ftqOffset;
    logic [2:0]   io_commits_info_3_instrSize;
    logic         io_commits_info_3_fpWen;
    logic         io_commits_info_3_rfWen;
    logic         io_commits_info_3_needFlush;
    logic [3:0]   io_commits_info_3_traceBlockInPipe_itype;
    logic [3:0]   io_commits_info_3_traceBlockInPipe_iretire;
    logic         io_commits_info_3_traceBlockInPipe_ilastsize;
    logic [49:0]  io_commits_info_3_debug_pc;
    logic [31:0]  io_commits_info_3_debug_instr;
    logic [5:0]   io_commits_info_3_debug_ldest;
    logic [7:0]   io_commits_info_3_debug_pdest;
    logic [7:0]   io_commits_info_3_debug_otherPdest_0;
    logic [7:0]   io_commits_info_3_debug_otherPdest_1;
    logic [7:0]   io_commits_info_3_debug_otherPdest_2;
    logic [7:0]   io_commits_info_3_debug_otherPdest_3;
    logic [7:0]   io_commits_info_3_debug_otherPdest_4;
    logic [7:0]   io_commits_info_3_debug_otherPdest_5;
    logic [7:0]   io_commits_info_3_debug_otherPdest_6;
    logic [34:0]  io_commits_info_3_debug_fuType;
    logic         io_commits_info_3_dirtyFs;
    logic         io_commits_info_3_dirtyVs;
    logic         io_commits_info_4_walk_v;
    logic         io_commits_info_4_commit_v;
    logic         io_commits_info_4_commit_w;
    logic [6:0]   io_commits_info_4_realDestSize;
    logic         io_commits_info_4_interrupt_safe;
    logic         io_commits_info_4_wflags;
    logic [4:0]   io_commits_info_4_fflags;
    logic         io_commits_info_4_vxsat;
    logic         io_commits_info_4_isRVC;
    logic         io_commits_info_4_isVset;
    logic         io_commits_info_4_isHls;
    logic         io_commits_info_4_isVls;
    logic         io_commits_info_4_vls;
    logic         io_commits_info_4_mmio;
    logic [2:0]   io_commits_info_4_commitType;
    logic         io_commits_info_4_ftqIdx_flag;
    logic [5:0]   io_commits_info_4_ftqIdx_value;
    logic [3:0]   io_commits_info_4_ftqOffset;
    logic [2:0]   io_commits_info_4_instrSize;
    logic         io_commits_info_4_fpWen;
    logic         io_commits_info_4_rfWen;
    logic         io_commits_info_4_needFlush;
    logic [3:0]   io_commits_info_4_traceBlockInPipe_itype;
    logic [3:0]   io_commits_info_4_traceBlockInPipe_iretire;
    logic         io_commits_info_4_traceBlockInPipe_ilastsize;
    logic [49:0]  io_commits_info_4_debug_pc;
    logic [31:0]  io_commits_info_4_debug_instr;
    logic [5:0]   io_commits_info_4_debug_ldest;
    logic [7:0]   io_commits_info_4_debug_pdest;
    logic [7:0]   io_commits_info_4_debug_otherPdest_0;
    logic [7:0]   io_commits_info_4_debug_otherPdest_1;
    logic [7:0]   io_commits_info_4_debug_otherPdest_2;
    logic [7:0]   io_commits_info_4_debug_otherPdest_3;
    logic [7:0]   io_commits_info_4_debug_otherPdest_4;
    logic [7:0]   io_commits_info_4_debug_otherPdest_5;
    logic [7:0]   io_commits_info_4_debug_otherPdest_6;
    logic [34:0]  io_commits_info_4_debug_fuType;
    logic         io_commits_info_4_dirtyFs;
    logic         io_commits_info_4_dirtyVs;
    logic         io_commits_info_5_walk_v;
    logic         io_commits_info_5_commit_v;
    logic         io_commits_info_5_commit_w;
    logic [6:0]   io_commits_info_5_realDestSize;
    logic         io_commits_info_5_interrupt_safe;
    logic         io_commits_info_5_wflags;
    logic [4:0]   io_commits_info_5_fflags;
    logic         io_commits_info_5_vxsat;
    logic         io_commits_info_5_isRVC;
    logic         io_commits_info_5_isVset;
    logic         io_commits_info_5_isHls;
    logic         io_commits_info_5_isVls;
    logic         io_commits_info_5_vls;
    logic         io_commits_info_5_mmio;
    logic [2:0]   io_commits_info_5_commitType;
    logic         io_commits_info_5_ftqIdx_flag;
    logic [5:0]   io_commits_info_5_ftqIdx_value;
    logic [3:0]   io_commits_info_5_ftqOffset;
    logic [2:0]   io_commits_info_5_instrSize;
    logic         io_commits_info_5_fpWen;
    logic         io_commits_info_5_rfWen;
    logic         io_commits_info_5_needFlush;
    logic [3:0]   io_commits_info_5_traceBlockInPipe_itype;
    logic [3:0]   io_commits_info_5_traceBlockInPipe_iretire;
    logic         io_commits_info_5_traceBlockInPipe_ilastsize;
    logic [49:0]  io_commits_info_5_debug_pc;
    logic [31:0]  io_commits_info_5_debug_instr;
    logic [5:0]   io_commits_info_5_debug_ldest;
    logic [7:0]   io_commits_info_5_debug_pdest;
    logic [7:0]   io_commits_info_5_debug_otherPdest_0;
    logic [7:0]   io_commits_info_5_debug_otherPdest_1;
    logic [7:0]   io_commits_info_5_debug_otherPdest_2;
    logic [7:0]   io_commits_info_5_debug_otherPdest_3;
    logic [7:0]   io_commits_info_5_debug_otherPdest_4;
    logic [7:0]   io_commits_info_5_debug_otherPdest_5;
    logic [7:0]   io_commits_info_5_debug_otherPdest_6;
    logic [34:0]  io_commits_info_5_debug_fuType;
    logic         io_commits_info_5_dirtyFs;
    logic         io_commits_info_5_dirtyVs;
    logic         io_commits_info_6_walk_v;
    logic         io_commits_info_6_commit_v;
    logic         io_commits_info_6_commit_w;
    logic [6:0]   io_commits_info_6_realDestSize;
    logic         io_commits_info_6_interrupt_safe;
    logic         io_commits_info_6_wflags;
    logic [4:0]   io_commits_info_6_fflags;
    logic         io_commits_info_6_vxsat;
    logic         io_commits_info_6_isRVC;
    logic         io_commits_info_6_isVset;
    logic         io_commits_info_6_isHls;
    logic         io_commits_info_6_isVls;
    logic         io_commits_info_6_vls;
    logic         io_commits_info_6_mmio;
    logic [2:0]   io_commits_info_6_commitType;
    logic         io_commits_info_6_ftqIdx_flag;
    logic [5:0]   io_commits_info_6_ftqIdx_value;
    logic [3:0]   io_commits_info_6_ftqOffset;
    logic [2:0]   io_commits_info_6_instrSize;
    logic         io_commits_info_6_fpWen;
    logic         io_commits_info_6_rfWen;
    logic         io_commits_info_6_needFlush;
    logic [3:0]   io_commits_info_6_traceBlockInPipe_itype;
    logic [3:0]   io_commits_info_6_traceBlockInPipe_iretire;
    logic         io_commits_info_6_traceBlockInPipe_ilastsize;
    logic [49:0]  io_commits_info_6_debug_pc;
    logic [31:0]  io_commits_info_6_debug_instr;
    logic [5:0]   io_commits_info_6_debug_ldest;
    logic [7:0]   io_commits_info_6_debug_pdest;
    logic [7:0]   io_commits_info_6_debug_otherPdest_0;
    logic [7:0]   io_commits_info_6_debug_otherPdest_1;
    logic [7:0]   io_commits_info_6_debug_otherPdest_2;
    logic [7:0]   io_commits_info_6_debug_otherPdest_3;
    logic [7:0]   io_commits_info_6_debug_otherPdest_4;
    logic [7:0]   io_commits_info_6_debug_otherPdest_5;
    logic [7:0]   io_commits_info_6_debug_otherPdest_6;
    logic [34:0]  io_commits_info_6_debug_fuType;
    logic         io_commits_info_6_dirtyFs;
    logic         io_commits_info_6_dirtyVs;
    logic         io_commits_info_7_walk_v;
    logic         io_commits_info_7_commit_v;
    logic         io_commits_info_7_commit_w;
    logic [6:0]   io_commits_info_7_realDestSize;
    logic         io_commits_info_7_interrupt_safe;
    logic         io_commits_info_7_wflags;
    logic [4:0]   io_commits_info_7_fflags;
    logic         io_commits_info_7_vxsat;
    logic         io_commits_info_7_isRVC;
    logic         io_commits_info_7_isVset;
    logic         io_commits_info_7_isHls;
    logic         io_commits_info_7_isVls;
    logic         io_commits_info_7_vls;
    logic         io_commits_info_7_mmio;
    logic [2:0]   io_commits_info_7_commitType;
    logic         io_commits_info_7_ftqIdx_flag;
    logic [5:0]   io_commits_info_7_ftqIdx_value;
    logic [3:0]   io_commits_info_7_ftqOffset;
    logic [2:0]   io_commits_info_7_instrSize;
    logic         io_commits_info_7_fpWen;
    logic         io_commits_info_7_rfWen;
    logic         io_commits_info_7_needFlush;
    logic [3:0]   io_commits_info_7_traceBlockInPipe_itype;
    logic [3:0]   io_commits_info_7_traceBlockInPipe_iretire;
    logic         io_commits_info_7_traceBlockInPipe_ilastsize;
    logic [49:0]  io_commits_info_7_debug_pc;
    logic [31:0]  io_commits_info_7_debug_instr;
    logic [5:0]   io_commits_info_7_debug_ldest;
    logic [7:0]   io_commits_info_7_debug_pdest;
    logic [7:0]   io_commits_info_7_debug_otherPdest_0;
    logic [7:0]   io_commits_info_7_debug_otherPdest_1;
    logic [7:0]   io_commits_info_7_debug_otherPdest_2;
    logic [7:0]   io_commits_info_7_debug_otherPdest_3;
    logic [7:0]   io_commits_info_7_debug_otherPdest_4;
    logic [7:0]   io_commits_info_7_debug_otherPdest_5;
    logic [7:0]   io_commits_info_7_debug_otherPdest_6;
    logic [34:0]  io_commits_info_7_debug_fuType;
    logic         io_commits_info_7_dirtyFs;
    logic         io_commits_info_7_dirtyVs;
    logic         io_commits_robIdx_0_flag;
    logic [7:0]   io_commits_robIdx_0_value;
    logic         io_commits_robIdx_1_flag;
    logic [7:0]   io_commits_robIdx_1_value;
    logic         io_commits_robIdx_2_flag;
    logic [7:0]   io_commits_robIdx_2_value;
    logic         io_commits_robIdx_3_flag;
    logic [7:0]   io_commits_robIdx_3_value;
    logic         io_commits_robIdx_4_flag;
    logic [7:0]   io_commits_robIdx_4_value;
    logic         io_commits_robIdx_5_flag;
    logic [7:0]   io_commits_robIdx_5_value;
    logic         io_commits_robIdx_6_flag;
    logic [7:0]   io_commits_robIdx_6_value;
    logic         io_commits_robIdx_7_flag;
    logic [7:0]   io_commits_robIdx_7_value;
    logic         io_trace_blockCommit ;
    logic         io_trace_traceCommitInfo_blocks_0_valid;
    logic [5:0]   io_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value;
    logic [3:0]   io_trace_traceCommitInfo_blocks_0_bits_ftqOffset;
    logic [3:0]   io_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype;
    logic [3:0]   io_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire;
    logic         io_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize;
    logic         io_trace_traceCommitInfo_blocks_1_valid;
    logic [5:0]   io_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value;
    logic [3:0]   io_trace_traceCommitInfo_blocks_1_bits_ftqOffset;
    logic [3:0]   io_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype;
    logic [3:0]   io_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire;
    logic         io_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize;
    logic         io_trace_traceCommitInfo_blocks_2_valid;
    logic [5:0]   io_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value;
    logic [3:0]   io_trace_traceCommitInfo_blocks_2_bits_ftqOffset;
    logic [3:0]   io_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype;
    logic [3:0]   io_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire;
    logic         io_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize;
    logic         io_trace_traceCommitInfo_blocks_3_valid;
    logic [5:0]   io_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value;
    logic [3:0]   io_trace_traceCommitInfo_blocks_3_bits_ftqOffset;
    logic [3:0]   io_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype;
    logic [3:0]   io_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire;
    logic         io_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize;
    logic         io_trace_traceCommitInfo_blocks_4_valid;
    logic [5:0]   io_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value;
    logic [3:0]   io_trace_traceCommitInfo_blocks_4_bits_ftqOffset;
    logic [3:0]   io_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype;
    logic [3:0]   io_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire;
    logic         io_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize;
    logic         io_trace_traceCommitInfo_blocks_5_valid;
    logic [5:0]   io_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value;
    logic [3:0]   io_trace_traceCommitInfo_blocks_5_bits_ftqOffset;
    logic [3:0]   io_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype;
    logic [3:0]   io_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire;
    logic         io_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize;
    logic         io_trace_traceCommitInfo_blocks_6_valid;
    logic [5:0]   io_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value;
    logic [3:0]   io_trace_traceCommitInfo_blocks_6_bits_ftqOffset;
    logic [3:0]   io_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype;
    logic [3:0]   io_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire;
    logic         io_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize;
    logic         io_trace_traceCommitInfo_blocks_7_valid;
    logic [5:0]   io_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value;
    logic [3:0]   io_trace_traceCommitInfo_blocks_7_bits_ftqOffset;
    logic [3:0]   io_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype;
    logic [3:0]   io_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire;
    logic         io_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize;
    logic         io_rabCommits_isCommit;
    logic         io_rabCommits_commitValid_0;
    logic         io_rabCommits_commitValid_1;
    logic         io_rabCommits_commitValid_2;
    logic         io_rabCommits_commitValid_3;
    logic         io_rabCommits_commitValid_4;
    logic         io_rabCommits_commitValid_5;
    logic         io_rabCommits_isWalk ;
    logic         io_rabCommits_walkValid_0;
    logic         io_rabCommits_walkValid_1;
    logic         io_rabCommits_walkValid_2;
    logic         io_rabCommits_walkValid_3;
    logic         io_rabCommits_walkValid_4;
    logic         io_rabCommits_walkValid_5;
    logic [5:0]   io_rabCommits_info_0_ldest;
    logic [7:0]   io_rabCommits_info_0_pdest;
    logic         io_rabCommits_info_0_rfWen;
    logic         io_rabCommits_info_0_fpWen;
    logic         io_rabCommits_info_0_vecWen;
    logic         io_rabCommits_info_0_v0Wen;
    logic         io_rabCommits_info_0_vlWen;
    logic         io_rabCommits_info_0_isMove;
    logic [5:0]   io_rabCommits_info_1_ldest;
    logic [7:0]   io_rabCommits_info_1_pdest;
    logic         io_rabCommits_info_1_rfWen;
    logic         io_rabCommits_info_1_fpWen;
    logic         io_rabCommits_info_1_vecWen;
    logic         io_rabCommits_info_1_v0Wen;
    logic         io_rabCommits_info_1_vlWen;
    logic         io_rabCommits_info_1_isMove;
    logic [5:0]   io_rabCommits_info_2_ldest;
    logic [7:0]   io_rabCommits_info_2_pdest;
    logic         io_rabCommits_info_2_rfWen;
    logic         io_rabCommits_info_2_fpWen;
    logic         io_rabCommits_info_2_vecWen;
    logic         io_rabCommits_info_2_v0Wen;
    logic         io_rabCommits_info_2_vlWen;
    logic         io_rabCommits_info_2_isMove;
    logic [5:0]   io_rabCommits_info_3_ldest;
    logic [7:0]   io_rabCommits_info_3_pdest;
    logic         io_rabCommits_info_3_rfWen;
    logic         io_rabCommits_info_3_fpWen;
    logic         io_rabCommits_info_3_vecWen;
    logic         io_rabCommits_info_3_v0Wen;
    logic         io_rabCommits_info_3_vlWen;
    logic         io_rabCommits_info_3_isMove;
    logic [5:0]   io_rabCommits_info_4_ldest;
    logic [7:0]   io_rabCommits_info_4_pdest;
    logic         io_rabCommits_info_4_rfWen;
    logic         io_rabCommits_info_4_fpWen;
    logic         io_rabCommits_info_4_vecWen;
    logic         io_rabCommits_info_4_v0Wen;
    logic         io_rabCommits_info_4_vlWen;
    logic         io_rabCommits_info_4_isMove;
    logic [5:0]   io_rabCommits_info_5_ldest;
    logic [7:0]   io_rabCommits_info_5_pdest;
    logic         io_rabCommits_info_5_rfWen;
    logic         io_rabCommits_info_5_fpWen;
    logic         io_rabCommits_info_5_vecWen;
    logic         io_rabCommits_info_5_v0Wen;
    logic         io_rabCommits_info_5_vlWen;
    logic         io_rabCommits_info_5_isMove;
    logic         io_diffCommits_commitValid_0;
    logic         io_diffCommits_commitValid_1;
    logic         io_diffCommits_commitValid_2;
    logic         io_diffCommits_commitValid_3;
    logic         io_diffCommits_commitValid_4;
    logic         io_diffCommits_commitValid_5;
    logic         io_diffCommits_commitValid_6;
    logic         io_diffCommits_commitValid_7;
    logic         io_diffCommits_commitValid_8;
    logic         io_diffCommits_commitValid_9;
    logic         io_diffCommits_commitValid_10;
    logic         io_diffCommits_commitValid_11;
    logic         io_diffCommits_commitValid_12;
    logic         io_diffCommits_commitValid_13;
    logic         io_diffCommits_commitValid_14;
    logic         io_diffCommits_commitValid_15;
    logic         io_diffCommits_commitValid_16;
    logic         io_diffCommits_commitValid_17;
    logic         io_diffCommits_commitValid_18;
    logic         io_diffCommits_commitValid_19;
    logic         io_diffCommits_commitValid_20;
    logic         io_diffCommits_commitValid_21;
    logic         io_diffCommits_commitValid_22;
    logic         io_diffCommits_commitValid_23;
    logic         io_diffCommits_commitValid_24;
    logic         io_diffCommits_commitValid_25;
    logic         io_diffCommits_commitValid_26;
    logic         io_diffCommits_commitValid_27;
    logic         io_diffCommits_commitValid_28;
    logic         io_diffCommits_commitValid_29;
    logic         io_diffCommits_commitValid_30;
    logic         io_diffCommits_commitValid_31;
    logic         io_diffCommits_commitValid_32;
    logic         io_diffCommits_commitValid_33;
    logic         io_diffCommits_commitValid_34;
    logic         io_diffCommits_commitValid_35;
    logic         io_diffCommits_commitValid_36;
    logic         io_diffCommits_commitValid_37;
    logic         io_diffCommits_commitValid_38;
    logic         io_diffCommits_commitValid_39;
    logic         io_diffCommits_commitValid_40;
    logic         io_diffCommits_commitValid_41;
    logic         io_diffCommits_commitValid_42;
    logic         io_diffCommits_commitValid_43;
    logic         io_diffCommits_commitValid_44;
    logic         io_diffCommits_commitValid_45;
    logic         io_diffCommits_commitValid_46;
    logic         io_diffCommits_commitValid_47;
    logic         io_diffCommits_commitValid_48;
    logic         io_diffCommits_commitValid_49;
    logic         io_diffCommits_commitValid_50;
    logic         io_diffCommits_commitValid_51;
    logic         io_diffCommits_commitValid_52;
    logic         io_diffCommits_commitValid_53;
    logic         io_diffCommits_commitValid_54;
    logic         io_diffCommits_commitValid_55;
    logic         io_diffCommits_commitValid_56;
    logic         io_diffCommits_commitValid_57;
    logic         io_diffCommits_commitValid_58;
    logic         io_diffCommits_commitValid_59;
    logic         io_diffCommits_commitValid_60;
    logic         io_diffCommits_commitValid_61;
    logic         io_diffCommits_commitValid_62;
    logic         io_diffCommits_commitValid_63;
    logic         io_diffCommits_commitValid_64;
    logic         io_diffCommits_commitValid_65;
    logic         io_diffCommits_commitValid_66;
    logic         io_diffCommits_commitValid_67;
    logic         io_diffCommits_commitValid_68;
    logic         io_diffCommits_commitValid_69;
    logic         io_diffCommits_commitValid_70;
    logic         io_diffCommits_commitValid_71;
    logic         io_diffCommits_commitValid_72;
    logic         io_diffCommits_commitValid_73;
    logic         io_diffCommits_commitValid_74;
    logic         io_diffCommits_commitValid_75;
    logic         io_diffCommits_commitValid_76;
    logic         io_diffCommits_commitValid_77;
    logic         io_diffCommits_commitValid_78;
    logic         io_diffCommits_commitValid_79;
    logic         io_diffCommits_commitValid_80;
    logic         io_diffCommits_commitValid_81;
    logic         io_diffCommits_commitValid_82;
    logic         io_diffCommits_commitValid_83;
    logic         io_diffCommits_commitValid_84;
    logic         io_diffCommits_commitValid_85;
    logic         io_diffCommits_commitValid_86;
    logic         io_diffCommits_commitValid_87;
    logic         io_diffCommits_commitValid_88;
    logic         io_diffCommits_commitValid_89;
    logic         io_diffCommits_commitValid_90;
    logic         io_diffCommits_commitValid_91;
    logic         io_diffCommits_commitValid_92;
    logic         io_diffCommits_commitValid_93;
    logic         io_diffCommits_commitValid_94;
    logic         io_diffCommits_commitValid_95;
    logic         io_diffCommits_commitValid_96;
    logic         io_diffCommits_commitValid_97;
    logic         io_diffCommits_commitValid_98;
    logic         io_diffCommits_commitValid_99;
    logic         io_diffCommits_commitValid_100;
    logic         io_diffCommits_commitValid_101;
    logic         io_diffCommits_commitValid_102;
    logic         io_diffCommits_commitValid_103;
    logic         io_diffCommits_commitValid_104;
    logic         io_diffCommits_commitValid_105;
    logic         io_diffCommits_commitValid_106;
    logic         io_diffCommits_commitValid_107;
    logic         io_diffCommits_commitValid_108;
    logic         io_diffCommits_commitValid_109;
    logic         io_diffCommits_commitValid_110;
    logic         io_diffCommits_commitValid_111;
    logic         io_diffCommits_commitValid_112;
    logic         io_diffCommits_commitValid_113;
    logic         io_diffCommits_commitValid_114;
    logic         io_diffCommits_commitValid_115;
    logic         io_diffCommits_commitValid_116;
    logic         io_diffCommits_commitValid_117;
    logic         io_diffCommits_commitValid_118;
    logic         io_diffCommits_commitValid_119;
    logic         io_diffCommits_commitValid_120;
    logic         io_diffCommits_commitValid_121;
    logic         io_diffCommits_commitValid_122;
    logic         io_diffCommits_commitValid_123;
    logic         io_diffCommits_commitValid_124;
    logic         io_diffCommits_commitValid_125;
    logic         io_diffCommits_commitValid_126;
    logic         io_diffCommits_commitValid_127;
    logic         io_diffCommits_commitValid_128;
    logic         io_diffCommits_commitValid_129;
    logic         io_diffCommits_commitValid_130;
    logic         io_diffCommits_commitValid_131;
    logic         io_diffCommits_commitValid_132;
    logic         io_diffCommits_commitValid_133;
    logic         io_diffCommits_commitValid_134;
    logic         io_diffCommits_commitValid_135;
    logic         io_diffCommits_commitValid_136;
    logic         io_diffCommits_commitValid_137;
    logic         io_diffCommits_commitValid_138;
    logic         io_diffCommits_commitValid_139;
    logic         io_diffCommits_commitValid_140;
    logic         io_diffCommits_commitValid_141;
    logic         io_diffCommits_commitValid_142;
    logic         io_diffCommits_commitValid_143;
    logic         io_diffCommits_commitValid_144;
    logic         io_diffCommits_commitValid_145;
    logic         io_diffCommits_commitValid_146;
    logic         io_diffCommits_commitValid_147;
    logic         io_diffCommits_commitValid_148;
    logic         io_diffCommits_commitValid_149;
    logic         io_diffCommits_commitValid_150;
    logic         io_diffCommits_commitValid_151;
    logic         io_diffCommits_commitValid_152;
    logic         io_diffCommits_commitValid_153;
    logic         io_diffCommits_commitValid_154;
    logic         io_diffCommits_commitValid_155;
    logic         io_diffCommits_commitValid_156;
    logic         io_diffCommits_commitValid_157;
    logic         io_diffCommits_commitValid_158;
    logic         io_diffCommits_commitValid_159;
    logic         io_diffCommits_commitValid_160;
    logic         io_diffCommits_commitValid_161;
    logic         io_diffCommits_commitValid_162;
    logic         io_diffCommits_commitValid_163;
    logic         io_diffCommits_commitValid_164;
    logic         io_diffCommits_commitValid_165;
    logic         io_diffCommits_commitValid_166;
    logic         io_diffCommits_commitValid_167;
    logic         io_diffCommits_commitValid_168;
    logic         io_diffCommits_commitValid_169;
    logic         io_diffCommits_commitValid_170;
    logic         io_diffCommits_commitValid_171;
    logic         io_diffCommits_commitValid_172;
    logic         io_diffCommits_commitValid_173;
    logic         io_diffCommits_commitValid_174;
    logic         io_diffCommits_commitValid_175;
    logic         io_diffCommits_commitValid_176;
    logic         io_diffCommits_commitValid_177;
    logic         io_diffCommits_commitValid_178;
    logic         io_diffCommits_commitValid_179;
    logic         io_diffCommits_commitValid_180;
    logic         io_diffCommits_commitValid_181;
    logic         io_diffCommits_commitValid_182;
    logic         io_diffCommits_commitValid_183;
    logic         io_diffCommits_commitValid_184;
    logic         io_diffCommits_commitValid_185;
    logic         io_diffCommits_commitValid_186;
    logic         io_diffCommits_commitValid_187;
    logic         io_diffCommits_commitValid_188;
    logic         io_diffCommits_commitValid_189;
    logic         io_diffCommits_commitValid_190;
    logic         io_diffCommits_commitValid_191;
    logic         io_diffCommits_commitValid_192;
    logic         io_diffCommits_commitValid_193;
    logic         io_diffCommits_commitValid_194;
    logic         io_diffCommits_commitValid_195;
    logic         io_diffCommits_commitValid_196;
    logic         io_diffCommits_commitValid_197;
    logic         io_diffCommits_commitValid_198;
    logic         io_diffCommits_commitValid_199;
    logic         io_diffCommits_commitValid_200;
    logic         io_diffCommits_commitValid_201;
    logic         io_diffCommits_commitValid_202;
    logic         io_diffCommits_commitValid_203;
    logic         io_diffCommits_commitValid_204;
    logic         io_diffCommits_commitValid_205;
    logic         io_diffCommits_commitValid_206;
    logic         io_diffCommits_commitValid_207;
    logic         io_diffCommits_commitValid_208;
    logic         io_diffCommits_commitValid_209;
    logic         io_diffCommits_commitValid_210;
    logic         io_diffCommits_commitValid_211;
    logic         io_diffCommits_commitValid_212;
    logic         io_diffCommits_commitValid_213;
    logic         io_diffCommits_commitValid_214;
    logic         io_diffCommits_commitValid_215;
    logic         io_diffCommits_commitValid_216;
    logic         io_diffCommits_commitValid_217;
    logic         io_diffCommits_commitValid_218;
    logic         io_diffCommits_commitValid_219;
    logic         io_diffCommits_commitValid_220;
    logic         io_diffCommits_commitValid_221;
    logic         io_diffCommits_commitValid_222;
    logic         io_diffCommits_commitValid_223;
    logic         io_diffCommits_commitValid_224;
    logic         io_diffCommits_commitValid_225;
    logic         io_diffCommits_commitValid_226;
    logic         io_diffCommits_commitValid_227;
    logic         io_diffCommits_commitValid_228;
    logic         io_diffCommits_commitValid_229;
    logic         io_diffCommits_commitValid_230;
    logic         io_diffCommits_commitValid_231;
    logic         io_diffCommits_commitValid_232;
    logic         io_diffCommits_commitValid_233;
    logic         io_diffCommits_commitValid_234;
    logic         io_diffCommits_commitValid_235;
    logic         io_diffCommits_commitValid_236;
    logic         io_diffCommits_commitValid_237;
    logic         io_diffCommits_commitValid_238;
    logic         io_diffCommits_commitValid_239;
    logic         io_diffCommits_commitValid_240;
    logic         io_diffCommits_commitValid_241;
    logic         io_diffCommits_commitValid_242;
    logic         io_diffCommits_commitValid_243;
    logic         io_diffCommits_commitValid_244;
    logic         io_diffCommits_commitValid_245;
    logic         io_diffCommits_commitValid_246;
    logic         io_diffCommits_commitValid_247;
    logic         io_diffCommits_commitValid_248;
    logic         io_diffCommits_commitValid_249;
    logic         io_diffCommits_commitValid_250;
    logic         io_diffCommits_commitValid_251;
    logic         io_diffCommits_commitValid_252;
    logic         io_diffCommits_commitValid_253;
    logic         io_diffCommits_commitValid_254;
    logic [5:0]   io_diffCommits_info_0_ldest;
    logic [7:0]   io_diffCommits_info_0_pdest;
    logic         io_diffCommits_info_0_rfWen;
    logic         io_diffCommits_info_0_fpWen;
    logic         io_diffCommits_info_0_vecWen;
    logic         io_diffCommits_info_0_v0Wen;
    logic         io_diffCommits_info_0_vlWen;
    logic [5:0]   io_diffCommits_info_1_ldest;
    logic [7:0]   io_diffCommits_info_1_pdest;
    logic         io_diffCommits_info_1_rfWen;
    logic         io_diffCommits_info_1_fpWen;
    logic         io_diffCommits_info_1_vecWen;
    logic         io_diffCommits_info_1_v0Wen;
    logic         io_diffCommits_info_1_vlWen;
    logic [5:0]   io_diffCommits_info_2_ldest;
    logic [7:0]   io_diffCommits_info_2_pdest;
    logic         io_diffCommits_info_2_rfWen;
    logic         io_diffCommits_info_2_fpWen;
    logic         io_diffCommits_info_2_vecWen;
    logic         io_diffCommits_info_2_v0Wen;
    logic         io_diffCommits_info_2_vlWen;
    logic [5:0]   io_diffCommits_info_3_ldest;
    logic [7:0]   io_diffCommits_info_3_pdest;
    logic         io_diffCommits_info_3_rfWen;
    logic         io_diffCommits_info_3_fpWen;
    logic         io_diffCommits_info_3_vecWen;
    logic         io_diffCommits_info_3_v0Wen;
    logic         io_diffCommits_info_3_vlWen;
    logic [5:0]   io_diffCommits_info_4_ldest;
    logic [7:0]   io_diffCommits_info_4_pdest;
    logic         io_diffCommits_info_4_rfWen;
    logic         io_diffCommits_info_4_fpWen;
    logic         io_diffCommits_info_4_vecWen;
    logic         io_diffCommits_info_4_v0Wen;
    logic         io_diffCommits_info_4_vlWen;
    logic [5:0]   io_diffCommits_info_5_ldest;
    logic [7:0]   io_diffCommits_info_5_pdest;
    logic         io_diffCommits_info_5_rfWen;
    logic         io_diffCommits_info_5_fpWen;
    logic         io_diffCommits_info_5_vecWen;
    logic         io_diffCommits_info_5_v0Wen;
    logic         io_diffCommits_info_5_vlWen;
    logic [5:0]   io_diffCommits_info_6_ldest;
    logic [7:0]   io_diffCommits_info_6_pdest;
    logic         io_diffCommits_info_6_rfWen;
    logic         io_diffCommits_info_6_fpWen;
    logic         io_diffCommits_info_6_vecWen;
    logic         io_diffCommits_info_6_v0Wen;
    logic         io_diffCommits_info_6_vlWen;
    logic [5:0]   io_diffCommits_info_7_ldest;
    logic [7:0]   io_diffCommits_info_7_pdest;
    logic         io_diffCommits_info_7_rfWen;
    logic         io_diffCommits_info_7_fpWen;
    logic         io_diffCommits_info_7_vecWen;
    logic         io_diffCommits_info_7_v0Wen;
    logic         io_diffCommits_info_7_vlWen;
    logic [5:0]   io_diffCommits_info_8_ldest;
    logic [7:0]   io_diffCommits_info_8_pdest;
    logic         io_diffCommits_info_8_rfWen;
    logic         io_diffCommits_info_8_fpWen;
    logic         io_diffCommits_info_8_vecWen;
    logic         io_diffCommits_info_8_v0Wen;
    logic         io_diffCommits_info_8_vlWen;
    logic [5:0]   io_diffCommits_info_9_ldest;
    logic [7:0]   io_diffCommits_info_9_pdest;
    logic         io_diffCommits_info_9_rfWen;
    logic         io_diffCommits_info_9_fpWen;
    logic         io_diffCommits_info_9_vecWen;
    logic         io_diffCommits_info_9_v0Wen;
    logic         io_diffCommits_info_9_vlWen;
    logic [5:0]   io_diffCommits_info_10_ldest;
    logic [7:0]   io_diffCommits_info_10_pdest;
    logic         io_diffCommits_info_10_rfWen;
    logic         io_diffCommits_info_10_fpWen;
    logic         io_diffCommits_info_10_vecWen;
    logic         io_diffCommits_info_10_v0Wen;
    logic         io_diffCommits_info_10_vlWen;
    logic [5:0]   io_diffCommits_info_11_ldest;
    logic [7:0]   io_diffCommits_info_11_pdest;
    logic         io_diffCommits_info_11_rfWen;
    logic         io_diffCommits_info_11_fpWen;
    logic         io_diffCommits_info_11_vecWen;
    logic         io_diffCommits_info_11_v0Wen;
    logic         io_diffCommits_info_11_vlWen;
    logic [5:0]   io_diffCommits_info_12_ldest;
    logic [7:0]   io_diffCommits_info_12_pdest;
    logic         io_diffCommits_info_12_rfWen;
    logic         io_diffCommits_info_12_fpWen;
    logic         io_diffCommits_info_12_vecWen;
    logic         io_diffCommits_info_12_v0Wen;
    logic         io_diffCommits_info_12_vlWen;
    logic [5:0]   io_diffCommits_info_13_ldest;
    logic [7:0]   io_diffCommits_info_13_pdest;
    logic         io_diffCommits_info_13_rfWen;
    logic         io_diffCommits_info_13_fpWen;
    logic         io_diffCommits_info_13_vecWen;
    logic         io_diffCommits_info_13_v0Wen;
    logic         io_diffCommits_info_13_vlWen;
    logic [5:0]   io_diffCommits_info_14_ldest;
    logic [7:0]   io_diffCommits_info_14_pdest;
    logic         io_diffCommits_info_14_rfWen;
    logic         io_diffCommits_info_14_fpWen;
    logic         io_diffCommits_info_14_vecWen;
    logic         io_diffCommits_info_14_v0Wen;
    logic         io_diffCommits_info_14_vlWen;
    logic [5:0]   io_diffCommits_info_15_ldest;
    logic [7:0]   io_diffCommits_info_15_pdest;
    logic         io_diffCommits_info_15_rfWen;
    logic         io_diffCommits_info_15_fpWen;
    logic         io_diffCommits_info_15_vecWen;
    logic         io_diffCommits_info_15_v0Wen;
    logic         io_diffCommits_info_15_vlWen;
    logic [5:0]   io_diffCommits_info_16_ldest;
    logic [7:0]   io_diffCommits_info_16_pdest;
    logic         io_diffCommits_info_16_rfWen;
    logic         io_diffCommits_info_16_fpWen;
    logic         io_diffCommits_info_16_vecWen;
    logic         io_diffCommits_info_16_v0Wen;
    logic         io_diffCommits_info_16_vlWen;
    logic [5:0]   io_diffCommits_info_17_ldest;
    logic [7:0]   io_diffCommits_info_17_pdest;
    logic         io_diffCommits_info_17_rfWen;
    logic         io_diffCommits_info_17_fpWen;
    logic         io_diffCommits_info_17_vecWen;
    logic         io_diffCommits_info_17_v0Wen;
    logic         io_diffCommits_info_17_vlWen;
    logic [5:0]   io_diffCommits_info_18_ldest;
    logic [7:0]   io_diffCommits_info_18_pdest;
    logic         io_diffCommits_info_18_rfWen;
    logic         io_diffCommits_info_18_fpWen;
    logic         io_diffCommits_info_18_vecWen;
    logic         io_diffCommits_info_18_v0Wen;
    logic         io_diffCommits_info_18_vlWen;
    logic [5:0]   io_diffCommits_info_19_ldest;
    logic [7:0]   io_diffCommits_info_19_pdest;
    logic         io_diffCommits_info_19_rfWen;
    logic         io_diffCommits_info_19_fpWen;
    logic         io_diffCommits_info_19_vecWen;
    logic         io_diffCommits_info_19_v0Wen;
    logic         io_diffCommits_info_19_vlWen;
    logic [5:0]   io_diffCommits_info_20_ldest;
    logic [7:0]   io_diffCommits_info_20_pdest;
    logic         io_diffCommits_info_20_rfWen;
    logic         io_diffCommits_info_20_fpWen;
    logic         io_diffCommits_info_20_vecWen;
    logic         io_diffCommits_info_20_v0Wen;
    logic         io_diffCommits_info_20_vlWen;
    logic [5:0]   io_diffCommits_info_21_ldest;
    logic [7:0]   io_diffCommits_info_21_pdest;
    logic         io_diffCommits_info_21_rfWen;
    logic         io_diffCommits_info_21_fpWen;
    logic         io_diffCommits_info_21_vecWen;
    logic         io_diffCommits_info_21_v0Wen;
    logic         io_diffCommits_info_21_vlWen;
    logic [5:0]   io_diffCommits_info_22_ldest;
    logic [7:0]   io_diffCommits_info_22_pdest;
    logic         io_diffCommits_info_22_rfWen;
    logic         io_diffCommits_info_22_fpWen;
    logic         io_diffCommits_info_22_vecWen;
    logic         io_diffCommits_info_22_v0Wen;
    logic         io_diffCommits_info_22_vlWen;
    logic [5:0]   io_diffCommits_info_23_ldest;
    logic [7:0]   io_diffCommits_info_23_pdest;
    logic         io_diffCommits_info_23_rfWen;
    logic         io_diffCommits_info_23_fpWen;
    logic         io_diffCommits_info_23_vecWen;
    logic         io_diffCommits_info_23_v0Wen;
    logic         io_diffCommits_info_23_vlWen;
    logic [5:0]   io_diffCommits_info_24_ldest;
    logic [7:0]   io_diffCommits_info_24_pdest;
    logic         io_diffCommits_info_24_rfWen;
    logic         io_diffCommits_info_24_fpWen;
    logic         io_diffCommits_info_24_vecWen;
    logic         io_diffCommits_info_24_v0Wen;
    logic         io_diffCommits_info_24_vlWen;
    logic [5:0]   io_diffCommits_info_25_ldest;
    logic [7:0]   io_diffCommits_info_25_pdest;
    logic         io_diffCommits_info_25_rfWen;
    logic         io_diffCommits_info_25_fpWen;
    logic         io_diffCommits_info_25_vecWen;
    logic         io_diffCommits_info_25_v0Wen;
    logic         io_diffCommits_info_25_vlWen;
    logic [5:0]   io_diffCommits_info_26_ldest;
    logic [7:0]   io_diffCommits_info_26_pdest;
    logic         io_diffCommits_info_26_rfWen;
    logic         io_diffCommits_info_26_fpWen;
    logic         io_diffCommits_info_26_vecWen;
    logic         io_diffCommits_info_26_v0Wen;
    logic         io_diffCommits_info_26_vlWen;
    logic [5:0]   io_diffCommits_info_27_ldest;
    logic [7:0]   io_diffCommits_info_27_pdest;
    logic         io_diffCommits_info_27_rfWen;
    logic         io_diffCommits_info_27_fpWen;
    logic         io_diffCommits_info_27_vecWen;
    logic         io_diffCommits_info_27_v0Wen;
    logic         io_diffCommits_info_27_vlWen;
    logic [5:0]   io_diffCommits_info_28_ldest;
    logic [7:0]   io_diffCommits_info_28_pdest;
    logic         io_diffCommits_info_28_rfWen;
    logic         io_diffCommits_info_28_fpWen;
    logic         io_diffCommits_info_28_vecWen;
    logic         io_diffCommits_info_28_v0Wen;
    logic         io_diffCommits_info_28_vlWen;
    logic [5:0]   io_diffCommits_info_29_ldest;
    logic [7:0]   io_diffCommits_info_29_pdest;
    logic         io_diffCommits_info_29_rfWen;
    logic         io_diffCommits_info_29_fpWen;
    logic         io_diffCommits_info_29_vecWen;
    logic         io_diffCommits_info_29_v0Wen;
    logic         io_diffCommits_info_29_vlWen;
    logic [5:0]   io_diffCommits_info_30_ldest;
    logic [7:0]   io_diffCommits_info_30_pdest;
    logic         io_diffCommits_info_30_rfWen;
    logic         io_diffCommits_info_30_fpWen;
    logic         io_diffCommits_info_30_vecWen;
    logic         io_diffCommits_info_30_v0Wen;
    logic         io_diffCommits_info_30_vlWen;
    logic [5:0]   io_diffCommits_info_31_ldest;
    logic [7:0]   io_diffCommits_info_31_pdest;
    logic         io_diffCommits_info_31_rfWen;
    logic         io_diffCommits_info_31_fpWen;
    logic         io_diffCommits_info_31_vecWen;
    logic         io_diffCommits_info_31_v0Wen;
    logic         io_diffCommits_info_31_vlWen;
    logic [5:0]   io_diffCommits_info_32_ldest;
    logic [7:0]   io_diffCommits_info_32_pdest;
    logic         io_diffCommits_info_32_rfWen;
    logic         io_diffCommits_info_32_fpWen;
    logic         io_diffCommits_info_32_vecWen;
    logic         io_diffCommits_info_32_v0Wen;
    logic         io_diffCommits_info_32_vlWen;
    logic [5:0]   io_diffCommits_info_33_ldest;
    logic [7:0]   io_diffCommits_info_33_pdest;
    logic         io_diffCommits_info_33_rfWen;
    logic         io_diffCommits_info_33_fpWen;
    logic         io_diffCommits_info_33_vecWen;
    logic         io_diffCommits_info_33_v0Wen;
    logic         io_diffCommits_info_33_vlWen;
    logic [5:0]   io_diffCommits_info_34_ldest;
    logic [7:0]   io_diffCommits_info_34_pdest;
    logic         io_diffCommits_info_34_rfWen;
    logic         io_diffCommits_info_34_fpWen;
    logic         io_diffCommits_info_34_vecWen;
    logic         io_diffCommits_info_34_v0Wen;
    logic         io_diffCommits_info_34_vlWen;
    logic [5:0]   io_diffCommits_info_35_ldest;
    logic [7:0]   io_diffCommits_info_35_pdest;
    logic         io_diffCommits_info_35_rfWen;
    logic         io_diffCommits_info_35_fpWen;
    logic         io_diffCommits_info_35_vecWen;
    logic         io_diffCommits_info_35_v0Wen;
    logic         io_diffCommits_info_35_vlWen;
    logic [5:0]   io_diffCommits_info_36_ldest;
    logic [7:0]   io_diffCommits_info_36_pdest;
    logic         io_diffCommits_info_36_rfWen;
    logic         io_diffCommits_info_36_fpWen;
    logic         io_diffCommits_info_36_vecWen;
    logic         io_diffCommits_info_36_v0Wen;
    logic         io_diffCommits_info_36_vlWen;
    logic [5:0]   io_diffCommits_info_37_ldest;
    logic [7:0]   io_diffCommits_info_37_pdest;
    logic         io_diffCommits_info_37_rfWen;
    logic         io_diffCommits_info_37_fpWen;
    logic         io_diffCommits_info_37_vecWen;
    logic         io_diffCommits_info_37_v0Wen;
    logic         io_diffCommits_info_37_vlWen;
    logic [5:0]   io_diffCommits_info_38_ldest;
    logic [7:0]   io_diffCommits_info_38_pdest;
    logic         io_diffCommits_info_38_rfWen;
    logic         io_diffCommits_info_38_fpWen;
    logic         io_diffCommits_info_38_vecWen;
    logic         io_diffCommits_info_38_v0Wen;
    logic         io_diffCommits_info_38_vlWen;
    logic [5:0]   io_diffCommits_info_39_ldest;
    logic [7:0]   io_diffCommits_info_39_pdest;
    logic         io_diffCommits_info_39_rfWen;
    logic         io_diffCommits_info_39_fpWen;
    logic         io_diffCommits_info_39_vecWen;
    logic         io_diffCommits_info_39_v0Wen;
    logic         io_diffCommits_info_39_vlWen;
    logic [5:0]   io_diffCommits_info_40_ldest;
    logic [7:0]   io_diffCommits_info_40_pdest;
    logic         io_diffCommits_info_40_rfWen;
    logic         io_diffCommits_info_40_fpWen;
    logic         io_diffCommits_info_40_vecWen;
    logic         io_diffCommits_info_40_v0Wen;
    logic         io_diffCommits_info_40_vlWen;
    logic [5:0]   io_diffCommits_info_41_ldest;
    logic [7:0]   io_diffCommits_info_41_pdest;
    logic         io_diffCommits_info_41_rfWen;
    logic         io_diffCommits_info_41_fpWen;
    logic         io_diffCommits_info_41_vecWen;
    logic         io_diffCommits_info_41_v0Wen;
    logic         io_diffCommits_info_41_vlWen;
    logic [5:0]   io_diffCommits_info_42_ldest;
    logic [7:0]   io_diffCommits_info_42_pdest;
    logic         io_diffCommits_info_42_rfWen;
    logic         io_diffCommits_info_42_fpWen;
    logic         io_diffCommits_info_42_vecWen;
    logic         io_diffCommits_info_42_v0Wen;
    logic         io_diffCommits_info_42_vlWen;
    logic [5:0]   io_diffCommits_info_43_ldest;
    logic [7:0]   io_diffCommits_info_43_pdest;
    logic         io_diffCommits_info_43_rfWen;
    logic         io_diffCommits_info_43_fpWen;
    logic         io_diffCommits_info_43_vecWen;
    logic         io_diffCommits_info_43_v0Wen;
    logic         io_diffCommits_info_43_vlWen;
    logic [5:0]   io_diffCommits_info_44_ldest;
    logic [7:0]   io_diffCommits_info_44_pdest;
    logic         io_diffCommits_info_44_rfWen;
    logic         io_diffCommits_info_44_fpWen;
    logic         io_diffCommits_info_44_vecWen;
    logic         io_diffCommits_info_44_v0Wen;
    logic         io_diffCommits_info_44_vlWen;
    logic [5:0]   io_diffCommits_info_45_ldest;
    logic [7:0]   io_diffCommits_info_45_pdest;
    logic         io_diffCommits_info_45_rfWen;
    logic         io_diffCommits_info_45_fpWen;
    logic         io_diffCommits_info_45_vecWen;
    logic         io_diffCommits_info_45_v0Wen;
    logic         io_diffCommits_info_45_vlWen;
    logic [5:0]   io_diffCommits_info_46_ldest;
    logic [7:0]   io_diffCommits_info_46_pdest;
    logic         io_diffCommits_info_46_rfWen;
    logic         io_diffCommits_info_46_fpWen;
    logic         io_diffCommits_info_46_vecWen;
    logic         io_diffCommits_info_46_v0Wen;
    logic         io_diffCommits_info_46_vlWen;
    logic [5:0]   io_diffCommits_info_47_ldest;
    logic [7:0]   io_diffCommits_info_47_pdest;
    logic         io_diffCommits_info_47_rfWen;
    logic         io_diffCommits_info_47_fpWen;
    logic         io_diffCommits_info_47_vecWen;
    logic         io_diffCommits_info_47_v0Wen;
    logic         io_diffCommits_info_47_vlWen;
    logic [5:0]   io_diffCommits_info_48_ldest;
    logic [7:0]   io_diffCommits_info_48_pdest;
    logic         io_diffCommits_info_48_rfWen;
    logic         io_diffCommits_info_48_fpWen;
    logic         io_diffCommits_info_48_vecWen;
    logic         io_diffCommits_info_48_v0Wen;
    logic         io_diffCommits_info_48_vlWen;
    logic [5:0]   io_diffCommits_info_49_ldest;
    logic [7:0]   io_diffCommits_info_49_pdest;
    logic         io_diffCommits_info_49_rfWen;
    logic         io_diffCommits_info_49_fpWen;
    logic         io_diffCommits_info_49_vecWen;
    logic         io_diffCommits_info_49_v0Wen;
    logic         io_diffCommits_info_49_vlWen;
    logic [5:0]   io_diffCommits_info_50_ldest;
    logic [7:0]   io_diffCommits_info_50_pdest;
    logic         io_diffCommits_info_50_rfWen;
    logic         io_diffCommits_info_50_fpWen;
    logic         io_diffCommits_info_50_vecWen;
    logic         io_diffCommits_info_50_v0Wen;
    logic         io_diffCommits_info_50_vlWen;
    logic [5:0]   io_diffCommits_info_51_ldest;
    logic [7:0]   io_diffCommits_info_51_pdest;
    logic         io_diffCommits_info_51_rfWen;
    logic         io_diffCommits_info_51_fpWen;
    logic         io_diffCommits_info_51_vecWen;
    logic         io_diffCommits_info_51_v0Wen;
    logic         io_diffCommits_info_51_vlWen;
    logic [5:0]   io_diffCommits_info_52_ldest;
    logic [7:0]   io_diffCommits_info_52_pdest;
    logic         io_diffCommits_info_52_rfWen;
    logic         io_diffCommits_info_52_fpWen;
    logic         io_diffCommits_info_52_vecWen;
    logic         io_diffCommits_info_52_v0Wen;
    logic         io_diffCommits_info_52_vlWen;
    logic [5:0]   io_diffCommits_info_53_ldest;
    logic [7:0]   io_diffCommits_info_53_pdest;
    logic         io_diffCommits_info_53_rfWen;
    logic         io_diffCommits_info_53_fpWen;
    logic         io_diffCommits_info_53_vecWen;
    logic         io_diffCommits_info_53_v0Wen;
    logic         io_diffCommits_info_53_vlWen;
    logic [5:0]   io_diffCommits_info_54_ldest;
    logic [7:0]   io_diffCommits_info_54_pdest;
    logic         io_diffCommits_info_54_rfWen;
    logic         io_diffCommits_info_54_fpWen;
    logic         io_diffCommits_info_54_vecWen;
    logic         io_diffCommits_info_54_v0Wen;
    logic         io_diffCommits_info_54_vlWen;
    logic [5:0]   io_diffCommits_info_55_ldest;
    logic [7:0]   io_diffCommits_info_55_pdest;
    logic         io_diffCommits_info_55_rfWen;
    logic         io_diffCommits_info_55_fpWen;
    logic         io_diffCommits_info_55_vecWen;
    logic         io_diffCommits_info_55_v0Wen;
    logic         io_diffCommits_info_55_vlWen;
    logic [5:0]   io_diffCommits_info_56_ldest;
    logic [7:0]   io_diffCommits_info_56_pdest;
    logic         io_diffCommits_info_56_rfWen;
    logic         io_diffCommits_info_56_fpWen;
    logic         io_diffCommits_info_56_vecWen;
    logic         io_diffCommits_info_56_v0Wen;
    logic         io_diffCommits_info_56_vlWen;
    logic [5:0]   io_diffCommits_info_57_ldest;
    logic [7:0]   io_diffCommits_info_57_pdest;
    logic         io_diffCommits_info_57_rfWen;
    logic         io_diffCommits_info_57_fpWen;
    logic         io_diffCommits_info_57_vecWen;
    logic         io_diffCommits_info_57_v0Wen;
    logic         io_diffCommits_info_57_vlWen;
    logic [5:0]   io_diffCommits_info_58_ldest;
    logic [7:0]   io_diffCommits_info_58_pdest;
    logic         io_diffCommits_info_58_rfWen;
    logic         io_diffCommits_info_58_fpWen;
    logic         io_diffCommits_info_58_vecWen;
    logic         io_diffCommits_info_58_v0Wen;
    logic         io_diffCommits_info_58_vlWen;
    logic [5:0]   io_diffCommits_info_59_ldest;
    logic [7:0]   io_diffCommits_info_59_pdest;
    logic         io_diffCommits_info_59_rfWen;
    logic         io_diffCommits_info_59_fpWen;
    logic         io_diffCommits_info_59_vecWen;
    logic         io_diffCommits_info_59_v0Wen;
    logic         io_diffCommits_info_59_vlWen;
    logic [5:0]   io_diffCommits_info_60_ldest;
    logic [7:0]   io_diffCommits_info_60_pdest;
    logic         io_diffCommits_info_60_rfWen;
    logic         io_diffCommits_info_60_fpWen;
    logic         io_diffCommits_info_60_vecWen;
    logic         io_diffCommits_info_60_v0Wen;
    logic         io_diffCommits_info_60_vlWen;
    logic [5:0]   io_diffCommits_info_61_ldest;
    logic [7:0]   io_diffCommits_info_61_pdest;
    logic         io_diffCommits_info_61_rfWen;
    logic         io_diffCommits_info_61_fpWen;
    logic         io_diffCommits_info_61_vecWen;
    logic         io_diffCommits_info_61_v0Wen;
    logic         io_diffCommits_info_61_vlWen;
    logic [5:0]   io_diffCommits_info_62_ldest;
    logic [7:0]   io_diffCommits_info_62_pdest;
    logic         io_diffCommits_info_62_rfWen;
    logic         io_diffCommits_info_62_fpWen;
    logic         io_diffCommits_info_62_vecWen;
    logic         io_diffCommits_info_62_v0Wen;
    logic         io_diffCommits_info_62_vlWen;
    logic [5:0]   io_diffCommits_info_63_ldest;
    logic [7:0]   io_diffCommits_info_63_pdest;
    logic         io_diffCommits_info_63_rfWen;
    logic         io_diffCommits_info_63_fpWen;
    logic         io_diffCommits_info_63_vecWen;
    logic         io_diffCommits_info_63_v0Wen;
    logic         io_diffCommits_info_63_vlWen;
    logic [5:0]   io_diffCommits_info_64_ldest;
    logic [7:0]   io_diffCommits_info_64_pdest;
    logic         io_diffCommits_info_64_rfWen;
    logic         io_diffCommits_info_64_fpWen;
    logic         io_diffCommits_info_64_vecWen;
    logic         io_diffCommits_info_64_v0Wen;
    logic         io_diffCommits_info_64_vlWen;
    logic [5:0]   io_diffCommits_info_65_ldest;
    logic [7:0]   io_diffCommits_info_65_pdest;
    logic         io_diffCommits_info_65_rfWen;
    logic         io_diffCommits_info_65_fpWen;
    logic         io_diffCommits_info_65_vecWen;
    logic         io_diffCommits_info_65_v0Wen;
    logic         io_diffCommits_info_65_vlWen;
    logic [5:0]   io_diffCommits_info_66_ldest;
    logic [7:0]   io_diffCommits_info_66_pdest;
    logic         io_diffCommits_info_66_rfWen;
    logic         io_diffCommits_info_66_fpWen;
    logic         io_diffCommits_info_66_vecWen;
    logic         io_diffCommits_info_66_v0Wen;
    logic         io_diffCommits_info_66_vlWen;
    logic [5:0]   io_diffCommits_info_67_ldest;
    logic [7:0]   io_diffCommits_info_67_pdest;
    logic         io_diffCommits_info_67_rfWen;
    logic         io_diffCommits_info_67_fpWen;
    logic         io_diffCommits_info_67_vecWen;
    logic         io_diffCommits_info_67_v0Wen;
    logic         io_diffCommits_info_67_vlWen;
    logic [5:0]   io_diffCommits_info_68_ldest;
    logic [7:0]   io_diffCommits_info_68_pdest;
    logic         io_diffCommits_info_68_rfWen;
    logic         io_diffCommits_info_68_fpWen;
    logic         io_diffCommits_info_68_vecWen;
    logic         io_diffCommits_info_68_v0Wen;
    logic         io_diffCommits_info_68_vlWen;
    logic [5:0]   io_diffCommits_info_69_ldest;
    logic [7:0]   io_diffCommits_info_69_pdest;
    logic         io_diffCommits_info_69_rfWen;
    logic         io_diffCommits_info_69_fpWen;
    logic         io_diffCommits_info_69_vecWen;
    logic         io_diffCommits_info_69_v0Wen;
    logic         io_diffCommits_info_69_vlWen;
    logic [5:0]   io_diffCommits_info_70_ldest;
    logic [7:0]   io_diffCommits_info_70_pdest;
    logic         io_diffCommits_info_70_rfWen;
    logic         io_diffCommits_info_70_fpWen;
    logic         io_diffCommits_info_70_vecWen;
    logic         io_diffCommits_info_70_v0Wen;
    logic         io_diffCommits_info_70_vlWen;
    logic [5:0]   io_diffCommits_info_71_ldest;
    logic [7:0]   io_diffCommits_info_71_pdest;
    logic         io_diffCommits_info_71_rfWen;
    logic         io_diffCommits_info_71_fpWen;
    logic         io_diffCommits_info_71_vecWen;
    logic         io_diffCommits_info_71_v0Wen;
    logic         io_diffCommits_info_71_vlWen;
    logic [5:0]   io_diffCommits_info_72_ldest;
    logic [7:0]   io_diffCommits_info_72_pdest;
    logic         io_diffCommits_info_72_rfWen;
    logic         io_diffCommits_info_72_fpWen;
    logic         io_diffCommits_info_72_vecWen;
    logic         io_diffCommits_info_72_v0Wen;
    logic         io_diffCommits_info_72_vlWen;
    logic [5:0]   io_diffCommits_info_73_ldest;
    logic [7:0]   io_diffCommits_info_73_pdest;
    logic         io_diffCommits_info_73_rfWen;
    logic         io_diffCommits_info_73_fpWen;
    logic         io_diffCommits_info_73_vecWen;
    logic         io_diffCommits_info_73_v0Wen;
    logic         io_diffCommits_info_73_vlWen;
    logic [5:0]   io_diffCommits_info_74_ldest;
    logic [7:0]   io_diffCommits_info_74_pdest;
    logic         io_diffCommits_info_74_rfWen;
    logic         io_diffCommits_info_74_fpWen;
    logic         io_diffCommits_info_74_vecWen;
    logic         io_diffCommits_info_74_v0Wen;
    logic         io_diffCommits_info_74_vlWen;
    logic [5:0]   io_diffCommits_info_75_ldest;
    logic [7:0]   io_diffCommits_info_75_pdest;
    logic         io_diffCommits_info_75_rfWen;
    logic         io_diffCommits_info_75_fpWen;
    logic         io_diffCommits_info_75_vecWen;
    logic         io_diffCommits_info_75_v0Wen;
    logic         io_diffCommits_info_75_vlWen;
    logic [5:0]   io_diffCommits_info_76_ldest;
    logic [7:0]   io_diffCommits_info_76_pdest;
    logic         io_diffCommits_info_76_rfWen;
    logic         io_diffCommits_info_76_fpWen;
    logic         io_diffCommits_info_76_vecWen;
    logic         io_diffCommits_info_76_v0Wen;
    logic         io_diffCommits_info_76_vlWen;
    logic [5:0]   io_diffCommits_info_77_ldest;
    logic [7:0]   io_diffCommits_info_77_pdest;
    logic         io_diffCommits_info_77_rfWen;
    logic         io_diffCommits_info_77_fpWen;
    logic         io_diffCommits_info_77_vecWen;
    logic         io_diffCommits_info_77_v0Wen;
    logic         io_diffCommits_info_77_vlWen;
    logic [5:0]   io_diffCommits_info_78_ldest;
    logic [7:0]   io_diffCommits_info_78_pdest;
    logic         io_diffCommits_info_78_rfWen;
    logic         io_diffCommits_info_78_fpWen;
    logic         io_diffCommits_info_78_vecWen;
    logic         io_diffCommits_info_78_v0Wen;
    logic         io_diffCommits_info_78_vlWen;
    logic [5:0]   io_diffCommits_info_79_ldest;
    logic [7:0]   io_diffCommits_info_79_pdest;
    logic         io_diffCommits_info_79_rfWen;
    logic         io_diffCommits_info_79_fpWen;
    logic         io_diffCommits_info_79_vecWen;
    logic         io_diffCommits_info_79_v0Wen;
    logic         io_diffCommits_info_79_vlWen;
    logic [5:0]   io_diffCommits_info_80_ldest;
    logic [7:0]   io_diffCommits_info_80_pdest;
    logic         io_diffCommits_info_80_rfWen;
    logic         io_diffCommits_info_80_fpWen;
    logic         io_diffCommits_info_80_vecWen;
    logic         io_diffCommits_info_80_v0Wen;
    logic         io_diffCommits_info_80_vlWen;
    logic [5:0]   io_diffCommits_info_81_ldest;
    logic [7:0]   io_diffCommits_info_81_pdest;
    logic         io_diffCommits_info_81_rfWen;
    logic         io_diffCommits_info_81_fpWen;
    logic         io_diffCommits_info_81_vecWen;
    logic         io_diffCommits_info_81_v0Wen;
    logic         io_diffCommits_info_81_vlWen;
    logic [5:0]   io_diffCommits_info_82_ldest;
    logic [7:0]   io_diffCommits_info_82_pdest;
    logic         io_diffCommits_info_82_rfWen;
    logic         io_diffCommits_info_82_fpWen;
    logic         io_diffCommits_info_82_vecWen;
    logic         io_diffCommits_info_82_v0Wen;
    logic         io_diffCommits_info_82_vlWen;
    logic [5:0]   io_diffCommits_info_83_ldest;
    logic [7:0]   io_diffCommits_info_83_pdest;
    logic         io_diffCommits_info_83_rfWen;
    logic         io_diffCommits_info_83_fpWen;
    logic         io_diffCommits_info_83_vecWen;
    logic         io_diffCommits_info_83_v0Wen;
    logic         io_diffCommits_info_83_vlWen;
    logic [5:0]   io_diffCommits_info_84_ldest;
    logic [7:0]   io_diffCommits_info_84_pdest;
    logic         io_diffCommits_info_84_rfWen;
    logic         io_diffCommits_info_84_fpWen;
    logic         io_diffCommits_info_84_vecWen;
    logic         io_diffCommits_info_84_v0Wen;
    logic         io_diffCommits_info_84_vlWen;
    logic [5:0]   io_diffCommits_info_85_ldest;
    logic [7:0]   io_diffCommits_info_85_pdest;
    logic         io_diffCommits_info_85_rfWen;
    logic         io_diffCommits_info_85_fpWen;
    logic         io_diffCommits_info_85_vecWen;
    logic         io_diffCommits_info_85_v0Wen;
    logic         io_diffCommits_info_85_vlWen;
    logic [5:0]   io_diffCommits_info_86_ldest;
    logic [7:0]   io_diffCommits_info_86_pdest;
    logic         io_diffCommits_info_86_rfWen;
    logic         io_diffCommits_info_86_fpWen;
    logic         io_diffCommits_info_86_vecWen;
    logic         io_diffCommits_info_86_v0Wen;
    logic         io_diffCommits_info_86_vlWen;
    logic [5:0]   io_diffCommits_info_87_ldest;
    logic [7:0]   io_diffCommits_info_87_pdest;
    logic         io_diffCommits_info_87_rfWen;
    logic         io_diffCommits_info_87_fpWen;
    logic         io_diffCommits_info_87_vecWen;
    logic         io_diffCommits_info_87_v0Wen;
    logic         io_diffCommits_info_87_vlWen;
    logic [5:0]   io_diffCommits_info_88_ldest;
    logic [7:0]   io_diffCommits_info_88_pdest;
    logic         io_diffCommits_info_88_rfWen;
    logic         io_diffCommits_info_88_fpWen;
    logic         io_diffCommits_info_88_vecWen;
    logic         io_diffCommits_info_88_v0Wen;
    logic         io_diffCommits_info_88_vlWen;
    logic [5:0]   io_diffCommits_info_89_ldest;
    logic [7:0]   io_diffCommits_info_89_pdest;
    logic         io_diffCommits_info_89_rfWen;
    logic         io_diffCommits_info_89_fpWen;
    logic         io_diffCommits_info_89_vecWen;
    logic         io_diffCommits_info_89_v0Wen;
    logic         io_diffCommits_info_89_vlWen;
    logic [5:0]   io_diffCommits_info_90_ldest;
    logic [7:0]   io_diffCommits_info_90_pdest;
    logic         io_diffCommits_info_90_rfWen;
    logic         io_diffCommits_info_90_fpWen;
    logic         io_diffCommits_info_90_vecWen;
    logic         io_diffCommits_info_90_v0Wen;
    logic         io_diffCommits_info_90_vlWen;
    logic [5:0]   io_diffCommits_info_91_ldest;
    logic [7:0]   io_diffCommits_info_91_pdest;
    logic         io_diffCommits_info_91_rfWen;
    logic         io_diffCommits_info_91_fpWen;
    logic         io_diffCommits_info_91_vecWen;
    logic         io_diffCommits_info_91_v0Wen;
    logic         io_diffCommits_info_91_vlWen;
    logic [5:0]   io_diffCommits_info_92_ldest;
    logic [7:0]   io_diffCommits_info_92_pdest;
    logic         io_diffCommits_info_92_rfWen;
    logic         io_diffCommits_info_92_fpWen;
    logic         io_diffCommits_info_92_vecWen;
    logic         io_diffCommits_info_92_v0Wen;
    logic         io_diffCommits_info_92_vlWen;
    logic [5:0]   io_diffCommits_info_93_ldest;
    logic [7:0]   io_diffCommits_info_93_pdest;
    logic         io_diffCommits_info_93_rfWen;
    logic         io_diffCommits_info_93_fpWen;
    logic         io_diffCommits_info_93_vecWen;
    logic         io_diffCommits_info_93_v0Wen;
    logic         io_diffCommits_info_93_vlWen;
    logic [5:0]   io_diffCommits_info_94_ldest;
    logic [7:0]   io_diffCommits_info_94_pdest;
    logic         io_diffCommits_info_94_rfWen;
    logic         io_diffCommits_info_94_fpWen;
    logic         io_diffCommits_info_94_vecWen;
    logic         io_diffCommits_info_94_v0Wen;
    logic         io_diffCommits_info_94_vlWen;
    logic [5:0]   io_diffCommits_info_95_ldest;
    logic [7:0]   io_diffCommits_info_95_pdest;
    logic         io_diffCommits_info_95_rfWen;
    logic         io_diffCommits_info_95_fpWen;
    logic         io_diffCommits_info_95_vecWen;
    logic         io_diffCommits_info_95_v0Wen;
    logic         io_diffCommits_info_95_vlWen;
    logic [5:0]   io_diffCommits_info_96_ldest;
    logic [7:0]   io_diffCommits_info_96_pdest;
    logic         io_diffCommits_info_96_rfWen;
    logic         io_diffCommits_info_96_fpWen;
    logic         io_diffCommits_info_96_vecWen;
    logic         io_diffCommits_info_96_v0Wen;
    logic         io_diffCommits_info_96_vlWen;
    logic [5:0]   io_diffCommits_info_97_ldest;
    logic [7:0]   io_diffCommits_info_97_pdest;
    logic         io_diffCommits_info_97_rfWen;
    logic         io_diffCommits_info_97_fpWen;
    logic         io_diffCommits_info_97_vecWen;
    logic         io_diffCommits_info_97_v0Wen;
    logic         io_diffCommits_info_97_vlWen;
    logic [5:0]   io_diffCommits_info_98_ldest;
    logic [7:0]   io_diffCommits_info_98_pdest;
    logic         io_diffCommits_info_98_rfWen;
    logic         io_diffCommits_info_98_fpWen;
    logic         io_diffCommits_info_98_vecWen;
    logic         io_diffCommits_info_98_v0Wen;
    logic         io_diffCommits_info_98_vlWen;
    logic [5:0]   io_diffCommits_info_99_ldest;
    logic [7:0]   io_diffCommits_info_99_pdest;
    logic         io_diffCommits_info_99_rfWen;
    logic         io_diffCommits_info_99_fpWen;
    logic         io_diffCommits_info_99_vecWen;
    logic         io_diffCommits_info_99_v0Wen;
    logic         io_diffCommits_info_99_vlWen;
    logic [5:0]   io_diffCommits_info_100_ldest;
    logic [7:0]   io_diffCommits_info_100_pdest;
    logic         io_diffCommits_info_100_rfWen;
    logic         io_diffCommits_info_100_fpWen;
    logic         io_diffCommits_info_100_vecWen;
    logic         io_diffCommits_info_100_v0Wen;
    logic         io_diffCommits_info_100_vlWen;
    logic [5:0]   io_diffCommits_info_101_ldest;
    logic [7:0]   io_diffCommits_info_101_pdest;
    logic         io_diffCommits_info_101_rfWen;
    logic         io_diffCommits_info_101_fpWen;
    logic         io_diffCommits_info_101_vecWen;
    logic         io_diffCommits_info_101_v0Wen;
    logic         io_diffCommits_info_101_vlWen;
    logic [5:0]   io_diffCommits_info_102_ldest;
    logic [7:0]   io_diffCommits_info_102_pdest;
    logic         io_diffCommits_info_102_rfWen;
    logic         io_diffCommits_info_102_fpWen;
    logic         io_diffCommits_info_102_vecWen;
    logic         io_diffCommits_info_102_v0Wen;
    logic         io_diffCommits_info_102_vlWen;
    logic [5:0]   io_diffCommits_info_103_ldest;
    logic [7:0]   io_diffCommits_info_103_pdest;
    logic         io_diffCommits_info_103_rfWen;
    logic         io_diffCommits_info_103_fpWen;
    logic         io_diffCommits_info_103_vecWen;
    logic         io_diffCommits_info_103_v0Wen;
    logic         io_diffCommits_info_103_vlWen;
    logic [5:0]   io_diffCommits_info_104_ldest;
    logic [7:0]   io_diffCommits_info_104_pdest;
    logic         io_diffCommits_info_104_rfWen;
    logic         io_diffCommits_info_104_fpWen;
    logic         io_diffCommits_info_104_vecWen;
    logic         io_diffCommits_info_104_v0Wen;
    logic         io_diffCommits_info_104_vlWen;
    logic [5:0]   io_diffCommits_info_105_ldest;
    logic [7:0]   io_diffCommits_info_105_pdest;
    logic         io_diffCommits_info_105_rfWen;
    logic         io_diffCommits_info_105_fpWen;
    logic         io_diffCommits_info_105_vecWen;
    logic         io_diffCommits_info_105_v0Wen;
    logic         io_diffCommits_info_105_vlWen;
    logic [5:0]   io_diffCommits_info_106_ldest;
    logic [7:0]   io_diffCommits_info_106_pdest;
    logic         io_diffCommits_info_106_rfWen;
    logic         io_diffCommits_info_106_fpWen;
    logic         io_diffCommits_info_106_vecWen;
    logic         io_diffCommits_info_106_v0Wen;
    logic         io_diffCommits_info_106_vlWen;
    logic [5:0]   io_diffCommits_info_107_ldest;
    logic [7:0]   io_diffCommits_info_107_pdest;
    logic         io_diffCommits_info_107_rfWen;
    logic         io_diffCommits_info_107_fpWen;
    logic         io_diffCommits_info_107_vecWen;
    logic         io_diffCommits_info_107_v0Wen;
    logic         io_diffCommits_info_107_vlWen;
    logic [5:0]   io_diffCommits_info_108_ldest;
    logic [7:0]   io_diffCommits_info_108_pdest;
    logic         io_diffCommits_info_108_rfWen;
    logic         io_diffCommits_info_108_fpWen;
    logic         io_diffCommits_info_108_vecWen;
    logic         io_diffCommits_info_108_v0Wen;
    logic         io_diffCommits_info_108_vlWen;
    logic [5:0]   io_diffCommits_info_109_ldest;
    logic [7:0]   io_diffCommits_info_109_pdest;
    logic         io_diffCommits_info_109_rfWen;
    logic         io_diffCommits_info_109_fpWen;
    logic         io_diffCommits_info_109_vecWen;
    logic         io_diffCommits_info_109_v0Wen;
    logic         io_diffCommits_info_109_vlWen;
    logic [5:0]   io_diffCommits_info_110_ldest;
    logic [7:0]   io_diffCommits_info_110_pdest;
    logic         io_diffCommits_info_110_rfWen;
    logic         io_diffCommits_info_110_fpWen;
    logic         io_diffCommits_info_110_vecWen;
    logic         io_diffCommits_info_110_v0Wen;
    logic         io_diffCommits_info_110_vlWen;
    logic [5:0]   io_diffCommits_info_111_ldest;
    logic [7:0]   io_diffCommits_info_111_pdest;
    logic         io_diffCommits_info_111_rfWen;
    logic         io_diffCommits_info_111_fpWen;
    logic         io_diffCommits_info_111_vecWen;
    logic         io_diffCommits_info_111_v0Wen;
    logic         io_diffCommits_info_111_vlWen;
    logic [5:0]   io_diffCommits_info_112_ldest;
    logic [7:0]   io_diffCommits_info_112_pdest;
    logic         io_diffCommits_info_112_rfWen;
    logic         io_diffCommits_info_112_fpWen;
    logic         io_diffCommits_info_112_vecWen;
    logic         io_diffCommits_info_112_v0Wen;
    logic         io_diffCommits_info_112_vlWen;
    logic [5:0]   io_diffCommits_info_113_ldest;
    logic [7:0]   io_diffCommits_info_113_pdest;
    logic         io_diffCommits_info_113_rfWen;
    logic         io_diffCommits_info_113_fpWen;
    logic         io_diffCommits_info_113_vecWen;
    logic         io_diffCommits_info_113_v0Wen;
    logic         io_diffCommits_info_113_vlWen;
    logic [5:0]   io_diffCommits_info_114_ldest;
    logic [7:0]   io_diffCommits_info_114_pdest;
    logic         io_diffCommits_info_114_rfWen;
    logic         io_diffCommits_info_114_fpWen;
    logic         io_diffCommits_info_114_vecWen;
    logic         io_diffCommits_info_114_v0Wen;
    logic         io_diffCommits_info_114_vlWen;
    logic [5:0]   io_diffCommits_info_115_ldest;
    logic [7:0]   io_diffCommits_info_115_pdest;
    logic         io_diffCommits_info_115_rfWen;
    logic         io_diffCommits_info_115_fpWen;
    logic         io_diffCommits_info_115_vecWen;
    logic         io_diffCommits_info_115_v0Wen;
    logic         io_diffCommits_info_115_vlWen;
    logic [5:0]   io_diffCommits_info_116_ldest;
    logic [7:0]   io_diffCommits_info_116_pdest;
    logic         io_diffCommits_info_116_rfWen;
    logic         io_diffCommits_info_116_fpWen;
    logic         io_diffCommits_info_116_vecWen;
    logic         io_diffCommits_info_116_v0Wen;
    logic         io_diffCommits_info_116_vlWen;
    logic [5:0]   io_diffCommits_info_117_ldest;
    logic [7:0]   io_diffCommits_info_117_pdest;
    logic         io_diffCommits_info_117_rfWen;
    logic         io_diffCommits_info_117_fpWen;
    logic         io_diffCommits_info_117_vecWen;
    logic         io_diffCommits_info_117_v0Wen;
    logic         io_diffCommits_info_117_vlWen;
    logic [5:0]   io_diffCommits_info_118_ldest;
    logic [7:0]   io_diffCommits_info_118_pdest;
    logic         io_diffCommits_info_118_rfWen;
    logic         io_diffCommits_info_118_fpWen;
    logic         io_diffCommits_info_118_vecWen;
    logic         io_diffCommits_info_118_v0Wen;
    logic         io_diffCommits_info_118_vlWen;
    logic [5:0]   io_diffCommits_info_119_ldest;
    logic [7:0]   io_diffCommits_info_119_pdest;
    logic         io_diffCommits_info_119_rfWen;
    logic         io_diffCommits_info_119_fpWen;
    logic         io_diffCommits_info_119_vecWen;
    logic         io_diffCommits_info_119_v0Wen;
    logic         io_diffCommits_info_119_vlWen;
    logic [5:0]   io_diffCommits_info_120_ldest;
    logic [7:0]   io_diffCommits_info_120_pdest;
    logic         io_diffCommits_info_120_rfWen;
    logic         io_diffCommits_info_120_fpWen;
    logic         io_diffCommits_info_120_vecWen;
    logic         io_diffCommits_info_120_v0Wen;
    logic         io_diffCommits_info_120_vlWen;
    logic [5:0]   io_diffCommits_info_121_ldest;
    logic [7:0]   io_diffCommits_info_121_pdest;
    logic         io_diffCommits_info_121_rfWen;
    logic         io_diffCommits_info_121_fpWen;
    logic         io_diffCommits_info_121_vecWen;
    logic         io_diffCommits_info_121_v0Wen;
    logic         io_diffCommits_info_121_vlWen;
    logic [5:0]   io_diffCommits_info_122_ldest;
    logic [7:0]   io_diffCommits_info_122_pdest;
    logic         io_diffCommits_info_122_rfWen;
    logic         io_diffCommits_info_122_fpWen;
    logic         io_diffCommits_info_122_vecWen;
    logic         io_diffCommits_info_122_v0Wen;
    logic         io_diffCommits_info_122_vlWen;
    logic [5:0]   io_diffCommits_info_123_ldest;
    logic [7:0]   io_diffCommits_info_123_pdest;
    logic         io_diffCommits_info_123_rfWen;
    logic         io_diffCommits_info_123_fpWen;
    logic         io_diffCommits_info_123_vecWen;
    logic         io_diffCommits_info_123_v0Wen;
    logic         io_diffCommits_info_123_vlWen;
    logic [5:0]   io_diffCommits_info_124_ldest;
    logic [7:0]   io_diffCommits_info_124_pdest;
    logic         io_diffCommits_info_124_rfWen;
    logic         io_diffCommits_info_124_fpWen;
    logic         io_diffCommits_info_124_vecWen;
    logic         io_diffCommits_info_124_v0Wen;
    logic         io_diffCommits_info_124_vlWen;
    logic [5:0]   io_diffCommits_info_125_ldest;
    logic [7:0]   io_diffCommits_info_125_pdest;
    logic         io_diffCommits_info_125_rfWen;
    logic         io_diffCommits_info_125_fpWen;
    logic         io_diffCommits_info_125_vecWen;
    logic         io_diffCommits_info_125_v0Wen;
    logic         io_diffCommits_info_125_vlWen;
    logic [5:0]   io_diffCommits_info_126_ldest;
    logic [7:0]   io_diffCommits_info_126_pdest;
    logic         io_diffCommits_info_126_rfWen;
    logic         io_diffCommits_info_126_fpWen;
    logic         io_diffCommits_info_126_vecWen;
    logic         io_diffCommits_info_126_v0Wen;
    logic         io_diffCommits_info_126_vlWen;
    logic [5:0]   io_diffCommits_info_127_ldest;
    logic [7:0]   io_diffCommits_info_127_pdest;
    logic         io_diffCommits_info_127_rfWen;
    logic         io_diffCommits_info_127_fpWen;
    logic         io_diffCommits_info_127_vecWen;
    logic         io_diffCommits_info_127_v0Wen;
    logic         io_diffCommits_info_127_vlWen;
    logic [5:0]   io_diffCommits_info_128_ldest;
    logic [7:0]   io_diffCommits_info_128_pdest;
    logic         io_diffCommits_info_128_rfWen;
    logic         io_diffCommits_info_128_fpWen;
    logic         io_diffCommits_info_128_vecWen;
    logic         io_diffCommits_info_128_v0Wen;
    logic         io_diffCommits_info_128_vlWen;
    logic [5:0]   io_diffCommits_info_129_ldest;
    logic [7:0]   io_diffCommits_info_129_pdest;
    logic         io_diffCommits_info_129_rfWen;
    logic         io_diffCommits_info_129_fpWen;
    logic         io_diffCommits_info_129_vecWen;
    logic         io_diffCommits_info_129_v0Wen;
    logic         io_diffCommits_info_129_vlWen;
    logic [5:0]   io_diffCommits_info_130_ldest;
    logic [7:0]   io_diffCommits_info_130_pdest;
    logic         io_diffCommits_info_130_rfWen;
    logic         io_diffCommits_info_130_fpWen;
    logic         io_diffCommits_info_130_vecWen;
    logic         io_diffCommits_info_130_v0Wen;
    logic         io_diffCommits_info_130_vlWen;
    logic [5:0]   io_diffCommits_info_131_ldest;
    logic [7:0]   io_diffCommits_info_131_pdest;
    logic         io_diffCommits_info_131_rfWen;
    logic         io_diffCommits_info_131_fpWen;
    logic         io_diffCommits_info_131_vecWen;
    logic         io_diffCommits_info_131_v0Wen;
    logic         io_diffCommits_info_131_vlWen;
    logic [5:0]   io_diffCommits_info_132_ldest;
    logic [7:0]   io_diffCommits_info_132_pdest;
    logic         io_diffCommits_info_132_rfWen;
    logic         io_diffCommits_info_132_fpWen;
    logic         io_diffCommits_info_132_vecWen;
    logic         io_diffCommits_info_132_v0Wen;
    logic         io_diffCommits_info_132_vlWen;
    logic [5:0]   io_diffCommits_info_133_ldest;
    logic [7:0]   io_diffCommits_info_133_pdest;
    logic         io_diffCommits_info_133_rfWen;
    logic         io_diffCommits_info_133_fpWen;
    logic         io_diffCommits_info_133_vecWen;
    logic         io_diffCommits_info_133_v0Wen;
    logic         io_diffCommits_info_133_vlWen;
    logic [5:0]   io_diffCommits_info_134_ldest;
    logic [7:0]   io_diffCommits_info_134_pdest;
    logic         io_diffCommits_info_134_rfWen;
    logic         io_diffCommits_info_134_fpWen;
    logic         io_diffCommits_info_134_vecWen;
    logic         io_diffCommits_info_134_v0Wen;
    logic         io_diffCommits_info_134_vlWen;
    logic [5:0]   io_diffCommits_info_135_ldest;
    logic [7:0]   io_diffCommits_info_135_pdest;
    logic         io_diffCommits_info_135_rfWen;
    logic         io_diffCommits_info_135_fpWen;
    logic         io_diffCommits_info_135_vecWen;
    logic         io_diffCommits_info_135_v0Wen;
    logic         io_diffCommits_info_135_vlWen;
    logic [5:0]   io_diffCommits_info_136_ldest;
    logic [7:0]   io_diffCommits_info_136_pdest;
    logic         io_diffCommits_info_136_rfWen;
    logic         io_diffCommits_info_136_fpWen;
    logic         io_diffCommits_info_136_vecWen;
    logic         io_diffCommits_info_136_v0Wen;
    logic         io_diffCommits_info_136_vlWen;
    logic [5:0]   io_diffCommits_info_137_ldest;
    logic [7:0]   io_diffCommits_info_137_pdest;
    logic         io_diffCommits_info_137_rfWen;
    logic         io_diffCommits_info_137_fpWen;
    logic         io_diffCommits_info_137_vecWen;
    logic         io_diffCommits_info_137_v0Wen;
    logic         io_diffCommits_info_137_vlWen;
    logic [5:0]   io_diffCommits_info_138_ldest;
    logic [7:0]   io_diffCommits_info_138_pdest;
    logic         io_diffCommits_info_138_rfWen;
    logic         io_diffCommits_info_138_fpWen;
    logic         io_diffCommits_info_138_vecWen;
    logic         io_diffCommits_info_138_v0Wen;
    logic         io_diffCommits_info_138_vlWen;
    logic [5:0]   io_diffCommits_info_139_ldest;
    logic [7:0]   io_diffCommits_info_139_pdest;
    logic         io_diffCommits_info_139_rfWen;
    logic         io_diffCommits_info_139_fpWen;
    logic         io_diffCommits_info_139_vecWen;
    logic         io_diffCommits_info_139_v0Wen;
    logic         io_diffCommits_info_139_vlWen;
    logic [5:0]   io_diffCommits_info_140_ldest;
    logic [7:0]   io_diffCommits_info_140_pdest;
    logic         io_diffCommits_info_140_rfWen;
    logic         io_diffCommits_info_140_fpWen;
    logic         io_diffCommits_info_140_vecWen;
    logic         io_diffCommits_info_140_v0Wen;
    logic         io_diffCommits_info_140_vlWen;
    logic [5:0]   io_diffCommits_info_141_ldest;
    logic [7:0]   io_diffCommits_info_141_pdest;
    logic         io_diffCommits_info_141_rfWen;
    logic         io_diffCommits_info_141_fpWen;
    logic         io_diffCommits_info_141_vecWen;
    logic         io_diffCommits_info_141_v0Wen;
    logic         io_diffCommits_info_141_vlWen;
    logic [5:0]   io_diffCommits_info_142_ldest;
    logic [7:0]   io_diffCommits_info_142_pdest;
    logic         io_diffCommits_info_142_rfWen;
    logic         io_diffCommits_info_142_fpWen;
    logic         io_diffCommits_info_142_vecWen;
    logic         io_diffCommits_info_142_v0Wen;
    logic         io_diffCommits_info_142_vlWen;
    logic [5:0]   io_diffCommits_info_143_ldest;
    logic [7:0]   io_diffCommits_info_143_pdest;
    logic         io_diffCommits_info_143_rfWen;
    logic         io_diffCommits_info_143_fpWen;
    logic         io_diffCommits_info_143_vecWen;
    logic         io_diffCommits_info_143_v0Wen;
    logic         io_diffCommits_info_143_vlWen;
    logic [5:0]   io_diffCommits_info_144_ldest;
    logic [7:0]   io_diffCommits_info_144_pdest;
    logic         io_diffCommits_info_144_rfWen;
    logic         io_diffCommits_info_144_fpWen;
    logic         io_diffCommits_info_144_vecWen;
    logic         io_diffCommits_info_144_v0Wen;
    logic         io_diffCommits_info_144_vlWen;
    logic [5:0]   io_diffCommits_info_145_ldest;
    logic [7:0]   io_diffCommits_info_145_pdest;
    logic         io_diffCommits_info_145_rfWen;
    logic         io_diffCommits_info_145_fpWen;
    logic         io_diffCommits_info_145_vecWen;
    logic         io_diffCommits_info_145_v0Wen;
    logic         io_diffCommits_info_145_vlWen;
    logic [5:0]   io_diffCommits_info_146_ldest;
    logic [7:0]   io_diffCommits_info_146_pdest;
    logic         io_diffCommits_info_146_rfWen;
    logic         io_diffCommits_info_146_fpWen;
    logic         io_diffCommits_info_146_vecWen;
    logic         io_diffCommits_info_146_v0Wen;
    logic         io_diffCommits_info_146_vlWen;
    logic [5:0]   io_diffCommits_info_147_ldest;
    logic [7:0]   io_diffCommits_info_147_pdest;
    logic         io_diffCommits_info_147_rfWen;
    logic         io_diffCommits_info_147_fpWen;
    logic         io_diffCommits_info_147_vecWen;
    logic         io_diffCommits_info_147_v0Wen;
    logic         io_diffCommits_info_147_vlWen;
    logic [5:0]   io_diffCommits_info_148_ldest;
    logic [7:0]   io_diffCommits_info_148_pdest;
    logic         io_diffCommits_info_148_rfWen;
    logic         io_diffCommits_info_148_fpWen;
    logic         io_diffCommits_info_148_vecWen;
    logic         io_diffCommits_info_148_v0Wen;
    logic         io_diffCommits_info_148_vlWen;
    logic [5:0]   io_diffCommits_info_149_ldest;
    logic [7:0]   io_diffCommits_info_149_pdest;
    logic         io_diffCommits_info_149_rfWen;
    logic         io_diffCommits_info_149_fpWen;
    logic         io_diffCommits_info_149_vecWen;
    logic         io_diffCommits_info_149_v0Wen;
    logic         io_diffCommits_info_149_vlWen;
    logic [5:0]   io_diffCommits_info_150_ldest;
    logic [7:0]   io_diffCommits_info_150_pdest;
    logic         io_diffCommits_info_150_rfWen;
    logic         io_diffCommits_info_150_fpWen;
    logic         io_diffCommits_info_150_vecWen;
    logic         io_diffCommits_info_150_v0Wen;
    logic         io_diffCommits_info_150_vlWen;
    logic [5:0]   io_diffCommits_info_151_ldest;
    logic [7:0]   io_diffCommits_info_151_pdest;
    logic         io_diffCommits_info_151_rfWen;
    logic         io_diffCommits_info_151_fpWen;
    logic         io_diffCommits_info_151_vecWen;
    logic         io_diffCommits_info_151_v0Wen;
    logic         io_diffCommits_info_151_vlWen;
    logic [5:0]   io_diffCommits_info_152_ldest;
    logic [7:0]   io_diffCommits_info_152_pdest;
    logic         io_diffCommits_info_152_rfWen;
    logic         io_diffCommits_info_152_fpWen;
    logic         io_diffCommits_info_152_vecWen;
    logic         io_diffCommits_info_152_v0Wen;
    logic         io_diffCommits_info_152_vlWen;
    logic [5:0]   io_diffCommits_info_153_ldest;
    logic [7:0]   io_diffCommits_info_153_pdest;
    logic         io_diffCommits_info_153_rfWen;
    logic         io_diffCommits_info_153_fpWen;
    logic         io_diffCommits_info_153_vecWen;
    logic         io_diffCommits_info_153_v0Wen;
    logic         io_diffCommits_info_153_vlWen;
    logic [5:0]   io_diffCommits_info_154_ldest;
    logic [7:0]   io_diffCommits_info_154_pdest;
    logic         io_diffCommits_info_154_rfWen;
    logic         io_diffCommits_info_154_fpWen;
    logic         io_diffCommits_info_154_vecWen;
    logic         io_diffCommits_info_154_v0Wen;
    logic         io_diffCommits_info_154_vlWen;
    logic [5:0]   io_diffCommits_info_155_ldest;
    logic [7:0]   io_diffCommits_info_155_pdest;
    logic         io_diffCommits_info_155_rfWen;
    logic         io_diffCommits_info_155_fpWen;
    logic         io_diffCommits_info_155_vecWen;
    logic         io_diffCommits_info_155_v0Wen;
    logic         io_diffCommits_info_155_vlWen;
    logic [5:0]   io_diffCommits_info_156_ldest;
    logic [7:0]   io_diffCommits_info_156_pdest;
    logic         io_diffCommits_info_156_rfWen;
    logic         io_diffCommits_info_156_fpWen;
    logic         io_diffCommits_info_156_vecWen;
    logic         io_diffCommits_info_156_v0Wen;
    logic         io_diffCommits_info_156_vlWen;
    logic [5:0]   io_diffCommits_info_157_ldest;
    logic [7:0]   io_diffCommits_info_157_pdest;
    logic         io_diffCommits_info_157_rfWen;
    logic         io_diffCommits_info_157_fpWen;
    logic         io_diffCommits_info_157_vecWen;
    logic         io_diffCommits_info_157_v0Wen;
    logic         io_diffCommits_info_157_vlWen;
    logic [5:0]   io_diffCommits_info_158_ldest;
    logic [7:0]   io_diffCommits_info_158_pdest;
    logic         io_diffCommits_info_158_rfWen;
    logic         io_diffCommits_info_158_fpWen;
    logic         io_diffCommits_info_158_vecWen;
    logic         io_diffCommits_info_158_v0Wen;
    logic         io_diffCommits_info_158_vlWen;
    logic [5:0]   io_diffCommits_info_159_ldest;
    logic [7:0]   io_diffCommits_info_159_pdest;
    logic         io_diffCommits_info_159_rfWen;
    logic         io_diffCommits_info_159_fpWen;
    logic         io_diffCommits_info_159_vecWen;
    logic         io_diffCommits_info_159_v0Wen;
    logic         io_diffCommits_info_159_vlWen;
    logic [5:0]   io_diffCommits_info_160_ldest;
    logic [7:0]   io_diffCommits_info_160_pdest;
    logic         io_diffCommits_info_160_rfWen;
    logic         io_diffCommits_info_160_fpWen;
    logic         io_diffCommits_info_160_vecWen;
    logic         io_diffCommits_info_160_v0Wen;
    logic         io_diffCommits_info_160_vlWen;
    logic [5:0]   io_diffCommits_info_161_ldest;
    logic [7:0]   io_diffCommits_info_161_pdest;
    logic         io_diffCommits_info_161_rfWen;
    logic         io_diffCommits_info_161_fpWen;
    logic         io_diffCommits_info_161_vecWen;
    logic         io_diffCommits_info_161_v0Wen;
    logic         io_diffCommits_info_161_vlWen;
    logic [5:0]   io_diffCommits_info_162_ldest;
    logic [7:0]   io_diffCommits_info_162_pdest;
    logic         io_diffCommits_info_162_rfWen;
    logic         io_diffCommits_info_162_fpWen;
    logic         io_diffCommits_info_162_vecWen;
    logic         io_diffCommits_info_162_v0Wen;
    logic         io_diffCommits_info_162_vlWen;
    logic [5:0]   io_diffCommits_info_163_ldest;
    logic [7:0]   io_diffCommits_info_163_pdest;
    logic         io_diffCommits_info_163_rfWen;
    logic         io_diffCommits_info_163_fpWen;
    logic         io_diffCommits_info_163_vecWen;
    logic         io_diffCommits_info_163_v0Wen;
    logic         io_diffCommits_info_163_vlWen;
    logic [5:0]   io_diffCommits_info_164_ldest;
    logic [7:0]   io_diffCommits_info_164_pdest;
    logic         io_diffCommits_info_164_rfWen;
    logic         io_diffCommits_info_164_fpWen;
    logic         io_diffCommits_info_164_vecWen;
    logic         io_diffCommits_info_164_v0Wen;
    logic         io_diffCommits_info_164_vlWen;
    logic [5:0]   io_diffCommits_info_165_ldest;
    logic [7:0]   io_diffCommits_info_165_pdest;
    logic         io_diffCommits_info_165_rfWen;
    logic         io_diffCommits_info_165_fpWen;
    logic         io_diffCommits_info_165_vecWen;
    logic         io_diffCommits_info_165_v0Wen;
    logic         io_diffCommits_info_165_vlWen;
    logic [5:0]   io_diffCommits_info_166_ldest;
    logic [7:0]   io_diffCommits_info_166_pdest;
    logic         io_diffCommits_info_166_rfWen;
    logic         io_diffCommits_info_166_fpWen;
    logic         io_diffCommits_info_166_vecWen;
    logic         io_diffCommits_info_166_v0Wen;
    logic         io_diffCommits_info_166_vlWen;
    logic [5:0]   io_diffCommits_info_167_ldest;
    logic [7:0]   io_diffCommits_info_167_pdest;
    logic         io_diffCommits_info_167_rfWen;
    logic         io_diffCommits_info_167_fpWen;
    logic         io_diffCommits_info_167_vecWen;
    logic         io_diffCommits_info_167_v0Wen;
    logic         io_diffCommits_info_167_vlWen;
    logic [5:0]   io_diffCommits_info_168_ldest;
    logic [7:0]   io_diffCommits_info_168_pdest;
    logic         io_diffCommits_info_168_rfWen;
    logic         io_diffCommits_info_168_fpWen;
    logic         io_diffCommits_info_168_vecWen;
    logic         io_diffCommits_info_168_v0Wen;
    logic         io_diffCommits_info_168_vlWen;
    logic [5:0]   io_diffCommits_info_169_ldest;
    logic [7:0]   io_diffCommits_info_169_pdest;
    logic         io_diffCommits_info_169_rfWen;
    logic         io_diffCommits_info_169_fpWen;
    logic         io_diffCommits_info_169_vecWen;
    logic         io_diffCommits_info_169_v0Wen;
    logic         io_diffCommits_info_169_vlWen;
    logic [5:0]   io_diffCommits_info_170_ldest;
    logic [7:0]   io_diffCommits_info_170_pdest;
    logic         io_diffCommits_info_170_rfWen;
    logic         io_diffCommits_info_170_fpWen;
    logic         io_diffCommits_info_170_vecWen;
    logic         io_diffCommits_info_170_v0Wen;
    logic         io_diffCommits_info_170_vlWen;
    logic [5:0]   io_diffCommits_info_171_ldest;
    logic [7:0]   io_diffCommits_info_171_pdest;
    logic         io_diffCommits_info_171_rfWen;
    logic         io_diffCommits_info_171_fpWen;
    logic         io_diffCommits_info_171_vecWen;
    logic         io_diffCommits_info_171_v0Wen;
    logic         io_diffCommits_info_171_vlWen;
    logic [5:0]   io_diffCommits_info_172_ldest;
    logic [7:0]   io_diffCommits_info_172_pdest;
    logic         io_diffCommits_info_172_rfWen;
    logic         io_diffCommits_info_172_fpWen;
    logic         io_diffCommits_info_172_vecWen;
    logic         io_diffCommits_info_172_v0Wen;
    logic         io_diffCommits_info_172_vlWen;
    logic [5:0]   io_diffCommits_info_173_ldest;
    logic [7:0]   io_diffCommits_info_173_pdest;
    logic         io_diffCommits_info_173_rfWen;
    logic         io_diffCommits_info_173_fpWen;
    logic         io_diffCommits_info_173_vecWen;
    logic         io_diffCommits_info_173_v0Wen;
    logic         io_diffCommits_info_173_vlWen;
    logic [5:0]   io_diffCommits_info_174_ldest;
    logic [7:0]   io_diffCommits_info_174_pdest;
    logic         io_diffCommits_info_174_rfWen;
    logic         io_diffCommits_info_174_fpWen;
    logic         io_diffCommits_info_174_vecWen;
    logic         io_diffCommits_info_174_v0Wen;
    logic         io_diffCommits_info_174_vlWen;
    logic [5:0]   io_diffCommits_info_175_ldest;
    logic [7:0]   io_diffCommits_info_175_pdest;
    logic         io_diffCommits_info_175_rfWen;
    logic         io_diffCommits_info_175_fpWen;
    logic         io_diffCommits_info_175_vecWen;
    logic         io_diffCommits_info_175_v0Wen;
    logic         io_diffCommits_info_175_vlWen;
    logic [5:0]   io_diffCommits_info_176_ldest;
    logic [7:0]   io_diffCommits_info_176_pdest;
    logic         io_diffCommits_info_176_rfWen;
    logic         io_diffCommits_info_176_fpWen;
    logic         io_diffCommits_info_176_vecWen;
    logic         io_diffCommits_info_176_v0Wen;
    logic         io_diffCommits_info_176_vlWen;
    logic [5:0]   io_diffCommits_info_177_ldest;
    logic [7:0]   io_diffCommits_info_177_pdest;
    logic         io_diffCommits_info_177_rfWen;
    logic         io_diffCommits_info_177_fpWen;
    logic         io_diffCommits_info_177_vecWen;
    logic         io_diffCommits_info_177_v0Wen;
    logic         io_diffCommits_info_177_vlWen;
    logic [5:0]   io_diffCommits_info_178_ldest;
    logic [7:0]   io_diffCommits_info_178_pdest;
    logic         io_diffCommits_info_178_rfWen;
    logic         io_diffCommits_info_178_fpWen;
    logic         io_diffCommits_info_178_vecWen;
    logic         io_diffCommits_info_178_v0Wen;
    logic         io_diffCommits_info_178_vlWen;
    logic [5:0]   io_diffCommits_info_179_ldest;
    logic [7:0]   io_diffCommits_info_179_pdest;
    logic         io_diffCommits_info_179_rfWen;
    logic         io_diffCommits_info_179_fpWen;
    logic         io_diffCommits_info_179_vecWen;
    logic         io_diffCommits_info_179_v0Wen;
    logic         io_diffCommits_info_179_vlWen;
    logic [5:0]   io_diffCommits_info_180_ldest;
    logic [7:0]   io_diffCommits_info_180_pdest;
    logic         io_diffCommits_info_180_rfWen;
    logic         io_diffCommits_info_180_fpWen;
    logic         io_diffCommits_info_180_vecWen;
    logic         io_diffCommits_info_180_v0Wen;
    logic         io_diffCommits_info_180_vlWen;
    logic [5:0]   io_diffCommits_info_181_ldest;
    logic [7:0]   io_diffCommits_info_181_pdest;
    logic         io_diffCommits_info_181_rfWen;
    logic         io_diffCommits_info_181_fpWen;
    logic         io_diffCommits_info_181_vecWen;
    logic         io_diffCommits_info_181_v0Wen;
    logic         io_diffCommits_info_181_vlWen;
    logic [5:0]   io_diffCommits_info_182_ldest;
    logic [7:0]   io_diffCommits_info_182_pdest;
    logic         io_diffCommits_info_182_rfWen;
    logic         io_diffCommits_info_182_fpWen;
    logic         io_diffCommits_info_182_vecWen;
    logic         io_diffCommits_info_182_v0Wen;
    logic         io_diffCommits_info_182_vlWen;
    logic [5:0]   io_diffCommits_info_183_ldest;
    logic [7:0]   io_diffCommits_info_183_pdest;
    logic         io_diffCommits_info_183_rfWen;
    logic         io_diffCommits_info_183_fpWen;
    logic         io_diffCommits_info_183_vecWen;
    logic         io_diffCommits_info_183_v0Wen;
    logic         io_diffCommits_info_183_vlWen;
    logic [5:0]   io_diffCommits_info_184_ldest;
    logic [7:0]   io_diffCommits_info_184_pdest;
    logic         io_diffCommits_info_184_rfWen;
    logic         io_diffCommits_info_184_fpWen;
    logic         io_diffCommits_info_184_vecWen;
    logic         io_diffCommits_info_184_v0Wen;
    logic         io_diffCommits_info_184_vlWen;
    logic [5:0]   io_diffCommits_info_185_ldest;
    logic [7:0]   io_diffCommits_info_185_pdest;
    logic         io_diffCommits_info_185_rfWen;
    logic         io_diffCommits_info_185_fpWen;
    logic         io_diffCommits_info_185_vecWen;
    logic         io_diffCommits_info_185_v0Wen;
    logic         io_diffCommits_info_185_vlWen;
    logic [5:0]   io_diffCommits_info_186_ldest;
    logic [7:0]   io_diffCommits_info_186_pdest;
    logic         io_diffCommits_info_186_rfWen;
    logic         io_diffCommits_info_186_fpWen;
    logic         io_diffCommits_info_186_vecWen;
    logic         io_diffCommits_info_186_v0Wen;
    logic         io_diffCommits_info_186_vlWen;
    logic [5:0]   io_diffCommits_info_187_ldest;
    logic [7:0]   io_diffCommits_info_187_pdest;
    logic         io_diffCommits_info_187_rfWen;
    logic         io_diffCommits_info_187_fpWen;
    logic         io_diffCommits_info_187_vecWen;
    logic         io_diffCommits_info_187_v0Wen;
    logic         io_diffCommits_info_187_vlWen;
    logic [5:0]   io_diffCommits_info_188_ldest;
    logic [7:0]   io_diffCommits_info_188_pdest;
    logic         io_diffCommits_info_188_rfWen;
    logic         io_diffCommits_info_188_fpWen;
    logic         io_diffCommits_info_188_vecWen;
    logic         io_diffCommits_info_188_v0Wen;
    logic         io_diffCommits_info_188_vlWen;
    logic [5:0]   io_diffCommits_info_189_ldest;
    logic [7:0]   io_diffCommits_info_189_pdest;
    logic         io_diffCommits_info_189_rfWen;
    logic         io_diffCommits_info_189_fpWen;
    logic         io_diffCommits_info_189_vecWen;
    logic         io_diffCommits_info_189_v0Wen;
    logic         io_diffCommits_info_189_vlWen;
    logic [5:0]   io_diffCommits_info_190_ldest;
    logic [7:0]   io_diffCommits_info_190_pdest;
    logic         io_diffCommits_info_190_rfWen;
    logic         io_diffCommits_info_190_fpWen;
    logic         io_diffCommits_info_190_vecWen;
    logic         io_diffCommits_info_190_v0Wen;
    logic         io_diffCommits_info_190_vlWen;
    logic [5:0]   io_diffCommits_info_191_ldest;
    logic [7:0]   io_diffCommits_info_191_pdest;
    logic         io_diffCommits_info_191_rfWen;
    logic         io_diffCommits_info_191_fpWen;
    logic         io_diffCommits_info_191_vecWen;
    logic         io_diffCommits_info_191_v0Wen;
    logic         io_diffCommits_info_191_vlWen;
    logic [5:0]   io_diffCommits_info_192_ldest;
    logic [7:0]   io_diffCommits_info_192_pdest;
    logic         io_diffCommits_info_192_rfWen;
    logic         io_diffCommits_info_192_fpWen;
    logic         io_diffCommits_info_192_vecWen;
    logic         io_diffCommits_info_192_v0Wen;
    logic         io_diffCommits_info_192_vlWen;
    logic [5:0]   io_diffCommits_info_193_ldest;
    logic [7:0]   io_diffCommits_info_193_pdest;
    logic         io_diffCommits_info_193_rfWen;
    logic         io_diffCommits_info_193_fpWen;
    logic         io_diffCommits_info_193_vecWen;
    logic         io_diffCommits_info_193_v0Wen;
    logic         io_diffCommits_info_193_vlWen;
    logic [5:0]   io_diffCommits_info_194_ldest;
    logic [7:0]   io_diffCommits_info_194_pdest;
    logic         io_diffCommits_info_194_rfWen;
    logic         io_diffCommits_info_194_fpWen;
    logic         io_diffCommits_info_194_vecWen;
    logic         io_diffCommits_info_194_v0Wen;
    logic         io_diffCommits_info_194_vlWen;
    logic [5:0]   io_diffCommits_info_195_ldest;
    logic [7:0]   io_diffCommits_info_195_pdest;
    logic         io_diffCommits_info_195_rfWen;
    logic         io_diffCommits_info_195_fpWen;
    logic         io_diffCommits_info_195_vecWen;
    logic         io_diffCommits_info_195_v0Wen;
    logic         io_diffCommits_info_195_vlWen;
    logic [5:0]   io_diffCommits_info_196_ldest;
    logic [7:0]   io_diffCommits_info_196_pdest;
    logic         io_diffCommits_info_196_rfWen;
    logic         io_diffCommits_info_196_fpWen;
    logic         io_diffCommits_info_196_vecWen;
    logic         io_diffCommits_info_196_v0Wen;
    logic         io_diffCommits_info_196_vlWen;
    logic [5:0]   io_diffCommits_info_197_ldest;
    logic [7:0]   io_diffCommits_info_197_pdest;
    logic         io_diffCommits_info_197_rfWen;
    logic         io_diffCommits_info_197_fpWen;
    logic         io_diffCommits_info_197_vecWen;
    logic         io_diffCommits_info_197_v0Wen;
    logic         io_diffCommits_info_197_vlWen;
    logic [5:0]   io_diffCommits_info_198_ldest;
    logic [7:0]   io_diffCommits_info_198_pdest;
    logic         io_diffCommits_info_198_rfWen;
    logic         io_diffCommits_info_198_fpWen;
    logic         io_diffCommits_info_198_vecWen;
    logic         io_diffCommits_info_198_v0Wen;
    logic         io_diffCommits_info_198_vlWen;
    logic [5:0]   io_diffCommits_info_199_ldest;
    logic [7:0]   io_diffCommits_info_199_pdest;
    logic         io_diffCommits_info_199_rfWen;
    logic         io_diffCommits_info_199_fpWen;
    logic         io_diffCommits_info_199_vecWen;
    logic         io_diffCommits_info_199_v0Wen;
    logic         io_diffCommits_info_199_vlWen;
    logic [5:0]   io_diffCommits_info_200_ldest;
    logic [7:0]   io_diffCommits_info_200_pdest;
    logic         io_diffCommits_info_200_rfWen;
    logic         io_diffCommits_info_200_fpWen;
    logic         io_diffCommits_info_200_vecWen;
    logic         io_diffCommits_info_200_v0Wen;
    logic         io_diffCommits_info_200_vlWen;
    logic [5:0]   io_diffCommits_info_201_ldest;
    logic [7:0]   io_diffCommits_info_201_pdest;
    logic         io_diffCommits_info_201_rfWen;
    logic         io_diffCommits_info_201_fpWen;
    logic         io_diffCommits_info_201_vecWen;
    logic         io_diffCommits_info_201_v0Wen;
    logic         io_diffCommits_info_201_vlWen;
    logic [5:0]   io_diffCommits_info_202_ldest;
    logic [7:0]   io_diffCommits_info_202_pdest;
    logic         io_diffCommits_info_202_rfWen;
    logic         io_diffCommits_info_202_fpWen;
    logic         io_diffCommits_info_202_vecWen;
    logic         io_diffCommits_info_202_v0Wen;
    logic         io_diffCommits_info_202_vlWen;
    logic [5:0]   io_diffCommits_info_203_ldest;
    logic [7:0]   io_diffCommits_info_203_pdest;
    logic         io_diffCommits_info_203_rfWen;
    logic         io_diffCommits_info_203_fpWen;
    logic         io_diffCommits_info_203_vecWen;
    logic         io_diffCommits_info_203_v0Wen;
    logic         io_diffCommits_info_203_vlWen;
    logic [5:0]   io_diffCommits_info_204_ldest;
    logic [7:0]   io_diffCommits_info_204_pdest;
    logic         io_diffCommits_info_204_rfWen;
    logic         io_diffCommits_info_204_fpWen;
    logic         io_diffCommits_info_204_vecWen;
    logic         io_diffCommits_info_204_v0Wen;
    logic         io_diffCommits_info_204_vlWen;
    logic [5:0]   io_diffCommits_info_205_ldest;
    logic [7:0]   io_diffCommits_info_205_pdest;
    logic         io_diffCommits_info_205_rfWen;
    logic         io_diffCommits_info_205_fpWen;
    logic         io_diffCommits_info_205_vecWen;
    logic         io_diffCommits_info_205_v0Wen;
    logic         io_diffCommits_info_205_vlWen;
    logic [5:0]   io_diffCommits_info_206_ldest;
    logic [7:0]   io_diffCommits_info_206_pdest;
    logic         io_diffCommits_info_206_rfWen;
    logic         io_diffCommits_info_206_fpWen;
    logic         io_diffCommits_info_206_vecWen;
    logic         io_diffCommits_info_206_v0Wen;
    logic         io_diffCommits_info_206_vlWen;
    logic [5:0]   io_diffCommits_info_207_ldest;
    logic [7:0]   io_diffCommits_info_207_pdest;
    logic         io_diffCommits_info_207_rfWen;
    logic         io_diffCommits_info_207_fpWen;
    logic         io_diffCommits_info_207_vecWen;
    logic         io_diffCommits_info_207_v0Wen;
    logic         io_diffCommits_info_207_vlWen;
    logic [5:0]   io_diffCommits_info_208_ldest;
    logic [7:0]   io_diffCommits_info_208_pdest;
    logic         io_diffCommits_info_208_rfWen;
    logic         io_diffCommits_info_208_fpWen;
    logic         io_diffCommits_info_208_vecWen;
    logic         io_diffCommits_info_208_v0Wen;
    logic         io_diffCommits_info_208_vlWen;
    logic [5:0]   io_diffCommits_info_209_ldest;
    logic [7:0]   io_diffCommits_info_209_pdest;
    logic         io_diffCommits_info_209_rfWen;
    logic         io_diffCommits_info_209_fpWen;
    logic         io_diffCommits_info_209_vecWen;
    logic         io_diffCommits_info_209_v0Wen;
    logic         io_diffCommits_info_209_vlWen;
    logic [5:0]   io_diffCommits_info_210_ldest;
    logic [7:0]   io_diffCommits_info_210_pdest;
    logic         io_diffCommits_info_210_rfWen;
    logic         io_diffCommits_info_210_fpWen;
    logic         io_diffCommits_info_210_vecWen;
    logic         io_diffCommits_info_210_v0Wen;
    logic         io_diffCommits_info_210_vlWen;
    logic [5:0]   io_diffCommits_info_211_ldest;
    logic [7:0]   io_diffCommits_info_211_pdest;
    logic         io_diffCommits_info_211_rfWen;
    logic         io_diffCommits_info_211_fpWen;
    logic         io_diffCommits_info_211_vecWen;
    logic         io_diffCommits_info_211_v0Wen;
    logic         io_diffCommits_info_211_vlWen;
    logic [5:0]   io_diffCommits_info_212_ldest;
    logic [7:0]   io_diffCommits_info_212_pdest;
    logic         io_diffCommits_info_212_rfWen;
    logic         io_diffCommits_info_212_fpWen;
    logic         io_diffCommits_info_212_vecWen;
    logic         io_diffCommits_info_212_v0Wen;
    logic         io_diffCommits_info_212_vlWen;
    logic [5:0]   io_diffCommits_info_213_ldest;
    logic [7:0]   io_diffCommits_info_213_pdest;
    logic         io_diffCommits_info_213_rfWen;
    logic         io_diffCommits_info_213_fpWen;
    logic         io_diffCommits_info_213_vecWen;
    logic         io_diffCommits_info_213_v0Wen;
    logic         io_diffCommits_info_213_vlWen;
    logic [5:0]   io_diffCommits_info_214_ldest;
    logic [7:0]   io_diffCommits_info_214_pdest;
    logic         io_diffCommits_info_214_rfWen;
    logic         io_diffCommits_info_214_fpWen;
    logic         io_diffCommits_info_214_vecWen;
    logic         io_diffCommits_info_214_v0Wen;
    logic         io_diffCommits_info_214_vlWen;
    logic [5:0]   io_diffCommits_info_215_ldest;
    logic [7:0]   io_diffCommits_info_215_pdest;
    logic         io_diffCommits_info_215_rfWen;
    logic         io_diffCommits_info_215_fpWen;
    logic         io_diffCommits_info_215_vecWen;
    logic         io_diffCommits_info_215_v0Wen;
    logic         io_diffCommits_info_215_vlWen;
    logic [5:0]   io_diffCommits_info_216_ldest;
    logic [7:0]   io_diffCommits_info_216_pdest;
    logic         io_diffCommits_info_216_rfWen;
    logic         io_diffCommits_info_216_fpWen;
    logic         io_diffCommits_info_216_vecWen;
    logic         io_diffCommits_info_216_v0Wen;
    logic         io_diffCommits_info_216_vlWen;
    logic [5:0]   io_diffCommits_info_217_ldest;
    logic [7:0]   io_diffCommits_info_217_pdest;
    logic         io_diffCommits_info_217_rfWen;
    logic         io_diffCommits_info_217_fpWen;
    logic         io_diffCommits_info_217_vecWen;
    logic         io_diffCommits_info_217_v0Wen;
    logic         io_diffCommits_info_217_vlWen;
    logic [5:0]   io_diffCommits_info_218_ldest;
    logic [7:0]   io_diffCommits_info_218_pdest;
    logic         io_diffCommits_info_218_rfWen;
    logic         io_diffCommits_info_218_fpWen;
    logic         io_diffCommits_info_218_vecWen;
    logic         io_diffCommits_info_218_v0Wen;
    logic         io_diffCommits_info_218_vlWen;
    logic [5:0]   io_diffCommits_info_219_ldest;
    logic [7:0]   io_diffCommits_info_219_pdest;
    logic         io_diffCommits_info_219_rfWen;
    logic         io_diffCommits_info_219_fpWen;
    logic         io_diffCommits_info_219_vecWen;
    logic         io_diffCommits_info_219_v0Wen;
    logic         io_diffCommits_info_219_vlWen;
    logic [5:0]   io_diffCommits_info_220_ldest;
    logic [7:0]   io_diffCommits_info_220_pdest;
    logic         io_diffCommits_info_220_rfWen;
    logic         io_diffCommits_info_220_fpWen;
    logic         io_diffCommits_info_220_vecWen;
    logic         io_diffCommits_info_220_v0Wen;
    logic         io_diffCommits_info_220_vlWen;
    logic [5:0]   io_diffCommits_info_221_ldest;
    logic [7:0]   io_diffCommits_info_221_pdest;
    logic         io_diffCommits_info_221_rfWen;
    logic         io_diffCommits_info_221_fpWen;
    logic         io_diffCommits_info_221_vecWen;
    logic         io_diffCommits_info_221_v0Wen;
    logic         io_diffCommits_info_221_vlWen;
    logic [5:0]   io_diffCommits_info_222_ldest;
    logic [7:0]   io_diffCommits_info_222_pdest;
    logic         io_diffCommits_info_222_rfWen;
    logic         io_diffCommits_info_222_fpWen;
    logic         io_diffCommits_info_222_vecWen;
    logic         io_diffCommits_info_222_v0Wen;
    logic         io_diffCommits_info_222_vlWen;
    logic [5:0]   io_diffCommits_info_223_ldest;
    logic [7:0]   io_diffCommits_info_223_pdest;
    logic         io_diffCommits_info_223_rfWen;
    logic         io_diffCommits_info_223_fpWen;
    logic         io_diffCommits_info_223_vecWen;
    logic         io_diffCommits_info_223_v0Wen;
    logic         io_diffCommits_info_223_vlWen;
    logic [5:0]   io_diffCommits_info_224_ldest;
    logic [7:0]   io_diffCommits_info_224_pdest;
    logic         io_diffCommits_info_224_rfWen;
    logic         io_diffCommits_info_224_fpWen;
    logic         io_diffCommits_info_224_vecWen;
    logic         io_diffCommits_info_224_v0Wen;
    logic         io_diffCommits_info_224_vlWen;
    logic [5:0]   io_diffCommits_info_225_ldest;
    logic [7:0]   io_diffCommits_info_225_pdest;
    logic         io_diffCommits_info_225_rfWen;
    logic         io_diffCommits_info_225_fpWen;
    logic         io_diffCommits_info_225_vecWen;
    logic         io_diffCommits_info_225_v0Wen;
    logic         io_diffCommits_info_225_vlWen;
    logic [5:0]   io_diffCommits_info_226_ldest;
    logic [7:0]   io_diffCommits_info_226_pdest;
    logic         io_diffCommits_info_226_rfWen;
    logic         io_diffCommits_info_226_fpWen;
    logic         io_diffCommits_info_226_vecWen;
    logic         io_diffCommits_info_226_v0Wen;
    logic         io_diffCommits_info_226_vlWen;
    logic [5:0]   io_diffCommits_info_227_ldest;
    logic [7:0]   io_diffCommits_info_227_pdest;
    logic         io_diffCommits_info_227_rfWen;
    logic         io_diffCommits_info_227_fpWen;
    logic         io_diffCommits_info_227_vecWen;
    logic         io_diffCommits_info_227_v0Wen;
    logic         io_diffCommits_info_227_vlWen;
    logic [5:0]   io_diffCommits_info_228_ldest;
    logic [7:0]   io_diffCommits_info_228_pdest;
    logic         io_diffCommits_info_228_rfWen;
    logic         io_diffCommits_info_228_fpWen;
    logic         io_diffCommits_info_228_vecWen;
    logic         io_diffCommits_info_228_v0Wen;
    logic         io_diffCommits_info_228_vlWen;
    logic [5:0]   io_diffCommits_info_229_ldest;
    logic [7:0]   io_diffCommits_info_229_pdest;
    logic         io_diffCommits_info_229_rfWen;
    logic         io_diffCommits_info_229_fpWen;
    logic         io_diffCommits_info_229_vecWen;
    logic         io_diffCommits_info_229_v0Wen;
    logic         io_diffCommits_info_229_vlWen;
    logic [5:0]   io_diffCommits_info_230_ldest;
    logic [7:0]   io_diffCommits_info_230_pdest;
    logic         io_diffCommits_info_230_rfWen;
    logic         io_diffCommits_info_230_fpWen;
    logic         io_diffCommits_info_230_vecWen;
    logic         io_diffCommits_info_230_v0Wen;
    logic         io_diffCommits_info_230_vlWen;
    logic [5:0]   io_diffCommits_info_231_ldest;
    logic [7:0]   io_diffCommits_info_231_pdest;
    logic         io_diffCommits_info_231_rfWen;
    logic         io_diffCommits_info_231_fpWen;
    logic         io_diffCommits_info_231_vecWen;
    logic         io_diffCommits_info_231_v0Wen;
    logic         io_diffCommits_info_231_vlWen;
    logic [5:0]   io_diffCommits_info_232_ldest;
    logic [7:0]   io_diffCommits_info_232_pdest;
    logic         io_diffCommits_info_232_rfWen;
    logic         io_diffCommits_info_232_fpWen;
    logic         io_diffCommits_info_232_vecWen;
    logic         io_diffCommits_info_232_v0Wen;
    logic         io_diffCommits_info_232_vlWen;
    logic [5:0]   io_diffCommits_info_233_ldest;
    logic [7:0]   io_diffCommits_info_233_pdest;
    logic         io_diffCommits_info_233_rfWen;
    logic         io_diffCommits_info_233_fpWen;
    logic         io_diffCommits_info_233_vecWen;
    logic         io_diffCommits_info_233_v0Wen;
    logic         io_diffCommits_info_233_vlWen;
    logic [5:0]   io_diffCommits_info_234_ldest;
    logic [7:0]   io_diffCommits_info_234_pdest;
    logic         io_diffCommits_info_234_rfWen;
    logic         io_diffCommits_info_234_fpWen;
    logic         io_diffCommits_info_234_vecWen;
    logic         io_diffCommits_info_234_v0Wen;
    logic         io_diffCommits_info_234_vlWen;
    logic [5:0]   io_diffCommits_info_235_ldest;
    logic [7:0]   io_diffCommits_info_235_pdest;
    logic         io_diffCommits_info_235_rfWen;
    logic         io_diffCommits_info_235_fpWen;
    logic         io_diffCommits_info_235_vecWen;
    logic         io_diffCommits_info_235_v0Wen;
    logic         io_diffCommits_info_235_vlWen;
    logic [5:0]   io_diffCommits_info_236_ldest;
    logic [7:0]   io_diffCommits_info_236_pdest;
    logic         io_diffCommits_info_236_rfWen;
    logic         io_diffCommits_info_236_fpWen;
    logic         io_diffCommits_info_236_vecWen;
    logic         io_diffCommits_info_236_v0Wen;
    logic         io_diffCommits_info_236_vlWen;
    logic [5:0]   io_diffCommits_info_237_ldest;
    logic [7:0]   io_diffCommits_info_237_pdest;
    logic         io_diffCommits_info_237_rfWen;
    logic         io_diffCommits_info_237_fpWen;
    logic         io_diffCommits_info_237_vecWen;
    logic         io_diffCommits_info_237_v0Wen;
    logic         io_diffCommits_info_237_vlWen;
    logic [5:0]   io_diffCommits_info_238_ldest;
    logic [7:0]   io_diffCommits_info_238_pdest;
    logic         io_diffCommits_info_238_rfWen;
    logic         io_diffCommits_info_238_fpWen;
    logic         io_diffCommits_info_238_vecWen;
    logic         io_diffCommits_info_238_v0Wen;
    logic         io_diffCommits_info_238_vlWen;
    logic [5:0]   io_diffCommits_info_239_ldest;
    logic [7:0]   io_diffCommits_info_239_pdest;
    logic         io_diffCommits_info_239_rfWen;
    logic         io_diffCommits_info_239_fpWen;
    logic         io_diffCommits_info_239_vecWen;
    logic         io_diffCommits_info_239_v0Wen;
    logic         io_diffCommits_info_239_vlWen;
    logic [5:0]   io_diffCommits_info_240_ldest;
    logic [7:0]   io_diffCommits_info_240_pdest;
    logic         io_diffCommits_info_240_rfWen;
    logic         io_diffCommits_info_240_fpWen;
    logic         io_diffCommits_info_240_vecWen;
    logic         io_diffCommits_info_240_v0Wen;
    logic         io_diffCommits_info_240_vlWen;
    logic [5:0]   io_diffCommits_info_241_ldest;
    logic [7:0]   io_diffCommits_info_241_pdest;
    logic         io_diffCommits_info_241_rfWen;
    logic         io_diffCommits_info_241_fpWen;
    logic         io_diffCommits_info_241_vecWen;
    logic         io_diffCommits_info_241_v0Wen;
    logic         io_diffCommits_info_241_vlWen;
    logic [5:0]   io_diffCommits_info_242_ldest;
    logic [7:0]   io_diffCommits_info_242_pdest;
    logic         io_diffCommits_info_242_rfWen;
    logic         io_diffCommits_info_242_fpWen;
    logic         io_diffCommits_info_242_vecWen;
    logic         io_diffCommits_info_242_v0Wen;
    logic         io_diffCommits_info_242_vlWen;
    logic [5:0]   io_diffCommits_info_243_ldest;
    logic [7:0]   io_diffCommits_info_243_pdest;
    logic         io_diffCommits_info_243_rfWen;
    logic         io_diffCommits_info_243_fpWen;
    logic         io_diffCommits_info_243_vecWen;
    logic         io_diffCommits_info_243_v0Wen;
    logic         io_diffCommits_info_243_vlWen;
    logic [5:0]   io_diffCommits_info_244_ldest;
    logic [7:0]   io_diffCommits_info_244_pdest;
    logic         io_diffCommits_info_244_rfWen;
    logic         io_diffCommits_info_244_fpWen;
    logic         io_diffCommits_info_244_vecWen;
    logic         io_diffCommits_info_244_v0Wen;
    logic         io_diffCommits_info_244_vlWen;
    logic [5:0]   io_diffCommits_info_245_ldest;
    logic [7:0]   io_diffCommits_info_245_pdest;
    logic         io_diffCommits_info_245_rfWen;
    logic         io_diffCommits_info_245_fpWen;
    logic         io_diffCommits_info_245_vecWen;
    logic         io_diffCommits_info_245_v0Wen;
    logic         io_diffCommits_info_245_vlWen;
    logic [5:0]   io_diffCommits_info_246_ldest;
    logic [7:0]   io_diffCommits_info_246_pdest;
    logic         io_diffCommits_info_246_rfWen;
    logic         io_diffCommits_info_246_fpWen;
    logic         io_diffCommits_info_246_vecWen;
    logic         io_diffCommits_info_246_v0Wen;
    logic         io_diffCommits_info_246_vlWen;
    logic [5:0]   io_diffCommits_info_247_ldest;
    logic [7:0]   io_diffCommits_info_247_pdest;
    logic         io_diffCommits_info_247_rfWen;
    logic         io_diffCommits_info_247_fpWen;
    logic         io_diffCommits_info_247_vecWen;
    logic         io_diffCommits_info_247_v0Wen;
    logic         io_diffCommits_info_247_vlWen;
    logic [5:0]   io_diffCommits_info_248_ldest;
    logic [7:0]   io_diffCommits_info_248_pdest;
    logic         io_diffCommits_info_248_rfWen;
    logic         io_diffCommits_info_248_fpWen;
    logic         io_diffCommits_info_248_vecWen;
    logic         io_diffCommits_info_248_v0Wen;
    logic         io_diffCommits_info_248_vlWen;
    logic [5:0]   io_diffCommits_info_249_ldest;
    logic [7:0]   io_diffCommits_info_249_pdest;
    logic         io_diffCommits_info_249_rfWen;
    logic         io_diffCommits_info_249_fpWen;
    logic         io_diffCommits_info_249_vecWen;
    logic         io_diffCommits_info_249_v0Wen;
    logic         io_diffCommits_info_249_vlWen;
    logic [5:0]   io_diffCommits_info_250_ldest;
    logic [7:0]   io_diffCommits_info_250_pdest;
    logic         io_diffCommits_info_250_rfWen;
    logic         io_diffCommits_info_250_fpWen;
    logic         io_diffCommits_info_250_vecWen;
    logic         io_diffCommits_info_250_v0Wen;
    logic         io_diffCommits_info_250_vlWen;
    logic [5:0]   io_diffCommits_info_251_ldest;
    logic [7:0]   io_diffCommits_info_251_pdest;
    logic         io_diffCommits_info_251_rfWen;
    logic         io_diffCommits_info_251_fpWen;
    logic         io_diffCommits_info_251_vecWen;
    logic         io_diffCommits_info_251_v0Wen;
    logic         io_diffCommits_info_251_vlWen;
    logic [5:0]   io_diffCommits_info_252_ldest;
    logic [7:0]   io_diffCommits_info_252_pdest;
    logic         io_diffCommits_info_252_rfWen;
    logic         io_diffCommits_info_252_fpWen;
    logic         io_diffCommits_info_252_vecWen;
    logic         io_diffCommits_info_252_v0Wen;
    logic         io_diffCommits_info_252_vlWen;
    logic [5:0]   io_diffCommits_info_253_ldest;
    logic [7:0]   io_diffCommits_info_253_pdest;
    logic         io_diffCommits_info_253_rfWen;
    logic         io_diffCommits_info_253_fpWen;
    logic         io_diffCommits_info_253_vecWen;
    logic         io_diffCommits_info_253_v0Wen;
    logic         io_diffCommits_info_253_vlWen;
    logic [5:0]   io_diffCommits_info_254_ldest;
    logic [7:0]   io_diffCommits_info_254_pdest;
    logic         io_diffCommits_info_254_rfWen;
    logic         io_diffCommits_info_254_fpWen;
    logic         io_diffCommits_info_254_vecWen;
    logic         io_diffCommits_info_254_v0Wen;
    logic         io_diffCommits_info_254_vlWen;
    logic [5:0]   io_diffCommits_info_255_ldest;
    logic [7:0]   io_diffCommits_info_255_pdest;
    logic [5:0]   io_diffCommits_info_256_ldest;
    logic [7:0]   io_diffCommits_info_256_pdest;
    logic [5:0]   io_diffCommits_info_257_ldest;
    logic [7:0]   io_diffCommits_info_257_pdest;
    logic [5:0]   io_diffCommits_info_258_ldest;
    logic [7:0]   io_diffCommits_info_258_pdest;
    logic [5:0]   io_diffCommits_info_259_ldest;
    logic [7:0]   io_diffCommits_info_259_pdest;
    logic [5:0]   io_diffCommits_info_260_ldest;
    logic [7:0]   io_diffCommits_info_260_pdest;
    logic [5:0]   io_diffCommits_info_261_ldest;
    logic [7:0]   io_diffCommits_info_261_pdest;
    logic [5:0]   io_diffCommits_info_262_ldest;
    logic [7:0]   io_diffCommits_info_262_pdest;
    logic [5:0]   io_diffCommits_info_263_ldest;
    logic [7:0]   io_diffCommits_info_263_pdest;
    logic [5:0]   io_diffCommits_info_264_ldest;
    logic [7:0]   io_diffCommits_info_264_pdest;
    logic [5:0]   io_diffCommits_info_265_ldest;
    logic [7:0]   io_diffCommits_info_265_pdest;
    logic [5:0]   io_diffCommits_info_266_ldest;
    logic [7:0]   io_diffCommits_info_266_pdest;
    logic [5:0]   io_diffCommits_info_267_ldest;
    logic [7:0]   io_diffCommits_info_267_pdest;
    logic [5:0]   io_diffCommits_info_268_ldest;
    logic [7:0]   io_diffCommits_info_268_pdest;
    logic [5:0]   io_diffCommits_info_269_ldest;
    logic [7:0]   io_diffCommits_info_269_pdest;
    logic [5:0]   io_diffCommits_info_270_ldest;
    logic [7:0]   io_diffCommits_info_270_pdest;
    logic [5:0]   io_diffCommits_info_271_ldest;
    logic [7:0]   io_diffCommits_info_271_pdest;
    logic [5:0]   io_diffCommits_info_272_ldest;
    logic [7:0]   io_diffCommits_info_272_pdest;
    logic [5:0]   io_diffCommits_info_273_ldest;
    logic [7:0]   io_diffCommits_info_273_pdest;
    logic [5:0]   io_diffCommits_info_274_ldest;
    logic [7:0]   io_diffCommits_info_274_pdest;
    logic [5:0]   io_diffCommits_info_275_ldest;
    logic [7:0]   io_diffCommits_info_275_pdest;
    logic [5:0]   io_diffCommits_info_276_ldest;
    logic [7:0]   io_diffCommits_info_276_pdest;
    logic [5:0]   io_diffCommits_info_277_ldest;
    logic [7:0]   io_diffCommits_info_277_pdest;
    logic [5:0]   io_diffCommits_info_278_ldest;
    logic [7:0]   io_diffCommits_info_278_pdest;
    logic [5:0]   io_diffCommits_info_279_ldest;
    logic [7:0]   io_diffCommits_info_279_pdest;
    logic [5:0]   io_diffCommits_info_280_ldest;
    logic [7:0]   io_diffCommits_info_280_pdest;
    logic [5:0]   io_diffCommits_info_281_ldest;
    logic [7:0]   io_diffCommits_info_281_pdest;
    logic [5:0]   io_diffCommits_info_282_ldest;
    logic [7:0]   io_diffCommits_info_282_pdest;
    logic [5:0]   io_diffCommits_info_283_ldest;
    logic [7:0]   io_diffCommits_info_283_pdest;
    logic [5:0]   io_diffCommits_info_284_ldest;
    logic [7:0]   io_diffCommits_info_284_pdest;
    logic [5:0]   io_diffCommits_info_285_ldest;
    logic [7:0]   io_diffCommits_info_285_pdest;
    logic [5:0]   io_diffCommits_info_286_ldest;
    logic [7:0]   io_diffCommits_info_286_pdest;
    logic [5:0]   io_diffCommits_info_287_ldest;
    logic [7:0]   io_diffCommits_info_287_pdest;
    logic [5:0]   io_diffCommits_info_288_ldest;
    logic [7:0]   io_diffCommits_info_288_pdest;
    logic [5:0]   io_diffCommits_info_289_ldest;
    logic [7:0]   io_diffCommits_info_289_pdest;
    logic [5:0]   io_diffCommits_info_290_ldest;
    logic [7:0]   io_diffCommits_info_290_pdest;
    logic [5:0]   io_diffCommits_info_291_ldest;
    logic [7:0]   io_diffCommits_info_291_pdest;
    logic [5:0]   io_diffCommits_info_292_ldest;
    logic [7:0]   io_diffCommits_info_292_pdest;
    logic [5:0]   io_diffCommits_info_293_ldest;
    logic [7:0]   io_diffCommits_info_293_pdest;
    logic [5:0]   io_diffCommits_info_294_ldest;
    logic [7:0]   io_diffCommits_info_294_pdest;
    logic [5:0]   io_diffCommits_info_295_ldest;
    logic [7:0]   io_diffCommits_info_295_pdest;
    logic [5:0]   io_diffCommits_info_296_ldest;
    logic [7:0]   io_diffCommits_info_296_pdest;
    logic [5:0]   io_diffCommits_info_297_ldest;
    logic [7:0]   io_diffCommits_info_297_pdest;
    logic [5:0]   io_diffCommits_info_298_ldest;
    logic [7:0]   io_diffCommits_info_298_pdest;
    logic [5:0]   io_diffCommits_info_299_ldest;
    logic [7:0]   io_diffCommits_info_299_pdest;
    logic [5:0]   io_diffCommits_info_300_ldest;
    logic [7:0]   io_diffCommits_info_300_pdest;
    logic [5:0]   io_diffCommits_info_301_ldest;
    logic [7:0]   io_diffCommits_info_301_pdest;
    logic [5:0]   io_diffCommits_info_302_ldest;
    logic [7:0]   io_diffCommits_info_302_pdest;
    logic [5:0]   io_diffCommits_info_303_ldest;
    logic [7:0]   io_diffCommits_info_303_pdest;
    logic [5:0]   io_diffCommits_info_304_ldest;
    logic [7:0]   io_diffCommits_info_304_pdest;
    logic [5:0]   io_diffCommits_info_305_ldest;
    logic [7:0]   io_diffCommits_info_305_pdest;
    logic [5:0]   io_diffCommits_info_306_ldest;
    logic [7:0]   io_diffCommits_info_306_pdest;
    logic [5:0]   io_diffCommits_info_307_ldest;
    logic [7:0]   io_diffCommits_info_307_pdest;
    logic [5:0]   io_diffCommits_info_308_ldest;
    logic [7:0]   io_diffCommits_info_308_pdest;
    logic [5:0]   io_diffCommits_info_309_ldest;
    logic [7:0]   io_diffCommits_info_309_pdest;
    logic [5:0]   io_diffCommits_info_310_ldest;
    logic [7:0]   io_diffCommits_info_310_pdest;
    logic [5:0]   io_diffCommits_info_311_ldest;
    logic [7:0]   io_diffCommits_info_311_pdest;
    logic [5:0]   io_diffCommits_info_312_ldest;
    logic [7:0]   io_diffCommits_info_312_pdest;
    logic [5:0]   io_diffCommits_info_313_ldest;
    logic [7:0]   io_diffCommits_info_313_pdest;
    logic [5:0]   io_diffCommits_info_314_ldest;
    logic [7:0]   io_diffCommits_info_314_pdest;
    logic [5:0]   io_diffCommits_info_315_ldest;
    logic [7:0]   io_diffCommits_info_315_pdest;
    logic [5:0]   io_diffCommits_info_316_ldest;
    logic [7:0]   io_diffCommits_info_316_pdest;
    logic [5:0]   io_diffCommits_info_317_ldest;
    logic [7:0]   io_diffCommits_info_317_pdest;
    logic [5:0]   io_diffCommits_info_318_ldest;
    logic [7:0]   io_diffCommits_info_318_pdest;
    logic [5:0]   io_diffCommits_info_319_ldest;
    logic [7:0]   io_diffCommits_info_319_pdest;
    logic [5:0]   io_diffCommits_info_320_ldest;
    logic [7:0]   io_diffCommits_info_320_pdest;
    logic [5:0]   io_diffCommits_info_321_ldest;
    logic [7:0]   io_diffCommits_info_321_pdest;
    logic [5:0]   io_diffCommits_info_322_ldest;
    logic [7:0]   io_diffCommits_info_322_pdest;
    logic [5:0]   io_diffCommits_info_323_ldest;
    logic [7:0]   io_diffCommits_info_323_pdest;
    logic [5:0]   io_diffCommits_info_324_ldest;
    logic [7:0]   io_diffCommits_info_324_pdest;
    logic [5:0]   io_diffCommits_info_325_ldest;
    logic [7:0]   io_diffCommits_info_325_pdest;
    logic [5:0]   io_diffCommits_info_326_ldest;
    logic [7:0]   io_diffCommits_info_326_pdest;
    logic [5:0]   io_diffCommits_info_327_ldest;
    logic [7:0]   io_diffCommits_info_327_pdest;
    logic [5:0]   io_diffCommits_info_328_ldest;
    logic [7:0]   io_diffCommits_info_328_pdest;
    logic [5:0]   io_diffCommits_info_329_ldest;
    logic [7:0]   io_diffCommits_info_329_pdest;
    logic [5:0]   io_diffCommits_info_330_ldest;
    logic [7:0]   io_diffCommits_info_330_pdest;
    logic [5:0]   io_diffCommits_info_331_ldest;
    logic [7:0]   io_diffCommits_info_331_pdest;
    logic [5:0]   io_diffCommits_info_332_ldest;
    logic [7:0]   io_diffCommits_info_332_pdest;
    logic [5:0]   io_diffCommits_info_333_ldest;
    logic [7:0]   io_diffCommits_info_333_pdest;
    logic [5:0]   io_diffCommits_info_334_ldest;
    logic [7:0]   io_diffCommits_info_334_pdest;
    logic [5:0]   io_diffCommits_info_335_ldest;
    logic [7:0]   io_diffCommits_info_335_pdest;
    logic [5:0]   io_diffCommits_info_336_ldest;
    logic [7:0]   io_diffCommits_info_336_pdest;
    logic [5:0]   io_diffCommits_info_337_ldest;
    logic [7:0]   io_diffCommits_info_337_pdest;
    logic [5:0]   io_diffCommits_info_338_ldest;
    logic [7:0]   io_diffCommits_info_338_pdest;
    logic [5:0]   io_diffCommits_info_339_ldest;
    logic [7:0]   io_diffCommits_info_339_pdest;
    logic [5:0]   io_diffCommits_info_340_ldest;
    logic [7:0]   io_diffCommits_info_340_pdest;
    logic [5:0]   io_diffCommits_info_341_ldest;
    logic [7:0]   io_diffCommits_info_341_pdest;
    logic [5:0]   io_diffCommits_info_342_ldest;
    logic [7:0]   io_diffCommits_info_342_pdest;
    logic [5:0]   io_diffCommits_info_343_ldest;
    logic [7:0]   io_diffCommits_info_343_pdest;
    logic [5:0]   io_diffCommits_info_344_ldest;
    logic [7:0]   io_diffCommits_info_344_pdest;
    logic [5:0]   io_diffCommits_info_345_ldest;
    logic [7:0]   io_diffCommits_info_345_pdest;
    logic [5:0]   io_diffCommits_info_346_ldest;
    logic [7:0]   io_diffCommits_info_346_pdest;
    logic [5:0]   io_diffCommits_info_347_ldest;
    logic [7:0]   io_diffCommits_info_347_pdest;
    logic [5:0]   io_diffCommits_info_348_ldest;
    logic [7:0]   io_diffCommits_info_348_pdest;
    logic [5:0]   io_diffCommits_info_349_ldest;
    logic [7:0]   io_diffCommits_info_349_pdest;
    logic [5:0]   io_diffCommits_info_350_ldest;
    logic [7:0]   io_diffCommits_info_350_pdest;
    logic [5:0]   io_diffCommits_info_351_ldest;
    logic [7:0]   io_diffCommits_info_351_pdest;
    logic [5:0]   io_diffCommits_info_352_ldest;
    logic [7:0]   io_diffCommits_info_352_pdest;
    logic [5:0]   io_diffCommits_info_353_ldest;
    logic [7:0]   io_diffCommits_info_353_pdest;
    logic [5:0]   io_diffCommits_info_354_ldest;
    logic [7:0]   io_diffCommits_info_354_pdest;
    logic [5:0]   io_diffCommits_info_355_ldest;
    logic [7:0]   io_diffCommits_info_355_pdest;
    logic [5:0]   io_diffCommits_info_356_ldest;
    logic [7:0]   io_diffCommits_info_356_pdest;
    logic [5:0]   io_diffCommits_info_357_ldest;
    logic [7:0]   io_diffCommits_info_357_pdest;
    logic [5:0]   io_diffCommits_info_358_ldest;
    logic [7:0]   io_diffCommits_info_358_pdest;
    logic [5:0]   io_diffCommits_info_359_ldest;
    logic [7:0]   io_diffCommits_info_359_pdest;
    logic [5:0]   io_diffCommits_info_360_ldest;
    logic [7:0]   io_diffCommits_info_360_pdest;
    logic [5:0]   io_diffCommits_info_361_ldest;
    logic [7:0]   io_diffCommits_info_361_pdest;
    logic [5:0]   io_diffCommits_info_362_ldest;
    logic [7:0]   io_diffCommits_info_362_pdest;
    logic [5:0]   io_diffCommits_info_363_ldest;
    logic [7:0]   io_diffCommits_info_363_pdest;
    logic [5:0]   io_diffCommits_info_364_ldest;
    logic [7:0]   io_diffCommits_info_364_pdest;
    logic [5:0]   io_diffCommits_info_365_ldest;
    logic [7:0]   io_diffCommits_info_365_pdest;
    logic [5:0]   io_diffCommits_info_366_ldest;
    logic [7:0]   io_diffCommits_info_366_pdest;
    logic [5:0]   io_diffCommits_info_367_ldest;
    logic [7:0]   io_diffCommits_info_367_pdest;
    logic [5:0]   io_diffCommits_info_368_ldest;
    logic [7:0]   io_diffCommits_info_368_pdest;
    logic [5:0]   io_diffCommits_info_369_ldest;
    logic [7:0]   io_diffCommits_info_369_pdest;
    logic [5:0]   io_diffCommits_info_370_ldest;
    logic [7:0]   io_diffCommits_info_370_pdest;
    logic [5:0]   io_diffCommits_info_371_ldest;
    logic [7:0]   io_diffCommits_info_371_pdest;
    logic [5:0]   io_diffCommits_info_372_ldest;
    logic [7:0]   io_diffCommits_info_372_pdest;
    logic [5:0]   io_diffCommits_info_373_ldest;
    logic [7:0]   io_diffCommits_info_373_pdest;
    logic [5:0]   io_diffCommits_info_374_ldest;
    logic [7:0]   io_diffCommits_info_374_pdest;
    logic [5:0]   io_diffCommits_info_375_ldest;
    logic [7:0]   io_diffCommits_info_375_pdest;
    logic [5:0]   io_diffCommits_info_376_ldest;
    logic [7:0]   io_diffCommits_info_376_pdest;
    logic [5:0]   io_diffCommits_info_377_ldest;
    logic [7:0]   io_diffCommits_info_377_pdest;
    logic [5:0]   io_diffCommits_info_378_ldest;
    logic [7:0]   io_diffCommits_info_378_pdest;
    logic [5:0]   io_diffCommits_info_379_ldest;
    logic [7:0]   io_diffCommits_info_379_pdest;
    logic [5:0]   io_diffCommits_info_380_ldest;
    logic [7:0]   io_diffCommits_info_380_pdest;
    logic [5:0]   io_diffCommits_info_381_ldest;
    logic [7:0]   io_diffCommits_info_381_pdest;
    logic [5:0]   io_diffCommits_info_382_ldest;
    logic [7:0]   io_diffCommits_info_382_pdest;
    logic [5:0]   io_diffCommits_info_383_ldest;
    logic [7:0]   io_diffCommits_info_383_pdest;
    logic [5:0]   io_diffCommits_info_384_ldest;
    logic [7:0]   io_diffCommits_info_384_pdest;
    logic [5:0]   io_diffCommits_info_385_ldest;
    logic [7:0]   io_diffCommits_info_385_pdest;
    logic [5:0]   io_diffCommits_info_386_ldest;
    logic [7:0]   io_diffCommits_info_386_pdest;
    logic [5:0]   io_diffCommits_info_387_ldest;
    logic [7:0]   io_diffCommits_info_387_pdest;
    logic [5:0]   io_diffCommits_info_388_ldest;
    logic [7:0]   io_diffCommits_info_388_pdest;
    logic [5:0]   io_diffCommits_info_389_ldest;
    logic [7:0]   io_diffCommits_info_389_pdest;
    logic [3:0]   io_lsq_scommit       ;
    logic         io_lsq_pendingMMIOld ;
    logic         io_lsq_pendingst     ;
    logic         io_lsq_pendingPtr_flag;
    logic [7:0]   io_lsq_pendingPtr_value;
    logic         io_robDeqPtr_flag    ;
    logic [7:0]   io_robDeqPtr_value   ;
    logic         io_csr_fflags_valid  ;
    logic [4:0]   io_csr_fflags_bits   ;
    logic         io_csr_vxsat_valid   ;
    logic         io_csr_vxsat_bits    ;
    logic         io_csr_vstart_valid  ;
    logic [63:0]  io_csr_vstart_bits   ;
    logic         io_csr_dirty_fs      ;
    logic         io_csr_dirty_vs      ;
    logic [6:0]   io_csr_perfinfo_retiredInstr;
    logic         io_cpu_halt          ;
    logic         io_wfi_wfiReq        ;
    logic         io_toDecode_isResumeVType;
    logic         io_toDecode_walkToArchVType;
    logic         io_toDecode_walkVType_valid;
    logic         io_toDecode_walkVType_bits_illegal;
    logic         io_toDecode_walkVType_bits_vma;
    logic         io_toDecode_walkVType_bits_vta;
    logic [1:0]   io_toDecode_walkVType_bits_vsew;
    logic [2:0]   io_toDecode_walkVType_bits_vlmul;
    logic         io_toDecode_commitVType_vtype_valid;
    logic         io_toDecode_commitVType_vtype_bits_illegal;
    logic         io_toDecode_commitVType_vtype_bits_vma;
    logic         io_toDecode_commitVType_vtype_bits_vta;
    logic [1:0]   io_toDecode_commitVType_vtype_bits_vsew;
    logic [2:0]   io_toDecode_commitVType_vtype_bits_vlmul;
    logic         io_toDecode_commitVType_hasVsetvl;
    logic         io_readGPAMemAddr_valid;
    logic [5:0]   io_readGPAMemAddr_bits_ftqPtr_value;
    logic [3:0]   io_readGPAMemAddr_bits_ftqOffset;
    logic         io_toVecExcpMod_logicPhyRegMap_0_valid;
    logic [5:0]   io_toVecExcpMod_logicPhyRegMap_0_bits_lreg;
    logic [6:0]   io_toVecExcpMod_logicPhyRegMap_0_bits_preg;
    logic         io_toVecExcpMod_logicPhyRegMap_1_valid;
    logic [5:0]   io_toVecExcpMod_logicPhyRegMap_1_bits_lreg;
    logic [6:0]   io_toVecExcpMod_logicPhyRegMap_1_bits_preg;
    logic         io_toVecExcpMod_logicPhyRegMap_2_valid;
    logic [5:0]   io_toVecExcpMod_logicPhyRegMap_2_bits_lreg;
    logic [6:0]   io_toVecExcpMod_logicPhyRegMap_2_bits_preg;
    logic         io_toVecExcpMod_logicPhyRegMap_3_valid;
    logic [5:0]   io_toVecExcpMod_logicPhyRegMap_3_bits_lreg;
    logic [6:0]   io_toVecExcpMod_logicPhyRegMap_3_bits_preg;
    logic         io_toVecExcpMod_logicPhyRegMap_4_valid;
    logic [5:0]   io_toVecExcpMod_logicPhyRegMap_4_bits_lreg;
    logic [6:0]   io_toVecExcpMod_logicPhyRegMap_4_bits_preg;
    logic         io_toVecExcpMod_logicPhyRegMap_5_valid;
    logic [5:0]   io_toVecExcpMod_logicPhyRegMap_5_bits_lreg;
    logic [6:0]   io_toVecExcpMod_logicPhyRegMap_5_bits_preg;
    logic         io_toVecExcpMod_excpInfo_valid;
    logic [6:0]   io_toVecExcpMod_excpInfo_bits_vstart;
    logic [1:0]   io_toVecExcpMod_excpInfo_bits_vsew;
    logic [1:0]   io_toVecExcpMod_excpInfo_bits_veew;
    logic [2:0]   io_toVecExcpMod_excpInfo_bits_vlmul;
    logic [2:0]   io_toVecExcpMod_excpInfo_bits_nf;
    logic         io_toVecExcpMod_excpInfo_bits_isStride;
    logic         io_toVecExcpMod_excpInfo_bits_isIndexed;
    logic         io_toVecExcpMod_excpInfo_bits_isWhole;
    logic         io_toVecExcpMod_excpInfo_bits_isVlm;
    logic [49:0]  io_storeDebugInfo_1_pc;
    logic [5:0]   io_perf_0_value      ;
    logic [5:0]   io_perf_1_value      ;
    logic [5:0]   io_perf_2_value      ;
    logic [5:0]   io_perf_3_value      ;
    logic [5:0]   io_perf_4_value      ;
    logic [5:0]   io_perf_5_value      ;
    logic [5:0]   io_perf_6_value      ;
    logic [5:0]   io_perf_7_value      ;
    logic [5:0]   io_perf_8_value      ;
    logic [5:0]   io_perf_9_value      ;
    logic [5:0]   io_perf_10_value     ;
    logic [5:0]   io_perf_11_value     ;
    logic [5:0]   io_perf_12_value     ;
    logic [5:0]   io_perf_13_value     ;
    logic [5:0]   io_perf_14_value     ;
    logic [5:0]   io_perf_15_value     ;
    logic [5:0]   io_perf_16_value     ;
    logic [5:0]   io_perf_17_value     ;
    logic         io_error_0           ;

    clocking drv_cb @(posedge clk);
        `ifdef INTERFACE_ADD_DELAY
            default input #`DEF_SETUP_TIME output #`DEF_HOLD_TIME;
        `endif
        input  io_enq_canAccept;
        input  io_enq_canAcceptForDispatch;
        input  io_enq_isEmpty;
        input  io_flushOut_valid;
        input  io_flushOut_bits_isRVC;
        input  io_flushOut_bits_robIdx_flag;
        input  io_flushOut_bits_robIdx_value;
        input  io_flushOut_bits_ftqIdx_flag;
        input  io_flushOut_bits_ftqIdx_value;
        input  io_flushOut_bits_ftqOffset;
        input  io_flushOut_bits_level;
        input  io_exception_valid;
        input  io_exception_bits_instr;
        input  io_exception_bits_commitType;
        input  io_exception_bits_exceptionVec_0;
        input  io_exception_bits_exceptionVec_1;
        input  io_exception_bits_exceptionVec_2;
        input  io_exception_bits_exceptionVec_3;
        input  io_exception_bits_exceptionVec_4;
        input  io_exception_bits_exceptionVec_5;
        input  io_exception_bits_exceptionVec_6;
        input  io_exception_bits_exceptionVec_7;
        input  io_exception_bits_exceptionVec_8;
        input  io_exception_bits_exceptionVec_9;
        input  io_exception_bits_exceptionVec_10;
        input  io_exception_bits_exceptionVec_11;
        input  io_exception_bits_exceptionVec_12;
        input  io_exception_bits_exceptionVec_13;
        input  io_exception_bits_exceptionVec_14;
        input  io_exception_bits_exceptionVec_15;
        input  io_exception_bits_exceptionVec_16;
        input  io_exception_bits_exceptionVec_17;
        input  io_exception_bits_exceptionVec_18;
        input  io_exception_bits_exceptionVec_19;
        input  io_exception_bits_exceptionVec_20;
        input  io_exception_bits_exceptionVec_21;
        input  io_exception_bits_exceptionVec_22;
        input  io_exception_bits_exceptionVec_23;
        input  io_exception_bits_isPcBkpt;
        input  io_exception_bits_isFetchMalAddr;
        input  io_exception_bits_gpaddr;
        input  io_exception_bits_singleStep;
        input  io_exception_bits_crossPageIPFFix;
        input  io_exception_bits_isInterrupt;
        input  io_exception_bits_isHls;
        input  io_exception_bits_trigger;
        input  io_exception_bits_isForVSnonLeafPTE;
        input  io_commits_isCommit;
        input  io_commits_commitValid_0;
        input  io_commits_commitValid_1;
        input  io_commits_commitValid_2;
        input  io_commits_commitValid_3;
        input  io_commits_commitValid_4;
        input  io_commits_commitValid_5;
        input  io_commits_commitValid_6;
        input  io_commits_commitValid_7;
        input  io_commits_isWalk;
        input  io_commits_walkValid_0;
        input  io_commits_walkValid_1;
        input  io_commits_walkValid_2;
        input  io_commits_walkValid_3;
        input  io_commits_walkValid_4;
        input  io_commits_walkValid_5;
        input  io_commits_walkValid_6;
        input  io_commits_walkValid_7;
        input  io_commits_info_0_walk_v;
        input  io_commits_info_0_commit_v;
        input  io_commits_info_0_commit_w;
        input  io_commits_info_0_realDestSize;
        input  io_commits_info_0_interrupt_safe;
        input  io_commits_info_0_wflags;
        input  io_commits_info_0_fflags;
        input  io_commits_info_0_vxsat;
        input  io_commits_info_0_isRVC;
        input  io_commits_info_0_isVset;
        input  io_commits_info_0_isHls;
        input  io_commits_info_0_isVls;
        input  io_commits_info_0_vls;
        input  io_commits_info_0_mmio;
        input  io_commits_info_0_commitType;
        input  io_commits_info_0_ftqIdx_flag;
        input  io_commits_info_0_ftqIdx_value;
        input  io_commits_info_0_ftqOffset;
        input  io_commits_info_0_instrSize;
        input  io_commits_info_0_fpWen;
        input  io_commits_info_0_rfWen;
        input  io_commits_info_0_needFlush;
        input  io_commits_info_0_traceBlockInPipe_itype;
        input  io_commits_info_0_traceBlockInPipe_iretire;
        input  io_commits_info_0_traceBlockInPipe_ilastsize;
        input  io_commits_info_0_debug_pc;
        input  io_commits_info_0_debug_instr;
        input  io_commits_info_0_debug_ldest;
        input  io_commits_info_0_debug_pdest;
        input  io_commits_info_0_debug_otherPdest_0;
        input  io_commits_info_0_debug_otherPdest_1;
        input  io_commits_info_0_debug_otherPdest_2;
        input  io_commits_info_0_debug_otherPdest_3;
        input  io_commits_info_0_debug_otherPdest_4;
        input  io_commits_info_0_debug_otherPdest_5;
        input  io_commits_info_0_debug_otherPdest_6;
        input  io_commits_info_0_debug_fuType;
        input  io_commits_info_0_dirtyFs;
        input  io_commits_info_0_dirtyVs;
        input  io_commits_info_1_walk_v;
        input  io_commits_info_1_commit_v;
        input  io_commits_info_1_commit_w;
        input  io_commits_info_1_realDestSize;
        input  io_commits_info_1_interrupt_safe;
        input  io_commits_info_1_wflags;
        input  io_commits_info_1_fflags;
        input  io_commits_info_1_vxsat;
        input  io_commits_info_1_isRVC;
        input  io_commits_info_1_isVset;
        input  io_commits_info_1_isHls;
        input  io_commits_info_1_isVls;
        input  io_commits_info_1_vls;
        input  io_commits_info_1_mmio;
        input  io_commits_info_1_commitType;
        input  io_commits_info_1_ftqIdx_flag;
        input  io_commits_info_1_ftqIdx_value;
        input  io_commits_info_1_ftqOffset;
        input  io_commits_info_1_instrSize;
        input  io_commits_info_1_fpWen;
        input  io_commits_info_1_rfWen;
        input  io_commits_info_1_needFlush;
        input  io_commits_info_1_traceBlockInPipe_itype;
        input  io_commits_info_1_traceBlockInPipe_iretire;
        input  io_commits_info_1_traceBlockInPipe_ilastsize;
        input  io_commits_info_1_debug_pc;
        input  io_commits_info_1_debug_instr;
        input  io_commits_info_1_debug_ldest;
        input  io_commits_info_1_debug_pdest;
        input  io_commits_info_1_debug_otherPdest_0;
        input  io_commits_info_1_debug_otherPdest_1;
        input  io_commits_info_1_debug_otherPdest_2;
        input  io_commits_info_1_debug_otherPdest_3;
        input  io_commits_info_1_debug_otherPdest_4;
        input  io_commits_info_1_debug_otherPdest_5;
        input  io_commits_info_1_debug_otherPdest_6;
        input  io_commits_info_1_debug_fuType;
        input  io_commits_info_1_dirtyFs;
        input  io_commits_info_1_dirtyVs;
        input  io_commits_info_2_walk_v;
        input  io_commits_info_2_commit_v;
        input  io_commits_info_2_commit_w;
        input  io_commits_info_2_realDestSize;
        input  io_commits_info_2_interrupt_safe;
        input  io_commits_info_2_wflags;
        input  io_commits_info_2_fflags;
        input  io_commits_info_2_vxsat;
        input  io_commits_info_2_isRVC;
        input  io_commits_info_2_isVset;
        input  io_commits_info_2_isHls;
        input  io_commits_info_2_isVls;
        input  io_commits_info_2_vls;
        input  io_commits_info_2_mmio;
        input  io_commits_info_2_commitType;
        input  io_commits_info_2_ftqIdx_flag;
        input  io_commits_info_2_ftqIdx_value;
        input  io_commits_info_2_ftqOffset;
        input  io_commits_info_2_instrSize;
        input  io_commits_info_2_fpWen;
        input  io_commits_info_2_rfWen;
        input  io_commits_info_2_needFlush;
        input  io_commits_info_2_traceBlockInPipe_itype;
        input  io_commits_info_2_traceBlockInPipe_iretire;
        input  io_commits_info_2_traceBlockInPipe_ilastsize;
        input  io_commits_info_2_debug_pc;
        input  io_commits_info_2_debug_instr;
        input  io_commits_info_2_debug_ldest;
        input  io_commits_info_2_debug_pdest;
        input  io_commits_info_2_debug_otherPdest_0;
        input  io_commits_info_2_debug_otherPdest_1;
        input  io_commits_info_2_debug_otherPdest_2;
        input  io_commits_info_2_debug_otherPdest_3;
        input  io_commits_info_2_debug_otherPdest_4;
        input  io_commits_info_2_debug_otherPdest_5;
        input  io_commits_info_2_debug_otherPdest_6;
        input  io_commits_info_2_debug_fuType;
        input  io_commits_info_2_dirtyFs;
        input  io_commits_info_2_dirtyVs;
        input  io_commits_info_3_walk_v;
        input  io_commits_info_3_commit_v;
        input  io_commits_info_3_commit_w;
        input  io_commits_info_3_realDestSize;
        input  io_commits_info_3_interrupt_safe;
        input  io_commits_info_3_wflags;
        input  io_commits_info_3_fflags;
        input  io_commits_info_3_vxsat;
        input  io_commits_info_3_isRVC;
        input  io_commits_info_3_isVset;
        input  io_commits_info_3_isHls;
        input  io_commits_info_3_isVls;
        input  io_commits_info_3_vls;
        input  io_commits_info_3_mmio;
        input  io_commits_info_3_commitType;
        input  io_commits_info_3_ftqIdx_flag;
        input  io_commits_info_3_ftqIdx_value;
        input  io_commits_info_3_ftqOffset;
        input  io_commits_info_3_instrSize;
        input  io_commits_info_3_fpWen;
        input  io_commits_info_3_rfWen;
        input  io_commits_info_3_needFlush;
        input  io_commits_info_3_traceBlockInPipe_itype;
        input  io_commits_info_3_traceBlockInPipe_iretire;
        input  io_commits_info_3_traceBlockInPipe_ilastsize;
        input  io_commits_info_3_debug_pc;
        input  io_commits_info_3_debug_instr;
        input  io_commits_info_3_debug_ldest;
        input  io_commits_info_3_debug_pdest;
        input  io_commits_info_3_debug_otherPdest_0;
        input  io_commits_info_3_debug_otherPdest_1;
        input  io_commits_info_3_debug_otherPdest_2;
        input  io_commits_info_3_debug_otherPdest_3;
        input  io_commits_info_3_debug_otherPdest_4;
        input  io_commits_info_3_debug_otherPdest_5;
        input  io_commits_info_3_debug_otherPdest_6;
        input  io_commits_info_3_debug_fuType;
        input  io_commits_info_3_dirtyFs;
        input  io_commits_info_3_dirtyVs;
        input  io_commits_info_4_walk_v;
        input  io_commits_info_4_commit_v;
        input  io_commits_info_4_commit_w;
        input  io_commits_info_4_realDestSize;
        input  io_commits_info_4_interrupt_safe;
        input  io_commits_info_4_wflags;
        input  io_commits_info_4_fflags;
        input  io_commits_info_4_vxsat;
        input  io_commits_info_4_isRVC;
        input  io_commits_info_4_isVset;
        input  io_commits_info_4_isHls;
        input  io_commits_info_4_isVls;
        input  io_commits_info_4_vls;
        input  io_commits_info_4_mmio;
        input  io_commits_info_4_commitType;
        input  io_commits_info_4_ftqIdx_flag;
        input  io_commits_info_4_ftqIdx_value;
        input  io_commits_info_4_ftqOffset;
        input  io_commits_info_4_instrSize;
        input  io_commits_info_4_fpWen;
        input  io_commits_info_4_rfWen;
        input  io_commits_info_4_needFlush;
        input  io_commits_info_4_traceBlockInPipe_itype;
        input  io_commits_info_4_traceBlockInPipe_iretire;
        input  io_commits_info_4_traceBlockInPipe_ilastsize;
        input  io_commits_info_4_debug_pc;
        input  io_commits_info_4_debug_instr;
        input  io_commits_info_4_debug_ldest;
        input  io_commits_info_4_debug_pdest;
        input  io_commits_info_4_debug_otherPdest_0;
        input  io_commits_info_4_debug_otherPdest_1;
        input  io_commits_info_4_debug_otherPdest_2;
        input  io_commits_info_4_debug_otherPdest_3;
        input  io_commits_info_4_debug_otherPdest_4;
        input  io_commits_info_4_debug_otherPdest_5;
        input  io_commits_info_4_debug_otherPdest_6;
        input  io_commits_info_4_debug_fuType;
        input  io_commits_info_4_dirtyFs;
        input  io_commits_info_4_dirtyVs;
        input  io_commits_info_5_walk_v;
        input  io_commits_info_5_commit_v;
        input  io_commits_info_5_commit_w;
        input  io_commits_info_5_realDestSize;
        input  io_commits_info_5_interrupt_safe;
        input  io_commits_info_5_wflags;
        input  io_commits_info_5_fflags;
        input  io_commits_info_5_vxsat;
        input  io_commits_info_5_isRVC;
        input  io_commits_info_5_isVset;
        input  io_commits_info_5_isHls;
        input  io_commits_info_5_isVls;
        input  io_commits_info_5_vls;
        input  io_commits_info_5_mmio;
        input  io_commits_info_5_commitType;
        input  io_commits_info_5_ftqIdx_flag;
        input  io_commits_info_5_ftqIdx_value;
        input  io_commits_info_5_ftqOffset;
        input  io_commits_info_5_instrSize;
        input  io_commits_info_5_fpWen;
        input  io_commits_info_5_rfWen;
        input  io_commits_info_5_needFlush;
        input  io_commits_info_5_traceBlockInPipe_itype;
        input  io_commits_info_5_traceBlockInPipe_iretire;
        input  io_commits_info_5_traceBlockInPipe_ilastsize;
        input  io_commits_info_5_debug_pc;
        input  io_commits_info_5_debug_instr;
        input  io_commits_info_5_debug_ldest;
        input  io_commits_info_5_debug_pdest;
        input  io_commits_info_5_debug_otherPdest_0;
        input  io_commits_info_5_debug_otherPdest_1;
        input  io_commits_info_5_debug_otherPdest_2;
        input  io_commits_info_5_debug_otherPdest_3;
        input  io_commits_info_5_debug_otherPdest_4;
        input  io_commits_info_5_debug_otherPdest_5;
        input  io_commits_info_5_debug_otherPdest_6;
        input  io_commits_info_5_debug_fuType;
        input  io_commits_info_5_dirtyFs;
        input  io_commits_info_5_dirtyVs;
        input  io_commits_info_6_walk_v;
        input  io_commits_info_6_commit_v;
        input  io_commits_info_6_commit_w;
        input  io_commits_info_6_realDestSize;
        input  io_commits_info_6_interrupt_safe;
        input  io_commits_info_6_wflags;
        input  io_commits_info_6_fflags;
        input  io_commits_info_6_vxsat;
        input  io_commits_info_6_isRVC;
        input  io_commits_info_6_isVset;
        input  io_commits_info_6_isHls;
        input  io_commits_info_6_isVls;
        input  io_commits_info_6_vls;
        input  io_commits_info_6_mmio;
        input  io_commits_info_6_commitType;
        input  io_commits_info_6_ftqIdx_flag;
        input  io_commits_info_6_ftqIdx_value;
        input  io_commits_info_6_ftqOffset;
        input  io_commits_info_6_instrSize;
        input  io_commits_info_6_fpWen;
        input  io_commits_info_6_rfWen;
        input  io_commits_info_6_needFlush;
        input  io_commits_info_6_traceBlockInPipe_itype;
        input  io_commits_info_6_traceBlockInPipe_iretire;
        input  io_commits_info_6_traceBlockInPipe_ilastsize;
        input  io_commits_info_6_debug_pc;
        input  io_commits_info_6_debug_instr;
        input  io_commits_info_6_debug_ldest;
        input  io_commits_info_6_debug_pdest;
        input  io_commits_info_6_debug_otherPdest_0;
        input  io_commits_info_6_debug_otherPdest_1;
        input  io_commits_info_6_debug_otherPdest_2;
        input  io_commits_info_6_debug_otherPdest_3;
        input  io_commits_info_6_debug_otherPdest_4;
        input  io_commits_info_6_debug_otherPdest_5;
        input  io_commits_info_6_debug_otherPdest_6;
        input  io_commits_info_6_debug_fuType;
        input  io_commits_info_6_dirtyFs;
        input  io_commits_info_6_dirtyVs;
        input  io_commits_info_7_walk_v;
        input  io_commits_info_7_commit_v;
        input  io_commits_info_7_commit_w;
        input  io_commits_info_7_realDestSize;
        input  io_commits_info_7_interrupt_safe;
        input  io_commits_info_7_wflags;
        input  io_commits_info_7_fflags;
        input  io_commits_info_7_vxsat;
        input  io_commits_info_7_isRVC;
        input  io_commits_info_7_isVset;
        input  io_commits_info_7_isHls;
        input  io_commits_info_7_isVls;
        input  io_commits_info_7_vls;
        input  io_commits_info_7_mmio;
        input  io_commits_info_7_commitType;
        input  io_commits_info_7_ftqIdx_flag;
        input  io_commits_info_7_ftqIdx_value;
        input  io_commits_info_7_ftqOffset;
        input  io_commits_info_7_instrSize;
        input  io_commits_info_7_fpWen;
        input  io_commits_info_7_rfWen;
        input  io_commits_info_7_needFlush;
        input  io_commits_info_7_traceBlockInPipe_itype;
        input  io_commits_info_7_traceBlockInPipe_iretire;
        input  io_commits_info_7_traceBlockInPipe_ilastsize;
        input  io_commits_info_7_debug_pc;
        input  io_commits_info_7_debug_instr;
        input  io_commits_info_7_debug_ldest;
        input  io_commits_info_7_debug_pdest;
        input  io_commits_info_7_debug_otherPdest_0;
        input  io_commits_info_7_debug_otherPdest_1;
        input  io_commits_info_7_debug_otherPdest_2;
        input  io_commits_info_7_debug_otherPdest_3;
        input  io_commits_info_7_debug_otherPdest_4;
        input  io_commits_info_7_debug_otherPdest_5;
        input  io_commits_info_7_debug_otherPdest_6;
        input  io_commits_info_7_debug_fuType;
        input  io_commits_info_7_dirtyFs;
        input  io_commits_info_7_dirtyVs;
        input  io_commits_robIdx_0_flag;
        input  io_commits_robIdx_0_value;
        input  io_commits_robIdx_1_flag;
        input  io_commits_robIdx_1_value;
        input  io_commits_robIdx_2_flag;
        input  io_commits_robIdx_2_value;
        input  io_commits_robIdx_3_flag;
        input  io_commits_robIdx_3_value;
        input  io_commits_robIdx_4_flag;
        input  io_commits_robIdx_4_value;
        input  io_commits_robIdx_5_flag;
        input  io_commits_robIdx_5_value;
        input  io_commits_robIdx_6_flag;
        input  io_commits_robIdx_6_value;
        input  io_commits_robIdx_7_flag;
        input  io_commits_robIdx_7_value;
        output io_trace_blockCommit;
        input  io_trace_traceCommitInfo_blocks_0_valid;
        input  io_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value;
        input  io_trace_traceCommitInfo_blocks_0_bits_ftqOffset;
        input  io_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype;
        input  io_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire;
        input  io_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize;
        input  io_trace_traceCommitInfo_blocks_1_valid;
        input  io_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value;
        input  io_trace_traceCommitInfo_blocks_1_bits_ftqOffset;
        input  io_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype;
        input  io_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire;
        input  io_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize;
        input  io_trace_traceCommitInfo_blocks_2_valid;
        input  io_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value;
        input  io_trace_traceCommitInfo_blocks_2_bits_ftqOffset;
        input  io_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype;
        input  io_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire;
        input  io_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize;
        input  io_trace_traceCommitInfo_blocks_3_valid;
        input  io_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value;
        input  io_trace_traceCommitInfo_blocks_3_bits_ftqOffset;
        input  io_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype;
        input  io_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire;
        input  io_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize;
        input  io_trace_traceCommitInfo_blocks_4_valid;
        input  io_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value;
        input  io_trace_traceCommitInfo_blocks_4_bits_ftqOffset;
        input  io_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype;
        input  io_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire;
        input  io_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize;
        input  io_trace_traceCommitInfo_blocks_5_valid;
        input  io_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value;
        input  io_trace_traceCommitInfo_blocks_5_bits_ftqOffset;
        input  io_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype;
        input  io_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire;
        input  io_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize;
        input  io_trace_traceCommitInfo_blocks_6_valid;
        input  io_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value;
        input  io_trace_traceCommitInfo_blocks_6_bits_ftqOffset;
        input  io_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype;
        input  io_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire;
        input  io_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize;
        input  io_trace_traceCommitInfo_blocks_7_valid;
        input  io_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value;
        input  io_trace_traceCommitInfo_blocks_7_bits_ftqOffset;
        input  io_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype;
        input  io_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire;
        input  io_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize;
        input  io_rabCommits_isCommit;
        input  io_rabCommits_commitValid_0;
        input  io_rabCommits_commitValid_1;
        input  io_rabCommits_commitValid_2;
        input  io_rabCommits_commitValid_3;
        input  io_rabCommits_commitValid_4;
        input  io_rabCommits_commitValid_5;
        input  io_rabCommits_isWalk;
        input  io_rabCommits_walkValid_0;
        input  io_rabCommits_walkValid_1;
        input  io_rabCommits_walkValid_2;
        input  io_rabCommits_walkValid_3;
        input  io_rabCommits_walkValid_4;
        input  io_rabCommits_walkValid_5;
        input  io_rabCommits_info_0_ldest;
        input  io_rabCommits_info_0_pdest;
        input  io_rabCommits_info_0_rfWen;
        input  io_rabCommits_info_0_fpWen;
        input  io_rabCommits_info_0_vecWen;
        input  io_rabCommits_info_0_v0Wen;
        input  io_rabCommits_info_0_vlWen;
        input  io_rabCommits_info_0_isMove;
        input  io_rabCommits_info_1_ldest;
        input  io_rabCommits_info_1_pdest;
        input  io_rabCommits_info_1_rfWen;
        input  io_rabCommits_info_1_fpWen;
        input  io_rabCommits_info_1_vecWen;
        input  io_rabCommits_info_1_v0Wen;
        input  io_rabCommits_info_1_vlWen;
        input  io_rabCommits_info_1_isMove;
        input  io_rabCommits_info_2_ldest;
        input  io_rabCommits_info_2_pdest;
        input  io_rabCommits_info_2_rfWen;
        input  io_rabCommits_info_2_fpWen;
        input  io_rabCommits_info_2_vecWen;
        input  io_rabCommits_info_2_v0Wen;
        input  io_rabCommits_info_2_vlWen;
        input  io_rabCommits_info_2_isMove;
        input  io_rabCommits_info_3_ldest;
        input  io_rabCommits_info_3_pdest;
        input  io_rabCommits_info_3_rfWen;
        input  io_rabCommits_info_3_fpWen;
        input  io_rabCommits_info_3_vecWen;
        input  io_rabCommits_info_3_v0Wen;
        input  io_rabCommits_info_3_vlWen;
        input  io_rabCommits_info_3_isMove;
        input  io_rabCommits_info_4_ldest;
        input  io_rabCommits_info_4_pdest;
        input  io_rabCommits_info_4_rfWen;
        input  io_rabCommits_info_4_fpWen;
        input  io_rabCommits_info_4_vecWen;
        input  io_rabCommits_info_4_v0Wen;
        input  io_rabCommits_info_4_vlWen;
        input  io_rabCommits_info_4_isMove;
        input  io_rabCommits_info_5_ldest;
        input  io_rabCommits_info_5_pdest;
        input  io_rabCommits_info_5_rfWen;
        input  io_rabCommits_info_5_fpWen;
        input  io_rabCommits_info_5_vecWen;
        input  io_rabCommits_info_5_v0Wen;
        input  io_rabCommits_info_5_vlWen;
        input  io_rabCommits_info_5_isMove;
        input  io_diffCommits_commitValid_0;
        input  io_diffCommits_commitValid_1;
        input  io_diffCommits_commitValid_2;
        input  io_diffCommits_commitValid_3;
        input  io_diffCommits_commitValid_4;
        input  io_diffCommits_commitValid_5;
        input  io_diffCommits_commitValid_6;
        input  io_diffCommits_commitValid_7;
        input  io_diffCommits_commitValid_8;
        input  io_diffCommits_commitValid_9;
        input  io_diffCommits_commitValid_10;
        input  io_diffCommits_commitValid_11;
        input  io_diffCommits_commitValid_12;
        input  io_diffCommits_commitValid_13;
        input  io_diffCommits_commitValid_14;
        input  io_diffCommits_commitValid_15;
        input  io_diffCommits_commitValid_16;
        input  io_diffCommits_commitValid_17;
        input  io_diffCommits_commitValid_18;
        input  io_diffCommits_commitValid_19;
        input  io_diffCommits_commitValid_20;
        input  io_diffCommits_commitValid_21;
        input  io_diffCommits_commitValid_22;
        input  io_diffCommits_commitValid_23;
        input  io_diffCommits_commitValid_24;
        input  io_diffCommits_commitValid_25;
        input  io_diffCommits_commitValid_26;
        input  io_diffCommits_commitValid_27;
        input  io_diffCommits_commitValid_28;
        input  io_diffCommits_commitValid_29;
        input  io_diffCommits_commitValid_30;
        input  io_diffCommits_commitValid_31;
        input  io_diffCommits_commitValid_32;
        input  io_diffCommits_commitValid_33;
        input  io_diffCommits_commitValid_34;
        input  io_diffCommits_commitValid_35;
        input  io_diffCommits_commitValid_36;
        input  io_diffCommits_commitValid_37;
        input  io_diffCommits_commitValid_38;
        input  io_diffCommits_commitValid_39;
        input  io_diffCommits_commitValid_40;
        input  io_diffCommits_commitValid_41;
        input  io_diffCommits_commitValid_42;
        input  io_diffCommits_commitValid_43;
        input  io_diffCommits_commitValid_44;
        input  io_diffCommits_commitValid_45;
        input  io_diffCommits_commitValid_46;
        input  io_diffCommits_commitValid_47;
        input  io_diffCommits_commitValid_48;
        input  io_diffCommits_commitValid_49;
        input  io_diffCommits_commitValid_50;
        input  io_diffCommits_commitValid_51;
        input  io_diffCommits_commitValid_52;
        input  io_diffCommits_commitValid_53;
        input  io_diffCommits_commitValid_54;
        input  io_diffCommits_commitValid_55;
        input  io_diffCommits_commitValid_56;
        input  io_diffCommits_commitValid_57;
        input  io_diffCommits_commitValid_58;
        input  io_diffCommits_commitValid_59;
        input  io_diffCommits_commitValid_60;
        input  io_diffCommits_commitValid_61;
        input  io_diffCommits_commitValid_62;
        input  io_diffCommits_commitValid_63;
        input  io_diffCommits_commitValid_64;
        input  io_diffCommits_commitValid_65;
        input  io_diffCommits_commitValid_66;
        input  io_diffCommits_commitValid_67;
        input  io_diffCommits_commitValid_68;
        input  io_diffCommits_commitValid_69;
        input  io_diffCommits_commitValid_70;
        input  io_diffCommits_commitValid_71;
        input  io_diffCommits_commitValid_72;
        input  io_diffCommits_commitValid_73;
        input  io_diffCommits_commitValid_74;
        input  io_diffCommits_commitValid_75;
        input  io_diffCommits_commitValid_76;
        input  io_diffCommits_commitValid_77;
        input  io_diffCommits_commitValid_78;
        input  io_diffCommits_commitValid_79;
        input  io_diffCommits_commitValid_80;
        input  io_diffCommits_commitValid_81;
        input  io_diffCommits_commitValid_82;
        input  io_diffCommits_commitValid_83;
        input  io_diffCommits_commitValid_84;
        input  io_diffCommits_commitValid_85;
        input  io_diffCommits_commitValid_86;
        input  io_diffCommits_commitValid_87;
        input  io_diffCommits_commitValid_88;
        input  io_diffCommits_commitValid_89;
        input  io_diffCommits_commitValid_90;
        input  io_diffCommits_commitValid_91;
        input  io_diffCommits_commitValid_92;
        input  io_diffCommits_commitValid_93;
        input  io_diffCommits_commitValid_94;
        input  io_diffCommits_commitValid_95;
        input  io_diffCommits_commitValid_96;
        input  io_diffCommits_commitValid_97;
        input  io_diffCommits_commitValid_98;
        input  io_diffCommits_commitValid_99;
        input  io_diffCommits_commitValid_100;
        input  io_diffCommits_commitValid_101;
        input  io_diffCommits_commitValid_102;
        input  io_diffCommits_commitValid_103;
        input  io_diffCommits_commitValid_104;
        input  io_diffCommits_commitValid_105;
        input  io_diffCommits_commitValid_106;
        input  io_diffCommits_commitValid_107;
        input  io_diffCommits_commitValid_108;
        input  io_diffCommits_commitValid_109;
        input  io_diffCommits_commitValid_110;
        input  io_diffCommits_commitValid_111;
        input  io_diffCommits_commitValid_112;
        input  io_diffCommits_commitValid_113;
        input  io_diffCommits_commitValid_114;
        input  io_diffCommits_commitValid_115;
        input  io_diffCommits_commitValid_116;
        input  io_diffCommits_commitValid_117;
        input  io_diffCommits_commitValid_118;
        input  io_diffCommits_commitValid_119;
        input  io_diffCommits_commitValid_120;
        input  io_diffCommits_commitValid_121;
        input  io_diffCommits_commitValid_122;
        input  io_diffCommits_commitValid_123;
        input  io_diffCommits_commitValid_124;
        input  io_diffCommits_commitValid_125;
        input  io_diffCommits_commitValid_126;
        input  io_diffCommits_commitValid_127;
        input  io_diffCommits_commitValid_128;
        input  io_diffCommits_commitValid_129;
        input  io_diffCommits_commitValid_130;
        input  io_diffCommits_commitValid_131;
        input  io_diffCommits_commitValid_132;
        input  io_diffCommits_commitValid_133;
        input  io_diffCommits_commitValid_134;
        input  io_diffCommits_commitValid_135;
        input  io_diffCommits_commitValid_136;
        input  io_diffCommits_commitValid_137;
        input  io_diffCommits_commitValid_138;
        input  io_diffCommits_commitValid_139;
        input  io_diffCommits_commitValid_140;
        input  io_diffCommits_commitValid_141;
        input  io_diffCommits_commitValid_142;
        input  io_diffCommits_commitValid_143;
        input  io_diffCommits_commitValid_144;
        input  io_diffCommits_commitValid_145;
        input  io_diffCommits_commitValid_146;
        input  io_diffCommits_commitValid_147;
        input  io_diffCommits_commitValid_148;
        input  io_diffCommits_commitValid_149;
        input  io_diffCommits_commitValid_150;
        input  io_diffCommits_commitValid_151;
        input  io_diffCommits_commitValid_152;
        input  io_diffCommits_commitValid_153;
        input  io_diffCommits_commitValid_154;
        input  io_diffCommits_commitValid_155;
        input  io_diffCommits_commitValid_156;
        input  io_diffCommits_commitValid_157;
        input  io_diffCommits_commitValid_158;
        input  io_diffCommits_commitValid_159;
        input  io_diffCommits_commitValid_160;
        input  io_diffCommits_commitValid_161;
        input  io_diffCommits_commitValid_162;
        input  io_diffCommits_commitValid_163;
        input  io_diffCommits_commitValid_164;
        input  io_diffCommits_commitValid_165;
        input  io_diffCommits_commitValid_166;
        input  io_diffCommits_commitValid_167;
        input  io_diffCommits_commitValid_168;
        input  io_diffCommits_commitValid_169;
        input  io_diffCommits_commitValid_170;
        input  io_diffCommits_commitValid_171;
        input  io_diffCommits_commitValid_172;
        input  io_diffCommits_commitValid_173;
        input  io_diffCommits_commitValid_174;
        input  io_diffCommits_commitValid_175;
        input  io_diffCommits_commitValid_176;
        input  io_diffCommits_commitValid_177;
        input  io_diffCommits_commitValid_178;
        input  io_diffCommits_commitValid_179;
        input  io_diffCommits_commitValid_180;
        input  io_diffCommits_commitValid_181;
        input  io_diffCommits_commitValid_182;
        input  io_diffCommits_commitValid_183;
        input  io_diffCommits_commitValid_184;
        input  io_diffCommits_commitValid_185;
        input  io_diffCommits_commitValid_186;
        input  io_diffCommits_commitValid_187;
        input  io_diffCommits_commitValid_188;
        input  io_diffCommits_commitValid_189;
        input  io_diffCommits_commitValid_190;
        input  io_diffCommits_commitValid_191;
        input  io_diffCommits_commitValid_192;
        input  io_diffCommits_commitValid_193;
        input  io_diffCommits_commitValid_194;
        input  io_diffCommits_commitValid_195;
        input  io_diffCommits_commitValid_196;
        input  io_diffCommits_commitValid_197;
        input  io_diffCommits_commitValid_198;
        input  io_diffCommits_commitValid_199;
        input  io_diffCommits_commitValid_200;
        input  io_diffCommits_commitValid_201;
        input  io_diffCommits_commitValid_202;
        input  io_diffCommits_commitValid_203;
        input  io_diffCommits_commitValid_204;
        input  io_diffCommits_commitValid_205;
        input  io_diffCommits_commitValid_206;
        input  io_diffCommits_commitValid_207;
        input  io_diffCommits_commitValid_208;
        input  io_diffCommits_commitValid_209;
        input  io_diffCommits_commitValid_210;
        input  io_diffCommits_commitValid_211;
        input  io_diffCommits_commitValid_212;
        input  io_diffCommits_commitValid_213;
        input  io_diffCommits_commitValid_214;
        input  io_diffCommits_commitValid_215;
        input  io_diffCommits_commitValid_216;
        input  io_diffCommits_commitValid_217;
        input  io_diffCommits_commitValid_218;
        input  io_diffCommits_commitValid_219;
        input  io_diffCommits_commitValid_220;
        input  io_diffCommits_commitValid_221;
        input  io_diffCommits_commitValid_222;
        input  io_diffCommits_commitValid_223;
        input  io_diffCommits_commitValid_224;
        input  io_diffCommits_commitValid_225;
        input  io_diffCommits_commitValid_226;
        input  io_diffCommits_commitValid_227;
        input  io_diffCommits_commitValid_228;
        input  io_diffCommits_commitValid_229;
        input  io_diffCommits_commitValid_230;
        input  io_diffCommits_commitValid_231;
        input  io_diffCommits_commitValid_232;
        input  io_diffCommits_commitValid_233;
        input  io_diffCommits_commitValid_234;
        input  io_diffCommits_commitValid_235;
        input  io_diffCommits_commitValid_236;
        input  io_diffCommits_commitValid_237;
        input  io_diffCommits_commitValid_238;
        input  io_diffCommits_commitValid_239;
        input  io_diffCommits_commitValid_240;
        input  io_diffCommits_commitValid_241;
        input  io_diffCommits_commitValid_242;
        input  io_diffCommits_commitValid_243;
        input  io_diffCommits_commitValid_244;
        input  io_diffCommits_commitValid_245;
        input  io_diffCommits_commitValid_246;
        input  io_diffCommits_commitValid_247;
        input  io_diffCommits_commitValid_248;
        input  io_diffCommits_commitValid_249;
        input  io_diffCommits_commitValid_250;
        input  io_diffCommits_commitValid_251;
        input  io_diffCommits_commitValid_252;
        input  io_diffCommits_commitValid_253;
        input  io_diffCommits_commitValid_254;
        input  io_diffCommits_info_0_ldest;
        input  io_diffCommits_info_0_pdest;
        input  io_diffCommits_info_0_rfWen;
        input  io_diffCommits_info_0_fpWen;
        input  io_diffCommits_info_0_vecWen;
        input  io_diffCommits_info_0_v0Wen;
        input  io_diffCommits_info_0_vlWen;
        input  io_diffCommits_info_1_ldest;
        input  io_diffCommits_info_1_pdest;
        input  io_diffCommits_info_1_rfWen;
        input  io_diffCommits_info_1_fpWen;
        input  io_diffCommits_info_1_vecWen;
        input  io_diffCommits_info_1_v0Wen;
        input  io_diffCommits_info_1_vlWen;
        input  io_diffCommits_info_2_ldest;
        input  io_diffCommits_info_2_pdest;
        input  io_diffCommits_info_2_rfWen;
        input  io_diffCommits_info_2_fpWen;
        input  io_diffCommits_info_2_vecWen;
        input  io_diffCommits_info_2_v0Wen;
        input  io_diffCommits_info_2_vlWen;
        input  io_diffCommits_info_3_ldest;
        input  io_diffCommits_info_3_pdest;
        input  io_diffCommits_info_3_rfWen;
        input  io_diffCommits_info_3_fpWen;
        input  io_diffCommits_info_3_vecWen;
        input  io_diffCommits_info_3_v0Wen;
        input  io_diffCommits_info_3_vlWen;
        input  io_diffCommits_info_4_ldest;
        input  io_diffCommits_info_4_pdest;
        input  io_diffCommits_info_4_rfWen;
        input  io_diffCommits_info_4_fpWen;
        input  io_diffCommits_info_4_vecWen;
        input  io_diffCommits_info_4_v0Wen;
        input  io_diffCommits_info_4_vlWen;
        input  io_diffCommits_info_5_ldest;
        input  io_diffCommits_info_5_pdest;
        input  io_diffCommits_info_5_rfWen;
        input  io_diffCommits_info_5_fpWen;
        input  io_diffCommits_info_5_vecWen;
        input  io_diffCommits_info_5_v0Wen;
        input  io_diffCommits_info_5_vlWen;
        input  io_diffCommits_info_6_ldest;
        input  io_diffCommits_info_6_pdest;
        input  io_diffCommits_info_6_rfWen;
        input  io_diffCommits_info_6_fpWen;
        input  io_diffCommits_info_6_vecWen;
        input  io_diffCommits_info_6_v0Wen;
        input  io_diffCommits_info_6_vlWen;
        input  io_diffCommits_info_7_ldest;
        input  io_diffCommits_info_7_pdest;
        input  io_diffCommits_info_7_rfWen;
        input  io_diffCommits_info_7_fpWen;
        input  io_diffCommits_info_7_vecWen;
        input  io_diffCommits_info_7_v0Wen;
        input  io_diffCommits_info_7_vlWen;
        input  io_diffCommits_info_8_ldest;
        input  io_diffCommits_info_8_pdest;
        input  io_diffCommits_info_8_rfWen;
        input  io_diffCommits_info_8_fpWen;
        input  io_diffCommits_info_8_vecWen;
        input  io_diffCommits_info_8_v0Wen;
        input  io_diffCommits_info_8_vlWen;
        input  io_diffCommits_info_9_ldest;
        input  io_diffCommits_info_9_pdest;
        input  io_diffCommits_info_9_rfWen;
        input  io_diffCommits_info_9_fpWen;
        input  io_diffCommits_info_9_vecWen;
        input  io_diffCommits_info_9_v0Wen;
        input  io_diffCommits_info_9_vlWen;
        input  io_diffCommits_info_10_ldest;
        input  io_diffCommits_info_10_pdest;
        input  io_diffCommits_info_10_rfWen;
        input  io_diffCommits_info_10_fpWen;
        input  io_diffCommits_info_10_vecWen;
        input  io_diffCommits_info_10_v0Wen;
        input  io_diffCommits_info_10_vlWen;
        input  io_diffCommits_info_11_ldest;
        input  io_diffCommits_info_11_pdest;
        input  io_diffCommits_info_11_rfWen;
        input  io_diffCommits_info_11_fpWen;
        input  io_diffCommits_info_11_vecWen;
        input  io_diffCommits_info_11_v0Wen;
        input  io_diffCommits_info_11_vlWen;
        input  io_diffCommits_info_12_ldest;
        input  io_diffCommits_info_12_pdest;
        input  io_diffCommits_info_12_rfWen;
        input  io_diffCommits_info_12_fpWen;
        input  io_diffCommits_info_12_vecWen;
        input  io_diffCommits_info_12_v0Wen;
        input  io_diffCommits_info_12_vlWen;
        input  io_diffCommits_info_13_ldest;
        input  io_diffCommits_info_13_pdest;
        input  io_diffCommits_info_13_rfWen;
        input  io_diffCommits_info_13_fpWen;
        input  io_diffCommits_info_13_vecWen;
        input  io_diffCommits_info_13_v0Wen;
        input  io_diffCommits_info_13_vlWen;
        input  io_diffCommits_info_14_ldest;
        input  io_diffCommits_info_14_pdest;
        input  io_diffCommits_info_14_rfWen;
        input  io_diffCommits_info_14_fpWen;
        input  io_diffCommits_info_14_vecWen;
        input  io_diffCommits_info_14_v0Wen;
        input  io_diffCommits_info_14_vlWen;
        input  io_diffCommits_info_15_ldest;
        input  io_diffCommits_info_15_pdest;
        input  io_diffCommits_info_15_rfWen;
        input  io_diffCommits_info_15_fpWen;
        input  io_diffCommits_info_15_vecWen;
        input  io_diffCommits_info_15_v0Wen;
        input  io_diffCommits_info_15_vlWen;
        input  io_diffCommits_info_16_ldest;
        input  io_diffCommits_info_16_pdest;
        input  io_diffCommits_info_16_rfWen;
        input  io_diffCommits_info_16_fpWen;
        input  io_diffCommits_info_16_vecWen;
        input  io_diffCommits_info_16_v0Wen;
        input  io_diffCommits_info_16_vlWen;
        input  io_diffCommits_info_17_ldest;
        input  io_diffCommits_info_17_pdest;
        input  io_diffCommits_info_17_rfWen;
        input  io_diffCommits_info_17_fpWen;
        input  io_diffCommits_info_17_vecWen;
        input  io_diffCommits_info_17_v0Wen;
        input  io_diffCommits_info_17_vlWen;
        input  io_diffCommits_info_18_ldest;
        input  io_diffCommits_info_18_pdest;
        input  io_diffCommits_info_18_rfWen;
        input  io_diffCommits_info_18_fpWen;
        input  io_diffCommits_info_18_vecWen;
        input  io_diffCommits_info_18_v0Wen;
        input  io_diffCommits_info_18_vlWen;
        input  io_diffCommits_info_19_ldest;
        input  io_diffCommits_info_19_pdest;
        input  io_diffCommits_info_19_rfWen;
        input  io_diffCommits_info_19_fpWen;
        input  io_diffCommits_info_19_vecWen;
        input  io_diffCommits_info_19_v0Wen;
        input  io_diffCommits_info_19_vlWen;
        input  io_diffCommits_info_20_ldest;
        input  io_diffCommits_info_20_pdest;
        input  io_diffCommits_info_20_rfWen;
        input  io_diffCommits_info_20_fpWen;
        input  io_diffCommits_info_20_vecWen;
        input  io_diffCommits_info_20_v0Wen;
        input  io_diffCommits_info_20_vlWen;
        input  io_diffCommits_info_21_ldest;
        input  io_diffCommits_info_21_pdest;
        input  io_diffCommits_info_21_rfWen;
        input  io_diffCommits_info_21_fpWen;
        input  io_diffCommits_info_21_vecWen;
        input  io_diffCommits_info_21_v0Wen;
        input  io_diffCommits_info_21_vlWen;
        input  io_diffCommits_info_22_ldest;
        input  io_diffCommits_info_22_pdest;
        input  io_diffCommits_info_22_rfWen;
        input  io_diffCommits_info_22_fpWen;
        input  io_diffCommits_info_22_vecWen;
        input  io_diffCommits_info_22_v0Wen;
        input  io_diffCommits_info_22_vlWen;
        input  io_diffCommits_info_23_ldest;
        input  io_diffCommits_info_23_pdest;
        input  io_diffCommits_info_23_rfWen;
        input  io_diffCommits_info_23_fpWen;
        input  io_diffCommits_info_23_vecWen;
        input  io_diffCommits_info_23_v0Wen;
        input  io_diffCommits_info_23_vlWen;
        input  io_diffCommits_info_24_ldest;
        input  io_diffCommits_info_24_pdest;
        input  io_diffCommits_info_24_rfWen;
        input  io_diffCommits_info_24_fpWen;
        input  io_diffCommits_info_24_vecWen;
        input  io_diffCommits_info_24_v0Wen;
        input  io_diffCommits_info_24_vlWen;
        input  io_diffCommits_info_25_ldest;
        input  io_diffCommits_info_25_pdest;
        input  io_diffCommits_info_25_rfWen;
        input  io_diffCommits_info_25_fpWen;
        input  io_diffCommits_info_25_vecWen;
        input  io_diffCommits_info_25_v0Wen;
        input  io_diffCommits_info_25_vlWen;
        input  io_diffCommits_info_26_ldest;
        input  io_diffCommits_info_26_pdest;
        input  io_diffCommits_info_26_rfWen;
        input  io_diffCommits_info_26_fpWen;
        input  io_diffCommits_info_26_vecWen;
        input  io_diffCommits_info_26_v0Wen;
        input  io_diffCommits_info_26_vlWen;
        input  io_diffCommits_info_27_ldest;
        input  io_diffCommits_info_27_pdest;
        input  io_diffCommits_info_27_rfWen;
        input  io_diffCommits_info_27_fpWen;
        input  io_diffCommits_info_27_vecWen;
        input  io_diffCommits_info_27_v0Wen;
        input  io_diffCommits_info_27_vlWen;
        input  io_diffCommits_info_28_ldest;
        input  io_diffCommits_info_28_pdest;
        input  io_diffCommits_info_28_rfWen;
        input  io_diffCommits_info_28_fpWen;
        input  io_diffCommits_info_28_vecWen;
        input  io_diffCommits_info_28_v0Wen;
        input  io_diffCommits_info_28_vlWen;
        input  io_diffCommits_info_29_ldest;
        input  io_diffCommits_info_29_pdest;
        input  io_diffCommits_info_29_rfWen;
        input  io_diffCommits_info_29_fpWen;
        input  io_diffCommits_info_29_vecWen;
        input  io_diffCommits_info_29_v0Wen;
        input  io_diffCommits_info_29_vlWen;
        input  io_diffCommits_info_30_ldest;
        input  io_diffCommits_info_30_pdest;
        input  io_diffCommits_info_30_rfWen;
        input  io_diffCommits_info_30_fpWen;
        input  io_diffCommits_info_30_vecWen;
        input  io_diffCommits_info_30_v0Wen;
        input  io_diffCommits_info_30_vlWen;
        input  io_diffCommits_info_31_ldest;
        input  io_diffCommits_info_31_pdest;
        input  io_diffCommits_info_31_rfWen;
        input  io_diffCommits_info_31_fpWen;
        input  io_diffCommits_info_31_vecWen;
        input  io_diffCommits_info_31_v0Wen;
        input  io_diffCommits_info_31_vlWen;
        input  io_diffCommits_info_32_ldest;
        input  io_diffCommits_info_32_pdest;
        input  io_diffCommits_info_32_rfWen;
        input  io_diffCommits_info_32_fpWen;
        input  io_diffCommits_info_32_vecWen;
        input  io_diffCommits_info_32_v0Wen;
        input  io_diffCommits_info_32_vlWen;
        input  io_diffCommits_info_33_ldest;
        input  io_diffCommits_info_33_pdest;
        input  io_diffCommits_info_33_rfWen;
        input  io_diffCommits_info_33_fpWen;
        input  io_diffCommits_info_33_vecWen;
        input  io_diffCommits_info_33_v0Wen;
        input  io_diffCommits_info_33_vlWen;
        input  io_diffCommits_info_34_ldest;
        input  io_diffCommits_info_34_pdest;
        input  io_diffCommits_info_34_rfWen;
        input  io_diffCommits_info_34_fpWen;
        input  io_diffCommits_info_34_vecWen;
        input  io_diffCommits_info_34_v0Wen;
        input  io_diffCommits_info_34_vlWen;
        input  io_diffCommits_info_35_ldest;
        input  io_diffCommits_info_35_pdest;
        input  io_diffCommits_info_35_rfWen;
        input  io_diffCommits_info_35_fpWen;
        input  io_diffCommits_info_35_vecWen;
        input  io_diffCommits_info_35_v0Wen;
        input  io_diffCommits_info_35_vlWen;
        input  io_diffCommits_info_36_ldest;
        input  io_diffCommits_info_36_pdest;
        input  io_diffCommits_info_36_rfWen;
        input  io_diffCommits_info_36_fpWen;
        input  io_diffCommits_info_36_vecWen;
        input  io_diffCommits_info_36_v0Wen;
        input  io_diffCommits_info_36_vlWen;
        input  io_diffCommits_info_37_ldest;
        input  io_diffCommits_info_37_pdest;
        input  io_diffCommits_info_37_rfWen;
        input  io_diffCommits_info_37_fpWen;
        input  io_diffCommits_info_37_vecWen;
        input  io_diffCommits_info_37_v0Wen;
        input  io_diffCommits_info_37_vlWen;
        input  io_diffCommits_info_38_ldest;
        input  io_diffCommits_info_38_pdest;
        input  io_diffCommits_info_38_rfWen;
        input  io_diffCommits_info_38_fpWen;
        input  io_diffCommits_info_38_vecWen;
        input  io_diffCommits_info_38_v0Wen;
        input  io_diffCommits_info_38_vlWen;
        input  io_diffCommits_info_39_ldest;
        input  io_diffCommits_info_39_pdest;
        input  io_diffCommits_info_39_rfWen;
        input  io_diffCommits_info_39_fpWen;
        input  io_diffCommits_info_39_vecWen;
        input  io_diffCommits_info_39_v0Wen;
        input  io_diffCommits_info_39_vlWen;
        input  io_diffCommits_info_40_ldest;
        input  io_diffCommits_info_40_pdest;
        input  io_diffCommits_info_40_rfWen;
        input  io_diffCommits_info_40_fpWen;
        input  io_diffCommits_info_40_vecWen;
        input  io_diffCommits_info_40_v0Wen;
        input  io_diffCommits_info_40_vlWen;
        input  io_diffCommits_info_41_ldest;
        input  io_diffCommits_info_41_pdest;
        input  io_diffCommits_info_41_rfWen;
        input  io_diffCommits_info_41_fpWen;
        input  io_diffCommits_info_41_vecWen;
        input  io_diffCommits_info_41_v0Wen;
        input  io_diffCommits_info_41_vlWen;
        input  io_diffCommits_info_42_ldest;
        input  io_diffCommits_info_42_pdest;
        input  io_diffCommits_info_42_rfWen;
        input  io_diffCommits_info_42_fpWen;
        input  io_diffCommits_info_42_vecWen;
        input  io_diffCommits_info_42_v0Wen;
        input  io_diffCommits_info_42_vlWen;
        input  io_diffCommits_info_43_ldest;
        input  io_diffCommits_info_43_pdest;
        input  io_diffCommits_info_43_rfWen;
        input  io_diffCommits_info_43_fpWen;
        input  io_diffCommits_info_43_vecWen;
        input  io_diffCommits_info_43_v0Wen;
        input  io_diffCommits_info_43_vlWen;
        input  io_diffCommits_info_44_ldest;
        input  io_diffCommits_info_44_pdest;
        input  io_diffCommits_info_44_rfWen;
        input  io_diffCommits_info_44_fpWen;
        input  io_diffCommits_info_44_vecWen;
        input  io_diffCommits_info_44_v0Wen;
        input  io_diffCommits_info_44_vlWen;
        input  io_diffCommits_info_45_ldest;
        input  io_diffCommits_info_45_pdest;
        input  io_diffCommits_info_45_rfWen;
        input  io_diffCommits_info_45_fpWen;
        input  io_diffCommits_info_45_vecWen;
        input  io_diffCommits_info_45_v0Wen;
        input  io_diffCommits_info_45_vlWen;
        input  io_diffCommits_info_46_ldest;
        input  io_diffCommits_info_46_pdest;
        input  io_diffCommits_info_46_rfWen;
        input  io_diffCommits_info_46_fpWen;
        input  io_diffCommits_info_46_vecWen;
        input  io_diffCommits_info_46_v0Wen;
        input  io_diffCommits_info_46_vlWen;
        input  io_diffCommits_info_47_ldest;
        input  io_diffCommits_info_47_pdest;
        input  io_diffCommits_info_47_rfWen;
        input  io_diffCommits_info_47_fpWen;
        input  io_diffCommits_info_47_vecWen;
        input  io_diffCommits_info_47_v0Wen;
        input  io_diffCommits_info_47_vlWen;
        input  io_diffCommits_info_48_ldest;
        input  io_diffCommits_info_48_pdest;
        input  io_diffCommits_info_48_rfWen;
        input  io_diffCommits_info_48_fpWen;
        input  io_diffCommits_info_48_vecWen;
        input  io_diffCommits_info_48_v0Wen;
        input  io_diffCommits_info_48_vlWen;
        input  io_diffCommits_info_49_ldest;
        input  io_diffCommits_info_49_pdest;
        input  io_diffCommits_info_49_rfWen;
        input  io_diffCommits_info_49_fpWen;
        input  io_diffCommits_info_49_vecWen;
        input  io_diffCommits_info_49_v0Wen;
        input  io_diffCommits_info_49_vlWen;
        input  io_diffCommits_info_50_ldest;
        input  io_diffCommits_info_50_pdest;
        input  io_diffCommits_info_50_rfWen;
        input  io_diffCommits_info_50_fpWen;
        input  io_diffCommits_info_50_vecWen;
        input  io_diffCommits_info_50_v0Wen;
        input  io_diffCommits_info_50_vlWen;
        input  io_diffCommits_info_51_ldest;
        input  io_diffCommits_info_51_pdest;
        input  io_diffCommits_info_51_rfWen;
        input  io_diffCommits_info_51_fpWen;
        input  io_diffCommits_info_51_vecWen;
        input  io_diffCommits_info_51_v0Wen;
        input  io_diffCommits_info_51_vlWen;
        input  io_diffCommits_info_52_ldest;
        input  io_diffCommits_info_52_pdest;
        input  io_diffCommits_info_52_rfWen;
        input  io_diffCommits_info_52_fpWen;
        input  io_diffCommits_info_52_vecWen;
        input  io_diffCommits_info_52_v0Wen;
        input  io_diffCommits_info_52_vlWen;
        input  io_diffCommits_info_53_ldest;
        input  io_diffCommits_info_53_pdest;
        input  io_diffCommits_info_53_rfWen;
        input  io_diffCommits_info_53_fpWen;
        input  io_diffCommits_info_53_vecWen;
        input  io_diffCommits_info_53_v0Wen;
        input  io_diffCommits_info_53_vlWen;
        input  io_diffCommits_info_54_ldest;
        input  io_diffCommits_info_54_pdest;
        input  io_diffCommits_info_54_rfWen;
        input  io_diffCommits_info_54_fpWen;
        input  io_diffCommits_info_54_vecWen;
        input  io_diffCommits_info_54_v0Wen;
        input  io_diffCommits_info_54_vlWen;
        input  io_diffCommits_info_55_ldest;
        input  io_diffCommits_info_55_pdest;
        input  io_diffCommits_info_55_rfWen;
        input  io_diffCommits_info_55_fpWen;
        input  io_diffCommits_info_55_vecWen;
        input  io_diffCommits_info_55_v0Wen;
        input  io_diffCommits_info_55_vlWen;
        input  io_diffCommits_info_56_ldest;
        input  io_diffCommits_info_56_pdest;
        input  io_diffCommits_info_56_rfWen;
        input  io_diffCommits_info_56_fpWen;
        input  io_diffCommits_info_56_vecWen;
        input  io_diffCommits_info_56_v0Wen;
        input  io_diffCommits_info_56_vlWen;
        input  io_diffCommits_info_57_ldest;
        input  io_diffCommits_info_57_pdest;
        input  io_diffCommits_info_57_rfWen;
        input  io_diffCommits_info_57_fpWen;
        input  io_diffCommits_info_57_vecWen;
        input  io_diffCommits_info_57_v0Wen;
        input  io_diffCommits_info_57_vlWen;
        input  io_diffCommits_info_58_ldest;
        input  io_diffCommits_info_58_pdest;
        input  io_diffCommits_info_58_rfWen;
        input  io_diffCommits_info_58_fpWen;
        input  io_diffCommits_info_58_vecWen;
        input  io_diffCommits_info_58_v0Wen;
        input  io_diffCommits_info_58_vlWen;
        input  io_diffCommits_info_59_ldest;
        input  io_diffCommits_info_59_pdest;
        input  io_diffCommits_info_59_rfWen;
        input  io_diffCommits_info_59_fpWen;
        input  io_diffCommits_info_59_vecWen;
        input  io_diffCommits_info_59_v0Wen;
        input  io_diffCommits_info_59_vlWen;
        input  io_diffCommits_info_60_ldest;
        input  io_diffCommits_info_60_pdest;
        input  io_diffCommits_info_60_rfWen;
        input  io_diffCommits_info_60_fpWen;
        input  io_diffCommits_info_60_vecWen;
        input  io_diffCommits_info_60_v0Wen;
        input  io_diffCommits_info_60_vlWen;
        input  io_diffCommits_info_61_ldest;
        input  io_diffCommits_info_61_pdest;
        input  io_diffCommits_info_61_rfWen;
        input  io_diffCommits_info_61_fpWen;
        input  io_diffCommits_info_61_vecWen;
        input  io_diffCommits_info_61_v0Wen;
        input  io_diffCommits_info_61_vlWen;
        input  io_diffCommits_info_62_ldest;
        input  io_diffCommits_info_62_pdest;
        input  io_diffCommits_info_62_rfWen;
        input  io_diffCommits_info_62_fpWen;
        input  io_diffCommits_info_62_vecWen;
        input  io_diffCommits_info_62_v0Wen;
        input  io_diffCommits_info_62_vlWen;
        input  io_diffCommits_info_63_ldest;
        input  io_diffCommits_info_63_pdest;
        input  io_diffCommits_info_63_rfWen;
        input  io_diffCommits_info_63_fpWen;
        input  io_diffCommits_info_63_vecWen;
        input  io_diffCommits_info_63_v0Wen;
        input  io_diffCommits_info_63_vlWen;
        input  io_diffCommits_info_64_ldest;
        input  io_diffCommits_info_64_pdest;
        input  io_diffCommits_info_64_rfWen;
        input  io_diffCommits_info_64_fpWen;
        input  io_diffCommits_info_64_vecWen;
        input  io_diffCommits_info_64_v0Wen;
        input  io_diffCommits_info_64_vlWen;
        input  io_diffCommits_info_65_ldest;
        input  io_diffCommits_info_65_pdest;
        input  io_diffCommits_info_65_rfWen;
        input  io_diffCommits_info_65_fpWen;
        input  io_diffCommits_info_65_vecWen;
        input  io_diffCommits_info_65_v0Wen;
        input  io_diffCommits_info_65_vlWen;
        input  io_diffCommits_info_66_ldest;
        input  io_diffCommits_info_66_pdest;
        input  io_diffCommits_info_66_rfWen;
        input  io_diffCommits_info_66_fpWen;
        input  io_diffCommits_info_66_vecWen;
        input  io_diffCommits_info_66_v0Wen;
        input  io_diffCommits_info_66_vlWen;
        input  io_diffCommits_info_67_ldest;
        input  io_diffCommits_info_67_pdest;
        input  io_diffCommits_info_67_rfWen;
        input  io_diffCommits_info_67_fpWen;
        input  io_diffCommits_info_67_vecWen;
        input  io_diffCommits_info_67_v0Wen;
        input  io_diffCommits_info_67_vlWen;
        input  io_diffCommits_info_68_ldest;
        input  io_diffCommits_info_68_pdest;
        input  io_diffCommits_info_68_rfWen;
        input  io_diffCommits_info_68_fpWen;
        input  io_diffCommits_info_68_vecWen;
        input  io_diffCommits_info_68_v0Wen;
        input  io_diffCommits_info_68_vlWen;
        input  io_diffCommits_info_69_ldest;
        input  io_diffCommits_info_69_pdest;
        input  io_diffCommits_info_69_rfWen;
        input  io_diffCommits_info_69_fpWen;
        input  io_diffCommits_info_69_vecWen;
        input  io_diffCommits_info_69_v0Wen;
        input  io_diffCommits_info_69_vlWen;
        input  io_diffCommits_info_70_ldest;
        input  io_diffCommits_info_70_pdest;
        input  io_diffCommits_info_70_rfWen;
        input  io_diffCommits_info_70_fpWen;
        input  io_diffCommits_info_70_vecWen;
        input  io_diffCommits_info_70_v0Wen;
        input  io_diffCommits_info_70_vlWen;
        input  io_diffCommits_info_71_ldest;
        input  io_diffCommits_info_71_pdest;
        input  io_diffCommits_info_71_rfWen;
        input  io_diffCommits_info_71_fpWen;
        input  io_diffCommits_info_71_vecWen;
        input  io_diffCommits_info_71_v0Wen;
        input  io_diffCommits_info_71_vlWen;
        input  io_diffCommits_info_72_ldest;
        input  io_diffCommits_info_72_pdest;
        input  io_diffCommits_info_72_rfWen;
        input  io_diffCommits_info_72_fpWen;
        input  io_diffCommits_info_72_vecWen;
        input  io_diffCommits_info_72_v0Wen;
        input  io_diffCommits_info_72_vlWen;
        input  io_diffCommits_info_73_ldest;
        input  io_diffCommits_info_73_pdest;
        input  io_diffCommits_info_73_rfWen;
        input  io_diffCommits_info_73_fpWen;
        input  io_diffCommits_info_73_vecWen;
        input  io_diffCommits_info_73_v0Wen;
        input  io_diffCommits_info_73_vlWen;
        input  io_diffCommits_info_74_ldest;
        input  io_diffCommits_info_74_pdest;
        input  io_diffCommits_info_74_rfWen;
        input  io_diffCommits_info_74_fpWen;
        input  io_diffCommits_info_74_vecWen;
        input  io_diffCommits_info_74_v0Wen;
        input  io_diffCommits_info_74_vlWen;
        input  io_diffCommits_info_75_ldest;
        input  io_diffCommits_info_75_pdest;
        input  io_diffCommits_info_75_rfWen;
        input  io_diffCommits_info_75_fpWen;
        input  io_diffCommits_info_75_vecWen;
        input  io_diffCommits_info_75_v0Wen;
        input  io_diffCommits_info_75_vlWen;
        input  io_diffCommits_info_76_ldest;
        input  io_diffCommits_info_76_pdest;
        input  io_diffCommits_info_76_rfWen;
        input  io_diffCommits_info_76_fpWen;
        input  io_diffCommits_info_76_vecWen;
        input  io_diffCommits_info_76_v0Wen;
        input  io_diffCommits_info_76_vlWen;
        input  io_diffCommits_info_77_ldest;
        input  io_diffCommits_info_77_pdest;
        input  io_diffCommits_info_77_rfWen;
        input  io_diffCommits_info_77_fpWen;
        input  io_diffCommits_info_77_vecWen;
        input  io_diffCommits_info_77_v0Wen;
        input  io_diffCommits_info_77_vlWen;
        input  io_diffCommits_info_78_ldest;
        input  io_diffCommits_info_78_pdest;
        input  io_diffCommits_info_78_rfWen;
        input  io_diffCommits_info_78_fpWen;
        input  io_diffCommits_info_78_vecWen;
        input  io_diffCommits_info_78_v0Wen;
        input  io_diffCommits_info_78_vlWen;
        input  io_diffCommits_info_79_ldest;
        input  io_diffCommits_info_79_pdest;
        input  io_diffCommits_info_79_rfWen;
        input  io_diffCommits_info_79_fpWen;
        input  io_diffCommits_info_79_vecWen;
        input  io_diffCommits_info_79_v0Wen;
        input  io_diffCommits_info_79_vlWen;
        input  io_diffCommits_info_80_ldest;
        input  io_diffCommits_info_80_pdest;
        input  io_diffCommits_info_80_rfWen;
        input  io_diffCommits_info_80_fpWen;
        input  io_diffCommits_info_80_vecWen;
        input  io_diffCommits_info_80_v0Wen;
        input  io_diffCommits_info_80_vlWen;
        input  io_diffCommits_info_81_ldest;
        input  io_diffCommits_info_81_pdest;
        input  io_diffCommits_info_81_rfWen;
        input  io_diffCommits_info_81_fpWen;
        input  io_diffCommits_info_81_vecWen;
        input  io_diffCommits_info_81_v0Wen;
        input  io_diffCommits_info_81_vlWen;
        input  io_diffCommits_info_82_ldest;
        input  io_diffCommits_info_82_pdest;
        input  io_diffCommits_info_82_rfWen;
        input  io_diffCommits_info_82_fpWen;
        input  io_diffCommits_info_82_vecWen;
        input  io_diffCommits_info_82_v0Wen;
        input  io_diffCommits_info_82_vlWen;
        input  io_diffCommits_info_83_ldest;
        input  io_diffCommits_info_83_pdest;
        input  io_diffCommits_info_83_rfWen;
        input  io_diffCommits_info_83_fpWen;
        input  io_diffCommits_info_83_vecWen;
        input  io_diffCommits_info_83_v0Wen;
        input  io_diffCommits_info_83_vlWen;
        input  io_diffCommits_info_84_ldest;
        input  io_diffCommits_info_84_pdest;
        input  io_diffCommits_info_84_rfWen;
        input  io_diffCommits_info_84_fpWen;
        input  io_diffCommits_info_84_vecWen;
        input  io_diffCommits_info_84_v0Wen;
        input  io_diffCommits_info_84_vlWen;
        input  io_diffCommits_info_85_ldest;
        input  io_diffCommits_info_85_pdest;
        input  io_diffCommits_info_85_rfWen;
        input  io_diffCommits_info_85_fpWen;
        input  io_diffCommits_info_85_vecWen;
        input  io_diffCommits_info_85_v0Wen;
        input  io_diffCommits_info_85_vlWen;
        input  io_diffCommits_info_86_ldest;
        input  io_diffCommits_info_86_pdest;
        input  io_diffCommits_info_86_rfWen;
        input  io_diffCommits_info_86_fpWen;
        input  io_diffCommits_info_86_vecWen;
        input  io_diffCommits_info_86_v0Wen;
        input  io_diffCommits_info_86_vlWen;
        input  io_diffCommits_info_87_ldest;
        input  io_diffCommits_info_87_pdest;
        input  io_diffCommits_info_87_rfWen;
        input  io_diffCommits_info_87_fpWen;
        input  io_diffCommits_info_87_vecWen;
        input  io_diffCommits_info_87_v0Wen;
        input  io_diffCommits_info_87_vlWen;
        input  io_diffCommits_info_88_ldest;
        input  io_diffCommits_info_88_pdest;
        input  io_diffCommits_info_88_rfWen;
        input  io_diffCommits_info_88_fpWen;
        input  io_diffCommits_info_88_vecWen;
        input  io_diffCommits_info_88_v0Wen;
        input  io_diffCommits_info_88_vlWen;
        input  io_diffCommits_info_89_ldest;
        input  io_diffCommits_info_89_pdest;
        input  io_diffCommits_info_89_rfWen;
        input  io_diffCommits_info_89_fpWen;
        input  io_diffCommits_info_89_vecWen;
        input  io_diffCommits_info_89_v0Wen;
        input  io_diffCommits_info_89_vlWen;
        input  io_diffCommits_info_90_ldest;
        input  io_diffCommits_info_90_pdest;
        input  io_diffCommits_info_90_rfWen;
        input  io_diffCommits_info_90_fpWen;
        input  io_diffCommits_info_90_vecWen;
        input  io_diffCommits_info_90_v0Wen;
        input  io_diffCommits_info_90_vlWen;
        input  io_diffCommits_info_91_ldest;
        input  io_diffCommits_info_91_pdest;
        input  io_diffCommits_info_91_rfWen;
        input  io_diffCommits_info_91_fpWen;
        input  io_diffCommits_info_91_vecWen;
        input  io_diffCommits_info_91_v0Wen;
        input  io_diffCommits_info_91_vlWen;
        input  io_diffCommits_info_92_ldest;
        input  io_diffCommits_info_92_pdest;
        input  io_diffCommits_info_92_rfWen;
        input  io_diffCommits_info_92_fpWen;
        input  io_diffCommits_info_92_vecWen;
        input  io_diffCommits_info_92_v0Wen;
        input  io_diffCommits_info_92_vlWen;
        input  io_diffCommits_info_93_ldest;
        input  io_diffCommits_info_93_pdest;
        input  io_diffCommits_info_93_rfWen;
        input  io_diffCommits_info_93_fpWen;
        input  io_diffCommits_info_93_vecWen;
        input  io_diffCommits_info_93_v0Wen;
        input  io_diffCommits_info_93_vlWen;
        input  io_diffCommits_info_94_ldest;
        input  io_diffCommits_info_94_pdest;
        input  io_diffCommits_info_94_rfWen;
        input  io_diffCommits_info_94_fpWen;
        input  io_diffCommits_info_94_vecWen;
        input  io_diffCommits_info_94_v0Wen;
        input  io_diffCommits_info_94_vlWen;
        input  io_diffCommits_info_95_ldest;
        input  io_diffCommits_info_95_pdest;
        input  io_diffCommits_info_95_rfWen;
        input  io_diffCommits_info_95_fpWen;
        input  io_diffCommits_info_95_vecWen;
        input  io_diffCommits_info_95_v0Wen;
        input  io_diffCommits_info_95_vlWen;
        input  io_diffCommits_info_96_ldest;
        input  io_diffCommits_info_96_pdest;
        input  io_diffCommits_info_96_rfWen;
        input  io_diffCommits_info_96_fpWen;
        input  io_diffCommits_info_96_vecWen;
        input  io_diffCommits_info_96_v0Wen;
        input  io_diffCommits_info_96_vlWen;
        input  io_diffCommits_info_97_ldest;
        input  io_diffCommits_info_97_pdest;
        input  io_diffCommits_info_97_rfWen;
        input  io_diffCommits_info_97_fpWen;
        input  io_diffCommits_info_97_vecWen;
        input  io_diffCommits_info_97_v0Wen;
        input  io_diffCommits_info_97_vlWen;
        input  io_diffCommits_info_98_ldest;
        input  io_diffCommits_info_98_pdest;
        input  io_diffCommits_info_98_rfWen;
        input  io_diffCommits_info_98_fpWen;
        input  io_diffCommits_info_98_vecWen;
        input  io_diffCommits_info_98_v0Wen;
        input  io_diffCommits_info_98_vlWen;
        input  io_diffCommits_info_99_ldest;
        input  io_diffCommits_info_99_pdest;
        input  io_diffCommits_info_99_rfWen;
        input  io_diffCommits_info_99_fpWen;
        input  io_diffCommits_info_99_vecWen;
        input  io_diffCommits_info_99_v0Wen;
        input  io_diffCommits_info_99_vlWen;
        input  io_diffCommits_info_100_ldest;
        input  io_diffCommits_info_100_pdest;
        input  io_diffCommits_info_100_rfWen;
        input  io_diffCommits_info_100_fpWen;
        input  io_diffCommits_info_100_vecWen;
        input  io_diffCommits_info_100_v0Wen;
        input  io_diffCommits_info_100_vlWen;
        input  io_diffCommits_info_101_ldest;
        input  io_diffCommits_info_101_pdest;
        input  io_diffCommits_info_101_rfWen;
        input  io_diffCommits_info_101_fpWen;
        input  io_diffCommits_info_101_vecWen;
        input  io_diffCommits_info_101_v0Wen;
        input  io_diffCommits_info_101_vlWen;
        input  io_diffCommits_info_102_ldest;
        input  io_diffCommits_info_102_pdest;
        input  io_diffCommits_info_102_rfWen;
        input  io_diffCommits_info_102_fpWen;
        input  io_diffCommits_info_102_vecWen;
        input  io_diffCommits_info_102_v0Wen;
        input  io_diffCommits_info_102_vlWen;
        input  io_diffCommits_info_103_ldest;
        input  io_diffCommits_info_103_pdest;
        input  io_diffCommits_info_103_rfWen;
        input  io_diffCommits_info_103_fpWen;
        input  io_diffCommits_info_103_vecWen;
        input  io_diffCommits_info_103_v0Wen;
        input  io_diffCommits_info_103_vlWen;
        input  io_diffCommits_info_104_ldest;
        input  io_diffCommits_info_104_pdest;
        input  io_diffCommits_info_104_rfWen;
        input  io_diffCommits_info_104_fpWen;
        input  io_diffCommits_info_104_vecWen;
        input  io_diffCommits_info_104_v0Wen;
        input  io_diffCommits_info_104_vlWen;
        input  io_diffCommits_info_105_ldest;
        input  io_diffCommits_info_105_pdest;
        input  io_diffCommits_info_105_rfWen;
        input  io_diffCommits_info_105_fpWen;
        input  io_diffCommits_info_105_vecWen;
        input  io_diffCommits_info_105_v0Wen;
        input  io_diffCommits_info_105_vlWen;
        input  io_diffCommits_info_106_ldest;
        input  io_diffCommits_info_106_pdest;
        input  io_diffCommits_info_106_rfWen;
        input  io_diffCommits_info_106_fpWen;
        input  io_diffCommits_info_106_vecWen;
        input  io_diffCommits_info_106_v0Wen;
        input  io_diffCommits_info_106_vlWen;
        input  io_diffCommits_info_107_ldest;
        input  io_diffCommits_info_107_pdest;
        input  io_diffCommits_info_107_rfWen;
        input  io_diffCommits_info_107_fpWen;
        input  io_diffCommits_info_107_vecWen;
        input  io_diffCommits_info_107_v0Wen;
        input  io_diffCommits_info_107_vlWen;
        input  io_diffCommits_info_108_ldest;
        input  io_diffCommits_info_108_pdest;
        input  io_diffCommits_info_108_rfWen;
        input  io_diffCommits_info_108_fpWen;
        input  io_diffCommits_info_108_vecWen;
        input  io_diffCommits_info_108_v0Wen;
        input  io_diffCommits_info_108_vlWen;
        input  io_diffCommits_info_109_ldest;
        input  io_diffCommits_info_109_pdest;
        input  io_diffCommits_info_109_rfWen;
        input  io_diffCommits_info_109_fpWen;
        input  io_diffCommits_info_109_vecWen;
        input  io_diffCommits_info_109_v0Wen;
        input  io_diffCommits_info_109_vlWen;
        input  io_diffCommits_info_110_ldest;
        input  io_diffCommits_info_110_pdest;
        input  io_diffCommits_info_110_rfWen;
        input  io_diffCommits_info_110_fpWen;
        input  io_diffCommits_info_110_vecWen;
        input  io_diffCommits_info_110_v0Wen;
        input  io_diffCommits_info_110_vlWen;
        input  io_diffCommits_info_111_ldest;
        input  io_diffCommits_info_111_pdest;
        input  io_diffCommits_info_111_rfWen;
        input  io_diffCommits_info_111_fpWen;
        input  io_diffCommits_info_111_vecWen;
        input  io_diffCommits_info_111_v0Wen;
        input  io_diffCommits_info_111_vlWen;
        input  io_diffCommits_info_112_ldest;
        input  io_diffCommits_info_112_pdest;
        input  io_diffCommits_info_112_rfWen;
        input  io_diffCommits_info_112_fpWen;
        input  io_diffCommits_info_112_vecWen;
        input  io_diffCommits_info_112_v0Wen;
        input  io_diffCommits_info_112_vlWen;
        input  io_diffCommits_info_113_ldest;
        input  io_diffCommits_info_113_pdest;
        input  io_diffCommits_info_113_rfWen;
        input  io_diffCommits_info_113_fpWen;
        input  io_diffCommits_info_113_vecWen;
        input  io_diffCommits_info_113_v0Wen;
        input  io_diffCommits_info_113_vlWen;
        input  io_diffCommits_info_114_ldest;
        input  io_diffCommits_info_114_pdest;
        input  io_diffCommits_info_114_rfWen;
        input  io_diffCommits_info_114_fpWen;
        input  io_diffCommits_info_114_vecWen;
        input  io_diffCommits_info_114_v0Wen;
        input  io_diffCommits_info_114_vlWen;
        input  io_diffCommits_info_115_ldest;
        input  io_diffCommits_info_115_pdest;
        input  io_diffCommits_info_115_rfWen;
        input  io_diffCommits_info_115_fpWen;
        input  io_diffCommits_info_115_vecWen;
        input  io_diffCommits_info_115_v0Wen;
        input  io_diffCommits_info_115_vlWen;
        input  io_diffCommits_info_116_ldest;
        input  io_diffCommits_info_116_pdest;
        input  io_diffCommits_info_116_rfWen;
        input  io_diffCommits_info_116_fpWen;
        input  io_diffCommits_info_116_vecWen;
        input  io_diffCommits_info_116_v0Wen;
        input  io_diffCommits_info_116_vlWen;
        input  io_diffCommits_info_117_ldest;
        input  io_diffCommits_info_117_pdest;
        input  io_diffCommits_info_117_rfWen;
        input  io_diffCommits_info_117_fpWen;
        input  io_diffCommits_info_117_vecWen;
        input  io_diffCommits_info_117_v0Wen;
        input  io_diffCommits_info_117_vlWen;
        input  io_diffCommits_info_118_ldest;
        input  io_diffCommits_info_118_pdest;
        input  io_diffCommits_info_118_rfWen;
        input  io_diffCommits_info_118_fpWen;
        input  io_diffCommits_info_118_vecWen;
        input  io_diffCommits_info_118_v0Wen;
        input  io_diffCommits_info_118_vlWen;
        input  io_diffCommits_info_119_ldest;
        input  io_diffCommits_info_119_pdest;
        input  io_diffCommits_info_119_rfWen;
        input  io_diffCommits_info_119_fpWen;
        input  io_diffCommits_info_119_vecWen;
        input  io_diffCommits_info_119_v0Wen;
        input  io_diffCommits_info_119_vlWen;
        input  io_diffCommits_info_120_ldest;
        input  io_diffCommits_info_120_pdest;
        input  io_diffCommits_info_120_rfWen;
        input  io_diffCommits_info_120_fpWen;
        input  io_diffCommits_info_120_vecWen;
        input  io_diffCommits_info_120_v0Wen;
        input  io_diffCommits_info_120_vlWen;
        input  io_diffCommits_info_121_ldest;
        input  io_diffCommits_info_121_pdest;
        input  io_diffCommits_info_121_rfWen;
        input  io_diffCommits_info_121_fpWen;
        input  io_diffCommits_info_121_vecWen;
        input  io_diffCommits_info_121_v0Wen;
        input  io_diffCommits_info_121_vlWen;
        input  io_diffCommits_info_122_ldest;
        input  io_diffCommits_info_122_pdest;
        input  io_diffCommits_info_122_rfWen;
        input  io_diffCommits_info_122_fpWen;
        input  io_diffCommits_info_122_vecWen;
        input  io_diffCommits_info_122_v0Wen;
        input  io_diffCommits_info_122_vlWen;
        input  io_diffCommits_info_123_ldest;
        input  io_diffCommits_info_123_pdest;
        input  io_diffCommits_info_123_rfWen;
        input  io_diffCommits_info_123_fpWen;
        input  io_diffCommits_info_123_vecWen;
        input  io_diffCommits_info_123_v0Wen;
        input  io_diffCommits_info_123_vlWen;
        input  io_diffCommits_info_124_ldest;
        input  io_diffCommits_info_124_pdest;
        input  io_diffCommits_info_124_rfWen;
        input  io_diffCommits_info_124_fpWen;
        input  io_diffCommits_info_124_vecWen;
        input  io_diffCommits_info_124_v0Wen;
        input  io_diffCommits_info_124_vlWen;
        input  io_diffCommits_info_125_ldest;
        input  io_diffCommits_info_125_pdest;
        input  io_diffCommits_info_125_rfWen;
        input  io_diffCommits_info_125_fpWen;
        input  io_diffCommits_info_125_vecWen;
        input  io_diffCommits_info_125_v0Wen;
        input  io_diffCommits_info_125_vlWen;
        input  io_diffCommits_info_126_ldest;
        input  io_diffCommits_info_126_pdest;
        input  io_diffCommits_info_126_rfWen;
        input  io_diffCommits_info_126_fpWen;
        input  io_diffCommits_info_126_vecWen;
        input  io_diffCommits_info_126_v0Wen;
        input  io_diffCommits_info_126_vlWen;
        input  io_diffCommits_info_127_ldest;
        input  io_diffCommits_info_127_pdest;
        input  io_diffCommits_info_127_rfWen;
        input  io_diffCommits_info_127_fpWen;
        input  io_diffCommits_info_127_vecWen;
        input  io_diffCommits_info_127_v0Wen;
        input  io_diffCommits_info_127_vlWen;
        input  io_diffCommits_info_128_ldest;
        input  io_diffCommits_info_128_pdest;
        input  io_diffCommits_info_128_rfWen;
        input  io_diffCommits_info_128_fpWen;
        input  io_diffCommits_info_128_vecWen;
        input  io_diffCommits_info_128_v0Wen;
        input  io_diffCommits_info_128_vlWen;
        input  io_diffCommits_info_129_ldest;
        input  io_diffCommits_info_129_pdest;
        input  io_diffCommits_info_129_rfWen;
        input  io_diffCommits_info_129_fpWen;
        input  io_diffCommits_info_129_vecWen;
        input  io_diffCommits_info_129_v0Wen;
        input  io_diffCommits_info_129_vlWen;
        input  io_diffCommits_info_130_ldest;
        input  io_diffCommits_info_130_pdest;
        input  io_diffCommits_info_130_rfWen;
        input  io_diffCommits_info_130_fpWen;
        input  io_diffCommits_info_130_vecWen;
        input  io_diffCommits_info_130_v0Wen;
        input  io_diffCommits_info_130_vlWen;
        input  io_diffCommits_info_131_ldest;
        input  io_diffCommits_info_131_pdest;
        input  io_diffCommits_info_131_rfWen;
        input  io_diffCommits_info_131_fpWen;
        input  io_diffCommits_info_131_vecWen;
        input  io_diffCommits_info_131_v0Wen;
        input  io_diffCommits_info_131_vlWen;
        input  io_diffCommits_info_132_ldest;
        input  io_diffCommits_info_132_pdest;
        input  io_diffCommits_info_132_rfWen;
        input  io_diffCommits_info_132_fpWen;
        input  io_diffCommits_info_132_vecWen;
        input  io_diffCommits_info_132_v0Wen;
        input  io_diffCommits_info_132_vlWen;
        input  io_diffCommits_info_133_ldest;
        input  io_diffCommits_info_133_pdest;
        input  io_diffCommits_info_133_rfWen;
        input  io_diffCommits_info_133_fpWen;
        input  io_diffCommits_info_133_vecWen;
        input  io_diffCommits_info_133_v0Wen;
        input  io_diffCommits_info_133_vlWen;
        input  io_diffCommits_info_134_ldest;
        input  io_diffCommits_info_134_pdest;
        input  io_diffCommits_info_134_rfWen;
        input  io_diffCommits_info_134_fpWen;
        input  io_diffCommits_info_134_vecWen;
        input  io_diffCommits_info_134_v0Wen;
        input  io_diffCommits_info_134_vlWen;
        input  io_diffCommits_info_135_ldest;
        input  io_diffCommits_info_135_pdest;
        input  io_diffCommits_info_135_rfWen;
        input  io_diffCommits_info_135_fpWen;
        input  io_diffCommits_info_135_vecWen;
        input  io_diffCommits_info_135_v0Wen;
        input  io_diffCommits_info_135_vlWen;
        input  io_diffCommits_info_136_ldest;
        input  io_diffCommits_info_136_pdest;
        input  io_diffCommits_info_136_rfWen;
        input  io_diffCommits_info_136_fpWen;
        input  io_diffCommits_info_136_vecWen;
        input  io_diffCommits_info_136_v0Wen;
        input  io_diffCommits_info_136_vlWen;
        input  io_diffCommits_info_137_ldest;
        input  io_diffCommits_info_137_pdest;
        input  io_diffCommits_info_137_rfWen;
        input  io_diffCommits_info_137_fpWen;
        input  io_diffCommits_info_137_vecWen;
        input  io_diffCommits_info_137_v0Wen;
        input  io_diffCommits_info_137_vlWen;
        input  io_diffCommits_info_138_ldest;
        input  io_diffCommits_info_138_pdest;
        input  io_diffCommits_info_138_rfWen;
        input  io_diffCommits_info_138_fpWen;
        input  io_diffCommits_info_138_vecWen;
        input  io_diffCommits_info_138_v0Wen;
        input  io_diffCommits_info_138_vlWen;
        input  io_diffCommits_info_139_ldest;
        input  io_diffCommits_info_139_pdest;
        input  io_diffCommits_info_139_rfWen;
        input  io_diffCommits_info_139_fpWen;
        input  io_diffCommits_info_139_vecWen;
        input  io_diffCommits_info_139_v0Wen;
        input  io_diffCommits_info_139_vlWen;
        input  io_diffCommits_info_140_ldest;
        input  io_diffCommits_info_140_pdest;
        input  io_diffCommits_info_140_rfWen;
        input  io_diffCommits_info_140_fpWen;
        input  io_diffCommits_info_140_vecWen;
        input  io_diffCommits_info_140_v0Wen;
        input  io_diffCommits_info_140_vlWen;
        input  io_diffCommits_info_141_ldest;
        input  io_diffCommits_info_141_pdest;
        input  io_diffCommits_info_141_rfWen;
        input  io_diffCommits_info_141_fpWen;
        input  io_diffCommits_info_141_vecWen;
        input  io_diffCommits_info_141_v0Wen;
        input  io_diffCommits_info_141_vlWen;
        input  io_diffCommits_info_142_ldest;
        input  io_diffCommits_info_142_pdest;
        input  io_diffCommits_info_142_rfWen;
        input  io_diffCommits_info_142_fpWen;
        input  io_diffCommits_info_142_vecWen;
        input  io_diffCommits_info_142_v0Wen;
        input  io_diffCommits_info_142_vlWen;
        input  io_diffCommits_info_143_ldest;
        input  io_diffCommits_info_143_pdest;
        input  io_diffCommits_info_143_rfWen;
        input  io_diffCommits_info_143_fpWen;
        input  io_diffCommits_info_143_vecWen;
        input  io_diffCommits_info_143_v0Wen;
        input  io_diffCommits_info_143_vlWen;
        input  io_diffCommits_info_144_ldest;
        input  io_diffCommits_info_144_pdest;
        input  io_diffCommits_info_144_rfWen;
        input  io_diffCommits_info_144_fpWen;
        input  io_diffCommits_info_144_vecWen;
        input  io_diffCommits_info_144_v0Wen;
        input  io_diffCommits_info_144_vlWen;
        input  io_diffCommits_info_145_ldest;
        input  io_diffCommits_info_145_pdest;
        input  io_diffCommits_info_145_rfWen;
        input  io_diffCommits_info_145_fpWen;
        input  io_diffCommits_info_145_vecWen;
        input  io_diffCommits_info_145_v0Wen;
        input  io_diffCommits_info_145_vlWen;
        input  io_diffCommits_info_146_ldest;
        input  io_diffCommits_info_146_pdest;
        input  io_diffCommits_info_146_rfWen;
        input  io_diffCommits_info_146_fpWen;
        input  io_diffCommits_info_146_vecWen;
        input  io_diffCommits_info_146_v0Wen;
        input  io_diffCommits_info_146_vlWen;
        input  io_diffCommits_info_147_ldest;
        input  io_diffCommits_info_147_pdest;
        input  io_diffCommits_info_147_rfWen;
        input  io_diffCommits_info_147_fpWen;
        input  io_diffCommits_info_147_vecWen;
        input  io_diffCommits_info_147_v0Wen;
        input  io_diffCommits_info_147_vlWen;
        input  io_diffCommits_info_148_ldest;
        input  io_diffCommits_info_148_pdest;
        input  io_diffCommits_info_148_rfWen;
        input  io_diffCommits_info_148_fpWen;
        input  io_diffCommits_info_148_vecWen;
        input  io_diffCommits_info_148_v0Wen;
        input  io_diffCommits_info_148_vlWen;
        input  io_diffCommits_info_149_ldest;
        input  io_diffCommits_info_149_pdest;
        input  io_diffCommits_info_149_rfWen;
        input  io_diffCommits_info_149_fpWen;
        input  io_diffCommits_info_149_vecWen;
        input  io_diffCommits_info_149_v0Wen;
        input  io_diffCommits_info_149_vlWen;
        input  io_diffCommits_info_150_ldest;
        input  io_diffCommits_info_150_pdest;
        input  io_diffCommits_info_150_rfWen;
        input  io_diffCommits_info_150_fpWen;
        input  io_diffCommits_info_150_vecWen;
        input  io_diffCommits_info_150_v0Wen;
        input  io_diffCommits_info_150_vlWen;
        input  io_diffCommits_info_151_ldest;
        input  io_diffCommits_info_151_pdest;
        input  io_diffCommits_info_151_rfWen;
        input  io_diffCommits_info_151_fpWen;
        input  io_diffCommits_info_151_vecWen;
        input  io_diffCommits_info_151_v0Wen;
        input  io_diffCommits_info_151_vlWen;
        input  io_diffCommits_info_152_ldest;
        input  io_diffCommits_info_152_pdest;
        input  io_diffCommits_info_152_rfWen;
        input  io_diffCommits_info_152_fpWen;
        input  io_diffCommits_info_152_vecWen;
        input  io_diffCommits_info_152_v0Wen;
        input  io_diffCommits_info_152_vlWen;
        input  io_diffCommits_info_153_ldest;
        input  io_diffCommits_info_153_pdest;
        input  io_diffCommits_info_153_rfWen;
        input  io_diffCommits_info_153_fpWen;
        input  io_diffCommits_info_153_vecWen;
        input  io_diffCommits_info_153_v0Wen;
        input  io_diffCommits_info_153_vlWen;
        input  io_diffCommits_info_154_ldest;
        input  io_diffCommits_info_154_pdest;
        input  io_diffCommits_info_154_rfWen;
        input  io_diffCommits_info_154_fpWen;
        input  io_diffCommits_info_154_vecWen;
        input  io_diffCommits_info_154_v0Wen;
        input  io_diffCommits_info_154_vlWen;
        input  io_diffCommits_info_155_ldest;
        input  io_diffCommits_info_155_pdest;
        input  io_diffCommits_info_155_rfWen;
        input  io_diffCommits_info_155_fpWen;
        input  io_diffCommits_info_155_vecWen;
        input  io_diffCommits_info_155_v0Wen;
        input  io_diffCommits_info_155_vlWen;
        input  io_diffCommits_info_156_ldest;
        input  io_diffCommits_info_156_pdest;
        input  io_diffCommits_info_156_rfWen;
        input  io_diffCommits_info_156_fpWen;
        input  io_diffCommits_info_156_vecWen;
        input  io_diffCommits_info_156_v0Wen;
        input  io_diffCommits_info_156_vlWen;
        input  io_diffCommits_info_157_ldest;
        input  io_diffCommits_info_157_pdest;
        input  io_diffCommits_info_157_rfWen;
        input  io_diffCommits_info_157_fpWen;
        input  io_diffCommits_info_157_vecWen;
        input  io_diffCommits_info_157_v0Wen;
        input  io_diffCommits_info_157_vlWen;
        input  io_diffCommits_info_158_ldest;
        input  io_diffCommits_info_158_pdest;
        input  io_diffCommits_info_158_rfWen;
        input  io_diffCommits_info_158_fpWen;
        input  io_diffCommits_info_158_vecWen;
        input  io_diffCommits_info_158_v0Wen;
        input  io_diffCommits_info_158_vlWen;
        input  io_diffCommits_info_159_ldest;
        input  io_diffCommits_info_159_pdest;
        input  io_diffCommits_info_159_rfWen;
        input  io_diffCommits_info_159_fpWen;
        input  io_diffCommits_info_159_vecWen;
        input  io_diffCommits_info_159_v0Wen;
        input  io_diffCommits_info_159_vlWen;
        input  io_diffCommits_info_160_ldest;
        input  io_diffCommits_info_160_pdest;
        input  io_diffCommits_info_160_rfWen;
        input  io_diffCommits_info_160_fpWen;
        input  io_diffCommits_info_160_vecWen;
        input  io_diffCommits_info_160_v0Wen;
        input  io_diffCommits_info_160_vlWen;
        input  io_diffCommits_info_161_ldest;
        input  io_diffCommits_info_161_pdest;
        input  io_diffCommits_info_161_rfWen;
        input  io_diffCommits_info_161_fpWen;
        input  io_diffCommits_info_161_vecWen;
        input  io_diffCommits_info_161_v0Wen;
        input  io_diffCommits_info_161_vlWen;
        input  io_diffCommits_info_162_ldest;
        input  io_diffCommits_info_162_pdest;
        input  io_diffCommits_info_162_rfWen;
        input  io_diffCommits_info_162_fpWen;
        input  io_diffCommits_info_162_vecWen;
        input  io_diffCommits_info_162_v0Wen;
        input  io_diffCommits_info_162_vlWen;
        input  io_diffCommits_info_163_ldest;
        input  io_diffCommits_info_163_pdest;
        input  io_diffCommits_info_163_rfWen;
        input  io_diffCommits_info_163_fpWen;
        input  io_diffCommits_info_163_vecWen;
        input  io_diffCommits_info_163_v0Wen;
        input  io_diffCommits_info_163_vlWen;
        input  io_diffCommits_info_164_ldest;
        input  io_diffCommits_info_164_pdest;
        input  io_diffCommits_info_164_rfWen;
        input  io_diffCommits_info_164_fpWen;
        input  io_diffCommits_info_164_vecWen;
        input  io_diffCommits_info_164_v0Wen;
        input  io_diffCommits_info_164_vlWen;
        input  io_diffCommits_info_165_ldest;
        input  io_diffCommits_info_165_pdest;
        input  io_diffCommits_info_165_rfWen;
        input  io_diffCommits_info_165_fpWen;
        input  io_diffCommits_info_165_vecWen;
        input  io_diffCommits_info_165_v0Wen;
        input  io_diffCommits_info_165_vlWen;
        input  io_diffCommits_info_166_ldest;
        input  io_diffCommits_info_166_pdest;
        input  io_diffCommits_info_166_rfWen;
        input  io_diffCommits_info_166_fpWen;
        input  io_diffCommits_info_166_vecWen;
        input  io_diffCommits_info_166_v0Wen;
        input  io_diffCommits_info_166_vlWen;
        input  io_diffCommits_info_167_ldest;
        input  io_diffCommits_info_167_pdest;
        input  io_diffCommits_info_167_rfWen;
        input  io_diffCommits_info_167_fpWen;
        input  io_diffCommits_info_167_vecWen;
        input  io_diffCommits_info_167_v0Wen;
        input  io_diffCommits_info_167_vlWen;
        input  io_diffCommits_info_168_ldest;
        input  io_diffCommits_info_168_pdest;
        input  io_diffCommits_info_168_rfWen;
        input  io_diffCommits_info_168_fpWen;
        input  io_diffCommits_info_168_vecWen;
        input  io_diffCommits_info_168_v0Wen;
        input  io_diffCommits_info_168_vlWen;
        input  io_diffCommits_info_169_ldest;
        input  io_diffCommits_info_169_pdest;
        input  io_diffCommits_info_169_rfWen;
        input  io_diffCommits_info_169_fpWen;
        input  io_diffCommits_info_169_vecWen;
        input  io_diffCommits_info_169_v0Wen;
        input  io_diffCommits_info_169_vlWen;
        input  io_diffCommits_info_170_ldest;
        input  io_diffCommits_info_170_pdest;
        input  io_diffCommits_info_170_rfWen;
        input  io_diffCommits_info_170_fpWen;
        input  io_diffCommits_info_170_vecWen;
        input  io_diffCommits_info_170_v0Wen;
        input  io_diffCommits_info_170_vlWen;
        input  io_diffCommits_info_171_ldest;
        input  io_diffCommits_info_171_pdest;
        input  io_diffCommits_info_171_rfWen;
        input  io_diffCommits_info_171_fpWen;
        input  io_diffCommits_info_171_vecWen;
        input  io_diffCommits_info_171_v0Wen;
        input  io_diffCommits_info_171_vlWen;
        input  io_diffCommits_info_172_ldest;
        input  io_diffCommits_info_172_pdest;
        input  io_diffCommits_info_172_rfWen;
        input  io_diffCommits_info_172_fpWen;
        input  io_diffCommits_info_172_vecWen;
        input  io_diffCommits_info_172_v0Wen;
        input  io_diffCommits_info_172_vlWen;
        input  io_diffCommits_info_173_ldest;
        input  io_diffCommits_info_173_pdest;
        input  io_diffCommits_info_173_rfWen;
        input  io_diffCommits_info_173_fpWen;
        input  io_diffCommits_info_173_vecWen;
        input  io_diffCommits_info_173_v0Wen;
        input  io_diffCommits_info_173_vlWen;
        input  io_diffCommits_info_174_ldest;
        input  io_diffCommits_info_174_pdest;
        input  io_diffCommits_info_174_rfWen;
        input  io_diffCommits_info_174_fpWen;
        input  io_diffCommits_info_174_vecWen;
        input  io_diffCommits_info_174_v0Wen;
        input  io_diffCommits_info_174_vlWen;
        input  io_diffCommits_info_175_ldest;
        input  io_diffCommits_info_175_pdest;
        input  io_diffCommits_info_175_rfWen;
        input  io_diffCommits_info_175_fpWen;
        input  io_diffCommits_info_175_vecWen;
        input  io_diffCommits_info_175_v0Wen;
        input  io_diffCommits_info_175_vlWen;
        input  io_diffCommits_info_176_ldest;
        input  io_diffCommits_info_176_pdest;
        input  io_diffCommits_info_176_rfWen;
        input  io_diffCommits_info_176_fpWen;
        input  io_diffCommits_info_176_vecWen;
        input  io_diffCommits_info_176_v0Wen;
        input  io_diffCommits_info_176_vlWen;
        input  io_diffCommits_info_177_ldest;
        input  io_diffCommits_info_177_pdest;
        input  io_diffCommits_info_177_rfWen;
        input  io_diffCommits_info_177_fpWen;
        input  io_diffCommits_info_177_vecWen;
        input  io_diffCommits_info_177_v0Wen;
        input  io_diffCommits_info_177_vlWen;
        input  io_diffCommits_info_178_ldest;
        input  io_diffCommits_info_178_pdest;
        input  io_diffCommits_info_178_rfWen;
        input  io_diffCommits_info_178_fpWen;
        input  io_diffCommits_info_178_vecWen;
        input  io_diffCommits_info_178_v0Wen;
        input  io_diffCommits_info_178_vlWen;
        input  io_diffCommits_info_179_ldest;
        input  io_diffCommits_info_179_pdest;
        input  io_diffCommits_info_179_rfWen;
        input  io_diffCommits_info_179_fpWen;
        input  io_diffCommits_info_179_vecWen;
        input  io_diffCommits_info_179_v0Wen;
        input  io_diffCommits_info_179_vlWen;
        input  io_diffCommits_info_180_ldest;
        input  io_diffCommits_info_180_pdest;
        input  io_diffCommits_info_180_rfWen;
        input  io_diffCommits_info_180_fpWen;
        input  io_diffCommits_info_180_vecWen;
        input  io_diffCommits_info_180_v0Wen;
        input  io_diffCommits_info_180_vlWen;
        input  io_diffCommits_info_181_ldest;
        input  io_diffCommits_info_181_pdest;
        input  io_diffCommits_info_181_rfWen;
        input  io_diffCommits_info_181_fpWen;
        input  io_diffCommits_info_181_vecWen;
        input  io_diffCommits_info_181_v0Wen;
        input  io_diffCommits_info_181_vlWen;
        input  io_diffCommits_info_182_ldest;
        input  io_diffCommits_info_182_pdest;
        input  io_diffCommits_info_182_rfWen;
        input  io_diffCommits_info_182_fpWen;
        input  io_diffCommits_info_182_vecWen;
        input  io_diffCommits_info_182_v0Wen;
        input  io_diffCommits_info_182_vlWen;
        input  io_diffCommits_info_183_ldest;
        input  io_diffCommits_info_183_pdest;
        input  io_diffCommits_info_183_rfWen;
        input  io_diffCommits_info_183_fpWen;
        input  io_diffCommits_info_183_vecWen;
        input  io_diffCommits_info_183_v0Wen;
        input  io_diffCommits_info_183_vlWen;
        input  io_diffCommits_info_184_ldest;
        input  io_diffCommits_info_184_pdest;
        input  io_diffCommits_info_184_rfWen;
        input  io_diffCommits_info_184_fpWen;
        input  io_diffCommits_info_184_vecWen;
        input  io_diffCommits_info_184_v0Wen;
        input  io_diffCommits_info_184_vlWen;
        input  io_diffCommits_info_185_ldest;
        input  io_diffCommits_info_185_pdest;
        input  io_diffCommits_info_185_rfWen;
        input  io_diffCommits_info_185_fpWen;
        input  io_diffCommits_info_185_vecWen;
        input  io_diffCommits_info_185_v0Wen;
        input  io_diffCommits_info_185_vlWen;
        input  io_diffCommits_info_186_ldest;
        input  io_diffCommits_info_186_pdest;
        input  io_diffCommits_info_186_rfWen;
        input  io_diffCommits_info_186_fpWen;
        input  io_diffCommits_info_186_vecWen;
        input  io_diffCommits_info_186_v0Wen;
        input  io_diffCommits_info_186_vlWen;
        input  io_diffCommits_info_187_ldest;
        input  io_diffCommits_info_187_pdest;
        input  io_diffCommits_info_187_rfWen;
        input  io_diffCommits_info_187_fpWen;
        input  io_diffCommits_info_187_vecWen;
        input  io_diffCommits_info_187_v0Wen;
        input  io_diffCommits_info_187_vlWen;
        input  io_diffCommits_info_188_ldest;
        input  io_diffCommits_info_188_pdest;
        input  io_diffCommits_info_188_rfWen;
        input  io_diffCommits_info_188_fpWen;
        input  io_diffCommits_info_188_vecWen;
        input  io_diffCommits_info_188_v0Wen;
        input  io_diffCommits_info_188_vlWen;
        input  io_diffCommits_info_189_ldest;
        input  io_diffCommits_info_189_pdest;
        input  io_diffCommits_info_189_rfWen;
        input  io_diffCommits_info_189_fpWen;
        input  io_diffCommits_info_189_vecWen;
        input  io_diffCommits_info_189_v0Wen;
        input  io_diffCommits_info_189_vlWen;
        input  io_diffCommits_info_190_ldest;
        input  io_diffCommits_info_190_pdest;
        input  io_diffCommits_info_190_rfWen;
        input  io_diffCommits_info_190_fpWen;
        input  io_diffCommits_info_190_vecWen;
        input  io_diffCommits_info_190_v0Wen;
        input  io_diffCommits_info_190_vlWen;
        input  io_diffCommits_info_191_ldest;
        input  io_diffCommits_info_191_pdest;
        input  io_diffCommits_info_191_rfWen;
        input  io_diffCommits_info_191_fpWen;
        input  io_diffCommits_info_191_vecWen;
        input  io_diffCommits_info_191_v0Wen;
        input  io_diffCommits_info_191_vlWen;
        input  io_diffCommits_info_192_ldest;
        input  io_diffCommits_info_192_pdest;
        input  io_diffCommits_info_192_rfWen;
        input  io_diffCommits_info_192_fpWen;
        input  io_diffCommits_info_192_vecWen;
        input  io_diffCommits_info_192_v0Wen;
        input  io_diffCommits_info_192_vlWen;
        input  io_diffCommits_info_193_ldest;
        input  io_diffCommits_info_193_pdest;
        input  io_diffCommits_info_193_rfWen;
        input  io_diffCommits_info_193_fpWen;
        input  io_diffCommits_info_193_vecWen;
        input  io_diffCommits_info_193_v0Wen;
        input  io_diffCommits_info_193_vlWen;
        input  io_diffCommits_info_194_ldest;
        input  io_diffCommits_info_194_pdest;
        input  io_diffCommits_info_194_rfWen;
        input  io_diffCommits_info_194_fpWen;
        input  io_diffCommits_info_194_vecWen;
        input  io_diffCommits_info_194_v0Wen;
        input  io_diffCommits_info_194_vlWen;
        input  io_diffCommits_info_195_ldest;
        input  io_diffCommits_info_195_pdest;
        input  io_diffCommits_info_195_rfWen;
        input  io_diffCommits_info_195_fpWen;
        input  io_diffCommits_info_195_vecWen;
        input  io_diffCommits_info_195_v0Wen;
        input  io_diffCommits_info_195_vlWen;
        input  io_diffCommits_info_196_ldest;
        input  io_diffCommits_info_196_pdest;
        input  io_diffCommits_info_196_rfWen;
        input  io_diffCommits_info_196_fpWen;
        input  io_diffCommits_info_196_vecWen;
        input  io_diffCommits_info_196_v0Wen;
        input  io_diffCommits_info_196_vlWen;
        input  io_diffCommits_info_197_ldest;
        input  io_diffCommits_info_197_pdest;
        input  io_diffCommits_info_197_rfWen;
        input  io_diffCommits_info_197_fpWen;
        input  io_diffCommits_info_197_vecWen;
        input  io_diffCommits_info_197_v0Wen;
        input  io_diffCommits_info_197_vlWen;
        input  io_diffCommits_info_198_ldest;
        input  io_diffCommits_info_198_pdest;
        input  io_diffCommits_info_198_rfWen;
        input  io_diffCommits_info_198_fpWen;
        input  io_diffCommits_info_198_vecWen;
        input  io_diffCommits_info_198_v0Wen;
        input  io_diffCommits_info_198_vlWen;
        input  io_diffCommits_info_199_ldest;
        input  io_diffCommits_info_199_pdest;
        input  io_diffCommits_info_199_rfWen;
        input  io_diffCommits_info_199_fpWen;
        input  io_diffCommits_info_199_vecWen;
        input  io_diffCommits_info_199_v0Wen;
        input  io_diffCommits_info_199_vlWen;
        input  io_diffCommits_info_200_ldest;
        input  io_diffCommits_info_200_pdest;
        input  io_diffCommits_info_200_rfWen;
        input  io_diffCommits_info_200_fpWen;
        input  io_diffCommits_info_200_vecWen;
        input  io_diffCommits_info_200_v0Wen;
        input  io_diffCommits_info_200_vlWen;
        input  io_diffCommits_info_201_ldest;
        input  io_diffCommits_info_201_pdest;
        input  io_diffCommits_info_201_rfWen;
        input  io_diffCommits_info_201_fpWen;
        input  io_diffCommits_info_201_vecWen;
        input  io_diffCommits_info_201_v0Wen;
        input  io_diffCommits_info_201_vlWen;
        input  io_diffCommits_info_202_ldest;
        input  io_diffCommits_info_202_pdest;
        input  io_diffCommits_info_202_rfWen;
        input  io_diffCommits_info_202_fpWen;
        input  io_diffCommits_info_202_vecWen;
        input  io_diffCommits_info_202_v0Wen;
        input  io_diffCommits_info_202_vlWen;
        input  io_diffCommits_info_203_ldest;
        input  io_diffCommits_info_203_pdest;
        input  io_diffCommits_info_203_rfWen;
        input  io_diffCommits_info_203_fpWen;
        input  io_diffCommits_info_203_vecWen;
        input  io_diffCommits_info_203_v0Wen;
        input  io_diffCommits_info_203_vlWen;
        input  io_diffCommits_info_204_ldest;
        input  io_diffCommits_info_204_pdest;
        input  io_diffCommits_info_204_rfWen;
        input  io_diffCommits_info_204_fpWen;
        input  io_diffCommits_info_204_vecWen;
        input  io_diffCommits_info_204_v0Wen;
        input  io_diffCommits_info_204_vlWen;
        input  io_diffCommits_info_205_ldest;
        input  io_diffCommits_info_205_pdest;
        input  io_diffCommits_info_205_rfWen;
        input  io_diffCommits_info_205_fpWen;
        input  io_diffCommits_info_205_vecWen;
        input  io_diffCommits_info_205_v0Wen;
        input  io_diffCommits_info_205_vlWen;
        input  io_diffCommits_info_206_ldest;
        input  io_diffCommits_info_206_pdest;
        input  io_diffCommits_info_206_rfWen;
        input  io_diffCommits_info_206_fpWen;
        input  io_diffCommits_info_206_vecWen;
        input  io_diffCommits_info_206_v0Wen;
        input  io_diffCommits_info_206_vlWen;
        input  io_diffCommits_info_207_ldest;
        input  io_diffCommits_info_207_pdest;
        input  io_diffCommits_info_207_rfWen;
        input  io_diffCommits_info_207_fpWen;
        input  io_diffCommits_info_207_vecWen;
        input  io_diffCommits_info_207_v0Wen;
        input  io_diffCommits_info_207_vlWen;
        input  io_diffCommits_info_208_ldest;
        input  io_diffCommits_info_208_pdest;
        input  io_diffCommits_info_208_rfWen;
        input  io_diffCommits_info_208_fpWen;
        input  io_diffCommits_info_208_vecWen;
        input  io_diffCommits_info_208_v0Wen;
        input  io_diffCommits_info_208_vlWen;
        input  io_diffCommits_info_209_ldest;
        input  io_diffCommits_info_209_pdest;
        input  io_diffCommits_info_209_rfWen;
        input  io_diffCommits_info_209_fpWen;
        input  io_diffCommits_info_209_vecWen;
        input  io_diffCommits_info_209_v0Wen;
        input  io_diffCommits_info_209_vlWen;
        input  io_diffCommits_info_210_ldest;
        input  io_diffCommits_info_210_pdest;
        input  io_diffCommits_info_210_rfWen;
        input  io_diffCommits_info_210_fpWen;
        input  io_diffCommits_info_210_vecWen;
        input  io_diffCommits_info_210_v0Wen;
        input  io_diffCommits_info_210_vlWen;
        input  io_diffCommits_info_211_ldest;
        input  io_diffCommits_info_211_pdest;
        input  io_diffCommits_info_211_rfWen;
        input  io_diffCommits_info_211_fpWen;
        input  io_diffCommits_info_211_vecWen;
        input  io_diffCommits_info_211_v0Wen;
        input  io_diffCommits_info_211_vlWen;
        input  io_diffCommits_info_212_ldest;
        input  io_diffCommits_info_212_pdest;
        input  io_diffCommits_info_212_rfWen;
        input  io_diffCommits_info_212_fpWen;
        input  io_diffCommits_info_212_vecWen;
        input  io_diffCommits_info_212_v0Wen;
        input  io_diffCommits_info_212_vlWen;
        input  io_diffCommits_info_213_ldest;
        input  io_diffCommits_info_213_pdest;
        input  io_diffCommits_info_213_rfWen;
        input  io_diffCommits_info_213_fpWen;
        input  io_diffCommits_info_213_vecWen;
        input  io_diffCommits_info_213_v0Wen;
        input  io_diffCommits_info_213_vlWen;
        input  io_diffCommits_info_214_ldest;
        input  io_diffCommits_info_214_pdest;
        input  io_diffCommits_info_214_rfWen;
        input  io_diffCommits_info_214_fpWen;
        input  io_diffCommits_info_214_vecWen;
        input  io_diffCommits_info_214_v0Wen;
        input  io_diffCommits_info_214_vlWen;
        input  io_diffCommits_info_215_ldest;
        input  io_diffCommits_info_215_pdest;
        input  io_diffCommits_info_215_rfWen;
        input  io_diffCommits_info_215_fpWen;
        input  io_diffCommits_info_215_vecWen;
        input  io_diffCommits_info_215_v0Wen;
        input  io_diffCommits_info_215_vlWen;
        input  io_diffCommits_info_216_ldest;
        input  io_diffCommits_info_216_pdest;
        input  io_diffCommits_info_216_rfWen;
        input  io_diffCommits_info_216_fpWen;
        input  io_diffCommits_info_216_vecWen;
        input  io_diffCommits_info_216_v0Wen;
        input  io_diffCommits_info_216_vlWen;
        input  io_diffCommits_info_217_ldest;
        input  io_diffCommits_info_217_pdest;
        input  io_diffCommits_info_217_rfWen;
        input  io_diffCommits_info_217_fpWen;
        input  io_diffCommits_info_217_vecWen;
        input  io_diffCommits_info_217_v0Wen;
        input  io_diffCommits_info_217_vlWen;
        input  io_diffCommits_info_218_ldest;
        input  io_diffCommits_info_218_pdest;
        input  io_diffCommits_info_218_rfWen;
        input  io_diffCommits_info_218_fpWen;
        input  io_diffCommits_info_218_vecWen;
        input  io_diffCommits_info_218_v0Wen;
        input  io_diffCommits_info_218_vlWen;
        input  io_diffCommits_info_219_ldest;
        input  io_diffCommits_info_219_pdest;
        input  io_diffCommits_info_219_rfWen;
        input  io_diffCommits_info_219_fpWen;
        input  io_diffCommits_info_219_vecWen;
        input  io_diffCommits_info_219_v0Wen;
        input  io_diffCommits_info_219_vlWen;
        input  io_diffCommits_info_220_ldest;
        input  io_diffCommits_info_220_pdest;
        input  io_diffCommits_info_220_rfWen;
        input  io_diffCommits_info_220_fpWen;
        input  io_diffCommits_info_220_vecWen;
        input  io_diffCommits_info_220_v0Wen;
        input  io_diffCommits_info_220_vlWen;
        input  io_diffCommits_info_221_ldest;
        input  io_diffCommits_info_221_pdest;
        input  io_diffCommits_info_221_rfWen;
        input  io_diffCommits_info_221_fpWen;
        input  io_diffCommits_info_221_vecWen;
        input  io_diffCommits_info_221_v0Wen;
        input  io_diffCommits_info_221_vlWen;
        input  io_diffCommits_info_222_ldest;
        input  io_diffCommits_info_222_pdest;
        input  io_diffCommits_info_222_rfWen;
        input  io_diffCommits_info_222_fpWen;
        input  io_diffCommits_info_222_vecWen;
        input  io_diffCommits_info_222_v0Wen;
        input  io_diffCommits_info_222_vlWen;
        input  io_diffCommits_info_223_ldest;
        input  io_diffCommits_info_223_pdest;
        input  io_diffCommits_info_223_rfWen;
        input  io_diffCommits_info_223_fpWen;
        input  io_diffCommits_info_223_vecWen;
        input  io_diffCommits_info_223_v0Wen;
        input  io_diffCommits_info_223_vlWen;
        input  io_diffCommits_info_224_ldest;
        input  io_diffCommits_info_224_pdest;
        input  io_diffCommits_info_224_rfWen;
        input  io_diffCommits_info_224_fpWen;
        input  io_diffCommits_info_224_vecWen;
        input  io_diffCommits_info_224_v0Wen;
        input  io_diffCommits_info_224_vlWen;
        input  io_diffCommits_info_225_ldest;
        input  io_diffCommits_info_225_pdest;
        input  io_diffCommits_info_225_rfWen;
        input  io_diffCommits_info_225_fpWen;
        input  io_diffCommits_info_225_vecWen;
        input  io_diffCommits_info_225_v0Wen;
        input  io_diffCommits_info_225_vlWen;
        input  io_diffCommits_info_226_ldest;
        input  io_diffCommits_info_226_pdest;
        input  io_diffCommits_info_226_rfWen;
        input  io_diffCommits_info_226_fpWen;
        input  io_diffCommits_info_226_vecWen;
        input  io_diffCommits_info_226_v0Wen;
        input  io_diffCommits_info_226_vlWen;
        input  io_diffCommits_info_227_ldest;
        input  io_diffCommits_info_227_pdest;
        input  io_diffCommits_info_227_rfWen;
        input  io_diffCommits_info_227_fpWen;
        input  io_diffCommits_info_227_vecWen;
        input  io_diffCommits_info_227_v0Wen;
        input  io_diffCommits_info_227_vlWen;
        input  io_diffCommits_info_228_ldest;
        input  io_diffCommits_info_228_pdest;
        input  io_diffCommits_info_228_rfWen;
        input  io_diffCommits_info_228_fpWen;
        input  io_diffCommits_info_228_vecWen;
        input  io_diffCommits_info_228_v0Wen;
        input  io_diffCommits_info_228_vlWen;
        input  io_diffCommits_info_229_ldest;
        input  io_diffCommits_info_229_pdest;
        input  io_diffCommits_info_229_rfWen;
        input  io_diffCommits_info_229_fpWen;
        input  io_diffCommits_info_229_vecWen;
        input  io_diffCommits_info_229_v0Wen;
        input  io_diffCommits_info_229_vlWen;
        input  io_diffCommits_info_230_ldest;
        input  io_diffCommits_info_230_pdest;
        input  io_diffCommits_info_230_rfWen;
        input  io_diffCommits_info_230_fpWen;
        input  io_diffCommits_info_230_vecWen;
        input  io_diffCommits_info_230_v0Wen;
        input  io_diffCommits_info_230_vlWen;
        input  io_diffCommits_info_231_ldest;
        input  io_diffCommits_info_231_pdest;
        input  io_diffCommits_info_231_rfWen;
        input  io_diffCommits_info_231_fpWen;
        input  io_diffCommits_info_231_vecWen;
        input  io_diffCommits_info_231_v0Wen;
        input  io_diffCommits_info_231_vlWen;
        input  io_diffCommits_info_232_ldest;
        input  io_diffCommits_info_232_pdest;
        input  io_diffCommits_info_232_rfWen;
        input  io_diffCommits_info_232_fpWen;
        input  io_diffCommits_info_232_vecWen;
        input  io_diffCommits_info_232_v0Wen;
        input  io_diffCommits_info_232_vlWen;
        input  io_diffCommits_info_233_ldest;
        input  io_diffCommits_info_233_pdest;
        input  io_diffCommits_info_233_rfWen;
        input  io_diffCommits_info_233_fpWen;
        input  io_diffCommits_info_233_vecWen;
        input  io_diffCommits_info_233_v0Wen;
        input  io_diffCommits_info_233_vlWen;
        input  io_diffCommits_info_234_ldest;
        input  io_diffCommits_info_234_pdest;
        input  io_diffCommits_info_234_rfWen;
        input  io_diffCommits_info_234_fpWen;
        input  io_diffCommits_info_234_vecWen;
        input  io_diffCommits_info_234_v0Wen;
        input  io_diffCommits_info_234_vlWen;
        input  io_diffCommits_info_235_ldest;
        input  io_diffCommits_info_235_pdest;
        input  io_diffCommits_info_235_rfWen;
        input  io_diffCommits_info_235_fpWen;
        input  io_diffCommits_info_235_vecWen;
        input  io_diffCommits_info_235_v0Wen;
        input  io_diffCommits_info_235_vlWen;
        input  io_diffCommits_info_236_ldest;
        input  io_diffCommits_info_236_pdest;
        input  io_diffCommits_info_236_rfWen;
        input  io_diffCommits_info_236_fpWen;
        input  io_diffCommits_info_236_vecWen;
        input  io_diffCommits_info_236_v0Wen;
        input  io_diffCommits_info_236_vlWen;
        input  io_diffCommits_info_237_ldest;
        input  io_diffCommits_info_237_pdest;
        input  io_diffCommits_info_237_rfWen;
        input  io_diffCommits_info_237_fpWen;
        input  io_diffCommits_info_237_vecWen;
        input  io_diffCommits_info_237_v0Wen;
        input  io_diffCommits_info_237_vlWen;
        input  io_diffCommits_info_238_ldest;
        input  io_diffCommits_info_238_pdest;
        input  io_diffCommits_info_238_rfWen;
        input  io_diffCommits_info_238_fpWen;
        input  io_diffCommits_info_238_vecWen;
        input  io_diffCommits_info_238_v0Wen;
        input  io_diffCommits_info_238_vlWen;
        input  io_diffCommits_info_239_ldest;
        input  io_diffCommits_info_239_pdest;
        input  io_diffCommits_info_239_rfWen;
        input  io_diffCommits_info_239_fpWen;
        input  io_diffCommits_info_239_vecWen;
        input  io_diffCommits_info_239_v0Wen;
        input  io_diffCommits_info_239_vlWen;
        input  io_diffCommits_info_240_ldest;
        input  io_diffCommits_info_240_pdest;
        input  io_diffCommits_info_240_rfWen;
        input  io_diffCommits_info_240_fpWen;
        input  io_diffCommits_info_240_vecWen;
        input  io_diffCommits_info_240_v0Wen;
        input  io_diffCommits_info_240_vlWen;
        input  io_diffCommits_info_241_ldest;
        input  io_diffCommits_info_241_pdest;
        input  io_diffCommits_info_241_rfWen;
        input  io_diffCommits_info_241_fpWen;
        input  io_diffCommits_info_241_vecWen;
        input  io_diffCommits_info_241_v0Wen;
        input  io_diffCommits_info_241_vlWen;
        input  io_diffCommits_info_242_ldest;
        input  io_diffCommits_info_242_pdest;
        input  io_diffCommits_info_242_rfWen;
        input  io_diffCommits_info_242_fpWen;
        input  io_diffCommits_info_242_vecWen;
        input  io_diffCommits_info_242_v0Wen;
        input  io_diffCommits_info_242_vlWen;
        input  io_diffCommits_info_243_ldest;
        input  io_diffCommits_info_243_pdest;
        input  io_diffCommits_info_243_rfWen;
        input  io_diffCommits_info_243_fpWen;
        input  io_diffCommits_info_243_vecWen;
        input  io_diffCommits_info_243_v0Wen;
        input  io_diffCommits_info_243_vlWen;
        input  io_diffCommits_info_244_ldest;
        input  io_diffCommits_info_244_pdest;
        input  io_diffCommits_info_244_rfWen;
        input  io_diffCommits_info_244_fpWen;
        input  io_diffCommits_info_244_vecWen;
        input  io_diffCommits_info_244_v0Wen;
        input  io_diffCommits_info_244_vlWen;
        input  io_diffCommits_info_245_ldest;
        input  io_diffCommits_info_245_pdest;
        input  io_diffCommits_info_245_rfWen;
        input  io_diffCommits_info_245_fpWen;
        input  io_diffCommits_info_245_vecWen;
        input  io_diffCommits_info_245_v0Wen;
        input  io_diffCommits_info_245_vlWen;
        input  io_diffCommits_info_246_ldest;
        input  io_diffCommits_info_246_pdest;
        input  io_diffCommits_info_246_rfWen;
        input  io_diffCommits_info_246_fpWen;
        input  io_diffCommits_info_246_vecWen;
        input  io_diffCommits_info_246_v0Wen;
        input  io_diffCommits_info_246_vlWen;
        input  io_diffCommits_info_247_ldest;
        input  io_diffCommits_info_247_pdest;
        input  io_diffCommits_info_247_rfWen;
        input  io_diffCommits_info_247_fpWen;
        input  io_diffCommits_info_247_vecWen;
        input  io_diffCommits_info_247_v0Wen;
        input  io_diffCommits_info_247_vlWen;
        input  io_diffCommits_info_248_ldest;
        input  io_diffCommits_info_248_pdest;
        input  io_diffCommits_info_248_rfWen;
        input  io_diffCommits_info_248_fpWen;
        input  io_diffCommits_info_248_vecWen;
        input  io_diffCommits_info_248_v0Wen;
        input  io_diffCommits_info_248_vlWen;
        input  io_diffCommits_info_249_ldest;
        input  io_diffCommits_info_249_pdest;
        input  io_diffCommits_info_249_rfWen;
        input  io_diffCommits_info_249_fpWen;
        input  io_diffCommits_info_249_vecWen;
        input  io_diffCommits_info_249_v0Wen;
        input  io_diffCommits_info_249_vlWen;
        input  io_diffCommits_info_250_ldest;
        input  io_diffCommits_info_250_pdest;
        input  io_diffCommits_info_250_rfWen;
        input  io_diffCommits_info_250_fpWen;
        input  io_diffCommits_info_250_vecWen;
        input  io_diffCommits_info_250_v0Wen;
        input  io_diffCommits_info_250_vlWen;
        input  io_diffCommits_info_251_ldest;
        input  io_diffCommits_info_251_pdest;
        input  io_diffCommits_info_251_rfWen;
        input  io_diffCommits_info_251_fpWen;
        input  io_diffCommits_info_251_vecWen;
        input  io_diffCommits_info_251_v0Wen;
        input  io_diffCommits_info_251_vlWen;
        input  io_diffCommits_info_252_ldest;
        input  io_diffCommits_info_252_pdest;
        input  io_diffCommits_info_252_rfWen;
        input  io_diffCommits_info_252_fpWen;
        input  io_diffCommits_info_252_vecWen;
        input  io_diffCommits_info_252_v0Wen;
        input  io_diffCommits_info_252_vlWen;
        input  io_diffCommits_info_253_ldest;
        input  io_diffCommits_info_253_pdest;
        input  io_diffCommits_info_253_rfWen;
        input  io_diffCommits_info_253_fpWen;
        input  io_diffCommits_info_253_vecWen;
        input  io_diffCommits_info_253_v0Wen;
        input  io_diffCommits_info_253_vlWen;
        input  io_diffCommits_info_254_ldest;
        input  io_diffCommits_info_254_pdest;
        input  io_diffCommits_info_254_rfWen;
        input  io_diffCommits_info_254_fpWen;
        input  io_diffCommits_info_254_vecWen;
        input  io_diffCommits_info_254_v0Wen;
        input  io_diffCommits_info_254_vlWen;
        input  io_diffCommits_info_255_ldest;
        input  io_diffCommits_info_255_pdest;
        input  io_diffCommits_info_256_ldest;
        input  io_diffCommits_info_256_pdest;
        input  io_diffCommits_info_257_ldest;
        input  io_diffCommits_info_257_pdest;
        input  io_diffCommits_info_258_ldest;
        input  io_diffCommits_info_258_pdest;
        input  io_diffCommits_info_259_ldest;
        input  io_diffCommits_info_259_pdest;
        input  io_diffCommits_info_260_ldest;
        input  io_diffCommits_info_260_pdest;
        input  io_diffCommits_info_261_ldest;
        input  io_diffCommits_info_261_pdest;
        input  io_diffCommits_info_262_ldest;
        input  io_diffCommits_info_262_pdest;
        input  io_diffCommits_info_263_ldest;
        input  io_diffCommits_info_263_pdest;
        input  io_diffCommits_info_264_ldest;
        input  io_diffCommits_info_264_pdest;
        input  io_diffCommits_info_265_ldest;
        input  io_diffCommits_info_265_pdest;
        input  io_diffCommits_info_266_ldest;
        input  io_diffCommits_info_266_pdest;
        input  io_diffCommits_info_267_ldest;
        input  io_diffCommits_info_267_pdest;
        input  io_diffCommits_info_268_ldest;
        input  io_diffCommits_info_268_pdest;
        input  io_diffCommits_info_269_ldest;
        input  io_diffCommits_info_269_pdest;
        input  io_diffCommits_info_270_ldest;
        input  io_diffCommits_info_270_pdest;
        input  io_diffCommits_info_271_ldest;
        input  io_diffCommits_info_271_pdest;
        input  io_diffCommits_info_272_ldest;
        input  io_diffCommits_info_272_pdest;
        input  io_diffCommits_info_273_ldest;
        input  io_diffCommits_info_273_pdest;
        input  io_diffCommits_info_274_ldest;
        input  io_diffCommits_info_274_pdest;
        input  io_diffCommits_info_275_ldest;
        input  io_diffCommits_info_275_pdest;
        input  io_diffCommits_info_276_ldest;
        input  io_diffCommits_info_276_pdest;
        input  io_diffCommits_info_277_ldest;
        input  io_diffCommits_info_277_pdest;
        input  io_diffCommits_info_278_ldest;
        input  io_diffCommits_info_278_pdest;
        input  io_diffCommits_info_279_ldest;
        input  io_diffCommits_info_279_pdest;
        input  io_diffCommits_info_280_ldest;
        input  io_diffCommits_info_280_pdest;
        input  io_diffCommits_info_281_ldest;
        input  io_diffCommits_info_281_pdest;
        input  io_diffCommits_info_282_ldest;
        input  io_diffCommits_info_282_pdest;
        input  io_diffCommits_info_283_ldest;
        input  io_diffCommits_info_283_pdest;
        input  io_diffCommits_info_284_ldest;
        input  io_diffCommits_info_284_pdest;
        input  io_diffCommits_info_285_ldest;
        input  io_diffCommits_info_285_pdest;
        input  io_diffCommits_info_286_ldest;
        input  io_diffCommits_info_286_pdest;
        input  io_diffCommits_info_287_ldest;
        input  io_diffCommits_info_287_pdest;
        input  io_diffCommits_info_288_ldest;
        input  io_diffCommits_info_288_pdest;
        input  io_diffCommits_info_289_ldest;
        input  io_diffCommits_info_289_pdest;
        input  io_diffCommits_info_290_ldest;
        input  io_diffCommits_info_290_pdest;
        input  io_diffCommits_info_291_ldest;
        input  io_diffCommits_info_291_pdest;
        input  io_diffCommits_info_292_ldest;
        input  io_diffCommits_info_292_pdest;
        input  io_diffCommits_info_293_ldest;
        input  io_diffCommits_info_293_pdest;
        input  io_diffCommits_info_294_ldest;
        input  io_diffCommits_info_294_pdest;
        input  io_diffCommits_info_295_ldest;
        input  io_diffCommits_info_295_pdest;
        input  io_diffCommits_info_296_ldest;
        input  io_diffCommits_info_296_pdest;
        input  io_diffCommits_info_297_ldest;
        input  io_diffCommits_info_297_pdest;
        input  io_diffCommits_info_298_ldest;
        input  io_diffCommits_info_298_pdest;
        input  io_diffCommits_info_299_ldest;
        input  io_diffCommits_info_299_pdest;
        input  io_diffCommits_info_300_ldest;
        input  io_diffCommits_info_300_pdest;
        input  io_diffCommits_info_301_ldest;
        input  io_diffCommits_info_301_pdest;
        input  io_diffCommits_info_302_ldest;
        input  io_diffCommits_info_302_pdest;
        input  io_diffCommits_info_303_ldest;
        input  io_diffCommits_info_303_pdest;
        input  io_diffCommits_info_304_ldest;
        input  io_diffCommits_info_304_pdest;
        input  io_diffCommits_info_305_ldest;
        input  io_diffCommits_info_305_pdest;
        input  io_diffCommits_info_306_ldest;
        input  io_diffCommits_info_306_pdest;
        input  io_diffCommits_info_307_ldest;
        input  io_diffCommits_info_307_pdest;
        input  io_diffCommits_info_308_ldest;
        input  io_diffCommits_info_308_pdest;
        input  io_diffCommits_info_309_ldest;
        input  io_diffCommits_info_309_pdest;
        input  io_diffCommits_info_310_ldest;
        input  io_diffCommits_info_310_pdest;
        input  io_diffCommits_info_311_ldest;
        input  io_diffCommits_info_311_pdest;
        input  io_diffCommits_info_312_ldest;
        input  io_diffCommits_info_312_pdest;
        input  io_diffCommits_info_313_ldest;
        input  io_diffCommits_info_313_pdest;
        input  io_diffCommits_info_314_ldest;
        input  io_diffCommits_info_314_pdest;
        input  io_diffCommits_info_315_ldest;
        input  io_diffCommits_info_315_pdest;
        input  io_diffCommits_info_316_ldest;
        input  io_diffCommits_info_316_pdest;
        input  io_diffCommits_info_317_ldest;
        input  io_diffCommits_info_317_pdest;
        input  io_diffCommits_info_318_ldest;
        input  io_diffCommits_info_318_pdest;
        input  io_diffCommits_info_319_ldest;
        input  io_diffCommits_info_319_pdest;
        input  io_diffCommits_info_320_ldest;
        input  io_diffCommits_info_320_pdest;
        input  io_diffCommits_info_321_ldest;
        input  io_diffCommits_info_321_pdest;
        input  io_diffCommits_info_322_ldest;
        input  io_diffCommits_info_322_pdest;
        input  io_diffCommits_info_323_ldest;
        input  io_diffCommits_info_323_pdest;
        input  io_diffCommits_info_324_ldest;
        input  io_diffCommits_info_324_pdest;
        input  io_diffCommits_info_325_ldest;
        input  io_diffCommits_info_325_pdest;
        input  io_diffCommits_info_326_ldest;
        input  io_diffCommits_info_326_pdest;
        input  io_diffCommits_info_327_ldest;
        input  io_diffCommits_info_327_pdest;
        input  io_diffCommits_info_328_ldest;
        input  io_diffCommits_info_328_pdest;
        input  io_diffCommits_info_329_ldest;
        input  io_diffCommits_info_329_pdest;
        input  io_diffCommits_info_330_ldest;
        input  io_diffCommits_info_330_pdest;
        input  io_diffCommits_info_331_ldest;
        input  io_diffCommits_info_331_pdest;
        input  io_diffCommits_info_332_ldest;
        input  io_diffCommits_info_332_pdest;
        input  io_diffCommits_info_333_ldest;
        input  io_diffCommits_info_333_pdest;
        input  io_diffCommits_info_334_ldest;
        input  io_diffCommits_info_334_pdest;
        input  io_diffCommits_info_335_ldest;
        input  io_diffCommits_info_335_pdest;
        input  io_diffCommits_info_336_ldest;
        input  io_diffCommits_info_336_pdest;
        input  io_diffCommits_info_337_ldest;
        input  io_diffCommits_info_337_pdest;
        input  io_diffCommits_info_338_ldest;
        input  io_diffCommits_info_338_pdest;
        input  io_diffCommits_info_339_ldest;
        input  io_diffCommits_info_339_pdest;
        input  io_diffCommits_info_340_ldest;
        input  io_diffCommits_info_340_pdest;
        input  io_diffCommits_info_341_ldest;
        input  io_diffCommits_info_341_pdest;
        input  io_diffCommits_info_342_ldest;
        input  io_diffCommits_info_342_pdest;
        input  io_diffCommits_info_343_ldest;
        input  io_diffCommits_info_343_pdest;
        input  io_diffCommits_info_344_ldest;
        input  io_diffCommits_info_344_pdest;
        input  io_diffCommits_info_345_ldest;
        input  io_diffCommits_info_345_pdest;
        input  io_diffCommits_info_346_ldest;
        input  io_diffCommits_info_346_pdest;
        input  io_diffCommits_info_347_ldest;
        input  io_diffCommits_info_347_pdest;
        input  io_diffCommits_info_348_ldest;
        input  io_diffCommits_info_348_pdest;
        input  io_diffCommits_info_349_ldest;
        input  io_diffCommits_info_349_pdest;
        input  io_diffCommits_info_350_ldest;
        input  io_diffCommits_info_350_pdest;
        input  io_diffCommits_info_351_ldest;
        input  io_diffCommits_info_351_pdest;
        input  io_diffCommits_info_352_ldest;
        input  io_diffCommits_info_352_pdest;
        input  io_diffCommits_info_353_ldest;
        input  io_diffCommits_info_353_pdest;
        input  io_diffCommits_info_354_ldest;
        input  io_diffCommits_info_354_pdest;
        input  io_diffCommits_info_355_ldest;
        input  io_diffCommits_info_355_pdest;
        input  io_diffCommits_info_356_ldest;
        input  io_diffCommits_info_356_pdest;
        input  io_diffCommits_info_357_ldest;
        input  io_diffCommits_info_357_pdest;
        input  io_diffCommits_info_358_ldest;
        input  io_diffCommits_info_358_pdest;
        input  io_diffCommits_info_359_ldest;
        input  io_diffCommits_info_359_pdest;
        input  io_diffCommits_info_360_ldest;
        input  io_diffCommits_info_360_pdest;
        input  io_diffCommits_info_361_ldest;
        input  io_diffCommits_info_361_pdest;
        input  io_diffCommits_info_362_ldest;
        input  io_diffCommits_info_362_pdest;
        input  io_diffCommits_info_363_ldest;
        input  io_diffCommits_info_363_pdest;
        input  io_diffCommits_info_364_ldest;
        input  io_diffCommits_info_364_pdest;
        input  io_diffCommits_info_365_ldest;
        input  io_diffCommits_info_365_pdest;
        input  io_diffCommits_info_366_ldest;
        input  io_diffCommits_info_366_pdest;
        input  io_diffCommits_info_367_ldest;
        input  io_diffCommits_info_367_pdest;
        input  io_diffCommits_info_368_ldest;
        input  io_diffCommits_info_368_pdest;
        input  io_diffCommits_info_369_ldest;
        input  io_diffCommits_info_369_pdest;
        input  io_diffCommits_info_370_ldest;
        input  io_diffCommits_info_370_pdest;
        input  io_diffCommits_info_371_ldest;
        input  io_diffCommits_info_371_pdest;
        input  io_diffCommits_info_372_ldest;
        input  io_diffCommits_info_372_pdest;
        input  io_diffCommits_info_373_ldest;
        input  io_diffCommits_info_373_pdest;
        input  io_diffCommits_info_374_ldest;
        input  io_diffCommits_info_374_pdest;
        input  io_diffCommits_info_375_ldest;
        input  io_diffCommits_info_375_pdest;
        input  io_diffCommits_info_376_ldest;
        input  io_diffCommits_info_376_pdest;
        input  io_diffCommits_info_377_ldest;
        input  io_diffCommits_info_377_pdest;
        input  io_diffCommits_info_378_ldest;
        input  io_diffCommits_info_378_pdest;
        input  io_diffCommits_info_379_ldest;
        input  io_diffCommits_info_379_pdest;
        input  io_diffCommits_info_380_ldest;
        input  io_diffCommits_info_380_pdest;
        input  io_diffCommits_info_381_ldest;
        input  io_diffCommits_info_381_pdest;
        input  io_diffCommits_info_382_ldest;
        input  io_diffCommits_info_382_pdest;
        input  io_diffCommits_info_383_ldest;
        input  io_diffCommits_info_383_pdest;
        input  io_diffCommits_info_384_ldest;
        input  io_diffCommits_info_384_pdest;
        input  io_diffCommits_info_385_ldest;
        input  io_diffCommits_info_385_pdest;
        input  io_diffCommits_info_386_ldest;
        input  io_diffCommits_info_386_pdest;
        input  io_diffCommits_info_387_ldest;
        input  io_diffCommits_info_387_pdest;
        input  io_diffCommits_info_388_ldest;
        input  io_diffCommits_info_388_pdest;
        input  io_diffCommits_info_389_ldest;
        input  io_diffCommits_info_389_pdest;
        input  io_lsq_scommit;
        input  io_lsq_pendingMMIOld;
        input  io_lsq_pendingst;
        input  io_lsq_pendingPtr_flag;
        input  io_lsq_pendingPtr_value;
        input  io_robDeqPtr_flag;
        input  io_robDeqPtr_value;
        input  io_csr_fflags_valid;
        input  io_csr_fflags_bits;
        input  io_csr_vxsat_valid;
        input  io_csr_vxsat_bits;
        input  io_csr_vstart_valid;
        input  io_csr_vstart_bits;
        input  io_csr_dirty_fs;
        input  io_csr_dirty_vs;
        input  io_csr_perfinfo_retiredInstr;
        input  io_cpu_halt;
        input  io_wfi_wfiReq;
        input  io_toDecode_isResumeVType;
        input  io_toDecode_walkToArchVType;
        input  io_toDecode_walkVType_valid;
        input  io_toDecode_walkVType_bits_illegal;
        input  io_toDecode_walkVType_bits_vma;
        input  io_toDecode_walkVType_bits_vta;
        input  io_toDecode_walkVType_bits_vsew;
        input  io_toDecode_walkVType_bits_vlmul;
        input  io_toDecode_commitVType_vtype_valid;
        input  io_toDecode_commitVType_vtype_bits_illegal;
        input  io_toDecode_commitVType_vtype_bits_vma;
        input  io_toDecode_commitVType_vtype_bits_vta;
        input  io_toDecode_commitVType_vtype_bits_vsew;
        input  io_toDecode_commitVType_vtype_bits_vlmul;
        input  io_toDecode_commitVType_hasVsetvl;
        input  io_readGPAMemAddr_valid;
        input  io_readGPAMemAddr_bits_ftqPtr_value;
        input  io_readGPAMemAddr_bits_ftqOffset;
        input  io_toVecExcpMod_logicPhyRegMap_0_valid;
        input  io_toVecExcpMod_logicPhyRegMap_0_bits_lreg;
        input  io_toVecExcpMod_logicPhyRegMap_0_bits_preg;
        input  io_toVecExcpMod_logicPhyRegMap_1_valid;
        input  io_toVecExcpMod_logicPhyRegMap_1_bits_lreg;
        input  io_toVecExcpMod_logicPhyRegMap_1_bits_preg;
        input  io_toVecExcpMod_logicPhyRegMap_2_valid;
        input  io_toVecExcpMod_logicPhyRegMap_2_bits_lreg;
        input  io_toVecExcpMod_logicPhyRegMap_2_bits_preg;
        input  io_toVecExcpMod_logicPhyRegMap_3_valid;
        input  io_toVecExcpMod_logicPhyRegMap_3_bits_lreg;
        input  io_toVecExcpMod_logicPhyRegMap_3_bits_preg;
        input  io_toVecExcpMod_logicPhyRegMap_4_valid;
        input  io_toVecExcpMod_logicPhyRegMap_4_bits_lreg;
        input  io_toVecExcpMod_logicPhyRegMap_4_bits_preg;
        input  io_toVecExcpMod_logicPhyRegMap_5_valid;
        input  io_toVecExcpMod_logicPhyRegMap_5_bits_lreg;
        input  io_toVecExcpMod_logicPhyRegMap_5_bits_preg;
        input  io_toVecExcpMod_excpInfo_valid;
        input  io_toVecExcpMod_excpInfo_bits_vstart;
        input  io_toVecExcpMod_excpInfo_bits_vsew;
        input  io_toVecExcpMod_excpInfo_bits_veew;
        input  io_toVecExcpMod_excpInfo_bits_vlmul;
        input  io_toVecExcpMod_excpInfo_bits_nf;
        input  io_toVecExcpMod_excpInfo_bits_isStride;
        input  io_toVecExcpMod_excpInfo_bits_isIndexed;
        input  io_toVecExcpMod_excpInfo_bits_isWhole;
        input  io_toVecExcpMod_excpInfo_bits_isVlm;
        input  io_storeDebugInfo_1_pc;
        input  io_perf_0_value;
        input  io_perf_1_value;
        input  io_perf_2_value;
        input  io_perf_3_value;
        input  io_perf_4_value;
        input  io_perf_5_value;
        input  io_perf_6_value;
        input  io_perf_7_value;
        input  io_perf_8_value;
        input  io_perf_9_value;
        input  io_perf_10_value;
        input  io_perf_11_value;
        input  io_perf_12_value;
        input  io_perf_13_value;
        input  io_perf_14_value;
        input  io_perf_15_value;
        input  io_perf_16_value;
        input  io_perf_17_value;
        input  io_error_0;

    endclocking:drv_cb

    clocking mon_cb @(posedge clk);
        `ifdef INTERFACE_ADD_DELAY
            default input #`DEF_SETUP_TIME output #`DEF_HOLD_TIME;
        `endif
        input  io_enq_canAccept;
        input  io_enq_canAcceptForDispatch;
        input  io_enq_isEmpty;
        input  io_flushOut_valid;
        input  io_flushOut_bits_isRVC;
        input  io_flushOut_bits_robIdx_flag;
        input  io_flushOut_bits_robIdx_value;
        input  io_flushOut_bits_ftqIdx_flag;
        input  io_flushOut_bits_ftqIdx_value;
        input  io_flushOut_bits_ftqOffset;
        input  io_flushOut_bits_level;
        input  io_exception_valid;
        input  io_exception_bits_instr;
        input  io_exception_bits_commitType;
        input  io_exception_bits_exceptionVec_0;
        input  io_exception_bits_exceptionVec_1;
        input  io_exception_bits_exceptionVec_2;
        input  io_exception_bits_exceptionVec_3;
        input  io_exception_bits_exceptionVec_4;
        input  io_exception_bits_exceptionVec_5;
        input  io_exception_bits_exceptionVec_6;
        input  io_exception_bits_exceptionVec_7;
        input  io_exception_bits_exceptionVec_8;
        input  io_exception_bits_exceptionVec_9;
        input  io_exception_bits_exceptionVec_10;
        input  io_exception_bits_exceptionVec_11;
        input  io_exception_bits_exceptionVec_12;
        input  io_exception_bits_exceptionVec_13;
        input  io_exception_bits_exceptionVec_14;
        input  io_exception_bits_exceptionVec_15;
        input  io_exception_bits_exceptionVec_16;
        input  io_exception_bits_exceptionVec_17;
        input  io_exception_bits_exceptionVec_18;
        input  io_exception_bits_exceptionVec_19;
        input  io_exception_bits_exceptionVec_20;
        input  io_exception_bits_exceptionVec_21;
        input  io_exception_bits_exceptionVec_22;
        input  io_exception_bits_exceptionVec_23;
        input  io_exception_bits_isPcBkpt;
        input  io_exception_bits_isFetchMalAddr;
        input  io_exception_bits_gpaddr;
        input  io_exception_bits_singleStep;
        input  io_exception_bits_crossPageIPFFix;
        input  io_exception_bits_isInterrupt;
        input  io_exception_bits_isHls;
        input  io_exception_bits_trigger;
        input  io_exception_bits_isForVSnonLeafPTE;
        input  io_commits_isCommit;
        input  io_commits_commitValid_0;
        input  io_commits_commitValid_1;
        input  io_commits_commitValid_2;
        input  io_commits_commitValid_3;
        input  io_commits_commitValid_4;
        input  io_commits_commitValid_5;
        input  io_commits_commitValid_6;
        input  io_commits_commitValid_7;
        input  io_commits_isWalk;
        input  io_commits_walkValid_0;
        input  io_commits_walkValid_1;
        input  io_commits_walkValid_2;
        input  io_commits_walkValid_3;
        input  io_commits_walkValid_4;
        input  io_commits_walkValid_5;
        input  io_commits_walkValid_6;
        input  io_commits_walkValid_7;
        input  io_commits_info_0_walk_v;
        input  io_commits_info_0_commit_v;
        input  io_commits_info_0_commit_w;
        input  io_commits_info_0_realDestSize;
        input  io_commits_info_0_interrupt_safe;
        input  io_commits_info_0_wflags;
        input  io_commits_info_0_fflags;
        input  io_commits_info_0_vxsat;
        input  io_commits_info_0_isRVC;
        input  io_commits_info_0_isVset;
        input  io_commits_info_0_isHls;
        input  io_commits_info_0_isVls;
        input  io_commits_info_0_vls;
        input  io_commits_info_0_mmio;
        input  io_commits_info_0_commitType;
        input  io_commits_info_0_ftqIdx_flag;
        input  io_commits_info_0_ftqIdx_value;
        input  io_commits_info_0_ftqOffset;
        input  io_commits_info_0_instrSize;
        input  io_commits_info_0_fpWen;
        input  io_commits_info_0_rfWen;
        input  io_commits_info_0_needFlush;
        input  io_commits_info_0_traceBlockInPipe_itype;
        input  io_commits_info_0_traceBlockInPipe_iretire;
        input  io_commits_info_0_traceBlockInPipe_ilastsize;
        input  io_commits_info_0_debug_pc;
        input  io_commits_info_0_debug_instr;
        input  io_commits_info_0_debug_ldest;
        input  io_commits_info_0_debug_pdest;
        input  io_commits_info_0_debug_otherPdest_0;
        input  io_commits_info_0_debug_otherPdest_1;
        input  io_commits_info_0_debug_otherPdest_2;
        input  io_commits_info_0_debug_otherPdest_3;
        input  io_commits_info_0_debug_otherPdest_4;
        input  io_commits_info_0_debug_otherPdest_5;
        input  io_commits_info_0_debug_otherPdest_6;
        input  io_commits_info_0_debug_fuType;
        input  io_commits_info_0_dirtyFs;
        input  io_commits_info_0_dirtyVs;
        input  io_commits_info_1_walk_v;
        input  io_commits_info_1_commit_v;
        input  io_commits_info_1_commit_w;
        input  io_commits_info_1_realDestSize;
        input  io_commits_info_1_interrupt_safe;
        input  io_commits_info_1_wflags;
        input  io_commits_info_1_fflags;
        input  io_commits_info_1_vxsat;
        input  io_commits_info_1_isRVC;
        input  io_commits_info_1_isVset;
        input  io_commits_info_1_isHls;
        input  io_commits_info_1_isVls;
        input  io_commits_info_1_vls;
        input  io_commits_info_1_mmio;
        input  io_commits_info_1_commitType;
        input  io_commits_info_1_ftqIdx_flag;
        input  io_commits_info_1_ftqIdx_value;
        input  io_commits_info_1_ftqOffset;
        input  io_commits_info_1_instrSize;
        input  io_commits_info_1_fpWen;
        input  io_commits_info_1_rfWen;
        input  io_commits_info_1_needFlush;
        input  io_commits_info_1_traceBlockInPipe_itype;
        input  io_commits_info_1_traceBlockInPipe_iretire;
        input  io_commits_info_1_traceBlockInPipe_ilastsize;
        input  io_commits_info_1_debug_pc;
        input  io_commits_info_1_debug_instr;
        input  io_commits_info_1_debug_ldest;
        input  io_commits_info_1_debug_pdest;
        input  io_commits_info_1_debug_otherPdest_0;
        input  io_commits_info_1_debug_otherPdest_1;
        input  io_commits_info_1_debug_otherPdest_2;
        input  io_commits_info_1_debug_otherPdest_3;
        input  io_commits_info_1_debug_otherPdest_4;
        input  io_commits_info_1_debug_otherPdest_5;
        input  io_commits_info_1_debug_otherPdest_6;
        input  io_commits_info_1_debug_fuType;
        input  io_commits_info_1_dirtyFs;
        input  io_commits_info_1_dirtyVs;
        input  io_commits_info_2_walk_v;
        input  io_commits_info_2_commit_v;
        input  io_commits_info_2_commit_w;
        input  io_commits_info_2_realDestSize;
        input  io_commits_info_2_interrupt_safe;
        input  io_commits_info_2_wflags;
        input  io_commits_info_2_fflags;
        input  io_commits_info_2_vxsat;
        input  io_commits_info_2_isRVC;
        input  io_commits_info_2_isVset;
        input  io_commits_info_2_isHls;
        input  io_commits_info_2_isVls;
        input  io_commits_info_2_vls;
        input  io_commits_info_2_mmio;
        input  io_commits_info_2_commitType;
        input  io_commits_info_2_ftqIdx_flag;
        input  io_commits_info_2_ftqIdx_value;
        input  io_commits_info_2_ftqOffset;
        input  io_commits_info_2_instrSize;
        input  io_commits_info_2_fpWen;
        input  io_commits_info_2_rfWen;
        input  io_commits_info_2_needFlush;
        input  io_commits_info_2_traceBlockInPipe_itype;
        input  io_commits_info_2_traceBlockInPipe_iretire;
        input  io_commits_info_2_traceBlockInPipe_ilastsize;
        input  io_commits_info_2_debug_pc;
        input  io_commits_info_2_debug_instr;
        input  io_commits_info_2_debug_ldest;
        input  io_commits_info_2_debug_pdest;
        input  io_commits_info_2_debug_otherPdest_0;
        input  io_commits_info_2_debug_otherPdest_1;
        input  io_commits_info_2_debug_otherPdest_2;
        input  io_commits_info_2_debug_otherPdest_3;
        input  io_commits_info_2_debug_otherPdest_4;
        input  io_commits_info_2_debug_otherPdest_5;
        input  io_commits_info_2_debug_otherPdest_6;
        input  io_commits_info_2_debug_fuType;
        input  io_commits_info_2_dirtyFs;
        input  io_commits_info_2_dirtyVs;
        input  io_commits_info_3_walk_v;
        input  io_commits_info_3_commit_v;
        input  io_commits_info_3_commit_w;
        input  io_commits_info_3_realDestSize;
        input  io_commits_info_3_interrupt_safe;
        input  io_commits_info_3_wflags;
        input  io_commits_info_3_fflags;
        input  io_commits_info_3_vxsat;
        input  io_commits_info_3_isRVC;
        input  io_commits_info_3_isVset;
        input  io_commits_info_3_isHls;
        input  io_commits_info_3_isVls;
        input  io_commits_info_3_vls;
        input  io_commits_info_3_mmio;
        input  io_commits_info_3_commitType;
        input  io_commits_info_3_ftqIdx_flag;
        input  io_commits_info_3_ftqIdx_value;
        input  io_commits_info_3_ftqOffset;
        input  io_commits_info_3_instrSize;
        input  io_commits_info_3_fpWen;
        input  io_commits_info_3_rfWen;
        input  io_commits_info_3_needFlush;
        input  io_commits_info_3_traceBlockInPipe_itype;
        input  io_commits_info_3_traceBlockInPipe_iretire;
        input  io_commits_info_3_traceBlockInPipe_ilastsize;
        input  io_commits_info_3_debug_pc;
        input  io_commits_info_3_debug_instr;
        input  io_commits_info_3_debug_ldest;
        input  io_commits_info_3_debug_pdest;
        input  io_commits_info_3_debug_otherPdest_0;
        input  io_commits_info_3_debug_otherPdest_1;
        input  io_commits_info_3_debug_otherPdest_2;
        input  io_commits_info_3_debug_otherPdest_3;
        input  io_commits_info_3_debug_otherPdest_4;
        input  io_commits_info_3_debug_otherPdest_5;
        input  io_commits_info_3_debug_otherPdest_6;
        input  io_commits_info_3_debug_fuType;
        input  io_commits_info_3_dirtyFs;
        input  io_commits_info_3_dirtyVs;
        input  io_commits_info_4_walk_v;
        input  io_commits_info_4_commit_v;
        input  io_commits_info_4_commit_w;
        input  io_commits_info_4_realDestSize;
        input  io_commits_info_4_interrupt_safe;
        input  io_commits_info_4_wflags;
        input  io_commits_info_4_fflags;
        input  io_commits_info_4_vxsat;
        input  io_commits_info_4_isRVC;
        input  io_commits_info_4_isVset;
        input  io_commits_info_4_isHls;
        input  io_commits_info_4_isVls;
        input  io_commits_info_4_vls;
        input  io_commits_info_4_mmio;
        input  io_commits_info_4_commitType;
        input  io_commits_info_4_ftqIdx_flag;
        input  io_commits_info_4_ftqIdx_value;
        input  io_commits_info_4_ftqOffset;
        input  io_commits_info_4_instrSize;
        input  io_commits_info_4_fpWen;
        input  io_commits_info_4_rfWen;
        input  io_commits_info_4_needFlush;
        input  io_commits_info_4_traceBlockInPipe_itype;
        input  io_commits_info_4_traceBlockInPipe_iretire;
        input  io_commits_info_4_traceBlockInPipe_ilastsize;
        input  io_commits_info_4_debug_pc;
        input  io_commits_info_4_debug_instr;
        input  io_commits_info_4_debug_ldest;
        input  io_commits_info_4_debug_pdest;
        input  io_commits_info_4_debug_otherPdest_0;
        input  io_commits_info_4_debug_otherPdest_1;
        input  io_commits_info_4_debug_otherPdest_2;
        input  io_commits_info_4_debug_otherPdest_3;
        input  io_commits_info_4_debug_otherPdest_4;
        input  io_commits_info_4_debug_otherPdest_5;
        input  io_commits_info_4_debug_otherPdest_6;
        input  io_commits_info_4_debug_fuType;
        input  io_commits_info_4_dirtyFs;
        input  io_commits_info_4_dirtyVs;
        input  io_commits_info_5_walk_v;
        input  io_commits_info_5_commit_v;
        input  io_commits_info_5_commit_w;
        input  io_commits_info_5_realDestSize;
        input  io_commits_info_5_interrupt_safe;
        input  io_commits_info_5_wflags;
        input  io_commits_info_5_fflags;
        input  io_commits_info_5_vxsat;
        input  io_commits_info_5_isRVC;
        input  io_commits_info_5_isVset;
        input  io_commits_info_5_isHls;
        input  io_commits_info_5_isVls;
        input  io_commits_info_5_vls;
        input  io_commits_info_5_mmio;
        input  io_commits_info_5_commitType;
        input  io_commits_info_5_ftqIdx_flag;
        input  io_commits_info_5_ftqIdx_value;
        input  io_commits_info_5_ftqOffset;
        input  io_commits_info_5_instrSize;
        input  io_commits_info_5_fpWen;
        input  io_commits_info_5_rfWen;
        input  io_commits_info_5_needFlush;
        input  io_commits_info_5_traceBlockInPipe_itype;
        input  io_commits_info_5_traceBlockInPipe_iretire;
        input  io_commits_info_5_traceBlockInPipe_ilastsize;
        input  io_commits_info_5_debug_pc;
        input  io_commits_info_5_debug_instr;
        input  io_commits_info_5_debug_ldest;
        input  io_commits_info_5_debug_pdest;
        input  io_commits_info_5_debug_otherPdest_0;
        input  io_commits_info_5_debug_otherPdest_1;
        input  io_commits_info_5_debug_otherPdest_2;
        input  io_commits_info_5_debug_otherPdest_3;
        input  io_commits_info_5_debug_otherPdest_4;
        input  io_commits_info_5_debug_otherPdest_5;
        input  io_commits_info_5_debug_otherPdest_6;
        input  io_commits_info_5_debug_fuType;
        input  io_commits_info_5_dirtyFs;
        input  io_commits_info_5_dirtyVs;
        input  io_commits_info_6_walk_v;
        input  io_commits_info_6_commit_v;
        input  io_commits_info_6_commit_w;
        input  io_commits_info_6_realDestSize;
        input  io_commits_info_6_interrupt_safe;
        input  io_commits_info_6_wflags;
        input  io_commits_info_6_fflags;
        input  io_commits_info_6_vxsat;
        input  io_commits_info_6_isRVC;
        input  io_commits_info_6_isVset;
        input  io_commits_info_6_isHls;
        input  io_commits_info_6_isVls;
        input  io_commits_info_6_vls;
        input  io_commits_info_6_mmio;
        input  io_commits_info_6_commitType;
        input  io_commits_info_6_ftqIdx_flag;
        input  io_commits_info_6_ftqIdx_value;
        input  io_commits_info_6_ftqOffset;
        input  io_commits_info_6_instrSize;
        input  io_commits_info_6_fpWen;
        input  io_commits_info_6_rfWen;
        input  io_commits_info_6_needFlush;
        input  io_commits_info_6_traceBlockInPipe_itype;
        input  io_commits_info_6_traceBlockInPipe_iretire;
        input  io_commits_info_6_traceBlockInPipe_ilastsize;
        input  io_commits_info_6_debug_pc;
        input  io_commits_info_6_debug_instr;
        input  io_commits_info_6_debug_ldest;
        input  io_commits_info_6_debug_pdest;
        input  io_commits_info_6_debug_otherPdest_0;
        input  io_commits_info_6_debug_otherPdest_1;
        input  io_commits_info_6_debug_otherPdest_2;
        input  io_commits_info_6_debug_otherPdest_3;
        input  io_commits_info_6_debug_otherPdest_4;
        input  io_commits_info_6_debug_otherPdest_5;
        input  io_commits_info_6_debug_otherPdest_6;
        input  io_commits_info_6_debug_fuType;
        input  io_commits_info_6_dirtyFs;
        input  io_commits_info_6_dirtyVs;
        input  io_commits_info_7_walk_v;
        input  io_commits_info_7_commit_v;
        input  io_commits_info_7_commit_w;
        input  io_commits_info_7_realDestSize;
        input  io_commits_info_7_interrupt_safe;
        input  io_commits_info_7_wflags;
        input  io_commits_info_7_fflags;
        input  io_commits_info_7_vxsat;
        input  io_commits_info_7_isRVC;
        input  io_commits_info_7_isVset;
        input  io_commits_info_7_isHls;
        input  io_commits_info_7_isVls;
        input  io_commits_info_7_vls;
        input  io_commits_info_7_mmio;
        input  io_commits_info_7_commitType;
        input  io_commits_info_7_ftqIdx_flag;
        input  io_commits_info_7_ftqIdx_value;
        input  io_commits_info_7_ftqOffset;
        input  io_commits_info_7_instrSize;
        input  io_commits_info_7_fpWen;
        input  io_commits_info_7_rfWen;
        input  io_commits_info_7_needFlush;
        input  io_commits_info_7_traceBlockInPipe_itype;
        input  io_commits_info_7_traceBlockInPipe_iretire;
        input  io_commits_info_7_traceBlockInPipe_ilastsize;
        input  io_commits_info_7_debug_pc;
        input  io_commits_info_7_debug_instr;
        input  io_commits_info_7_debug_ldest;
        input  io_commits_info_7_debug_pdest;
        input  io_commits_info_7_debug_otherPdest_0;
        input  io_commits_info_7_debug_otherPdest_1;
        input  io_commits_info_7_debug_otherPdest_2;
        input  io_commits_info_7_debug_otherPdest_3;
        input  io_commits_info_7_debug_otherPdest_4;
        input  io_commits_info_7_debug_otherPdest_5;
        input  io_commits_info_7_debug_otherPdest_6;
        input  io_commits_info_7_debug_fuType;
        input  io_commits_info_7_dirtyFs;
        input  io_commits_info_7_dirtyVs;
        input  io_commits_robIdx_0_flag;
        input  io_commits_robIdx_0_value;
        input  io_commits_robIdx_1_flag;
        input  io_commits_robIdx_1_value;
        input  io_commits_robIdx_2_flag;
        input  io_commits_robIdx_2_value;
        input  io_commits_robIdx_3_flag;
        input  io_commits_robIdx_3_value;
        input  io_commits_robIdx_4_flag;
        input  io_commits_robIdx_4_value;
        input  io_commits_robIdx_5_flag;
        input  io_commits_robIdx_5_value;
        input  io_commits_robIdx_6_flag;
        input  io_commits_robIdx_6_value;
        input  io_commits_robIdx_7_flag;
        input  io_commits_robIdx_7_value;
        input  io_trace_blockCommit;
        input  io_trace_traceCommitInfo_blocks_0_valid;
        input  io_trace_traceCommitInfo_blocks_0_bits_ftqIdx_value;
        input  io_trace_traceCommitInfo_blocks_0_bits_ftqOffset;
        input  io_trace_traceCommitInfo_blocks_0_bits_tracePipe_itype;
        input  io_trace_traceCommitInfo_blocks_0_bits_tracePipe_iretire;
        input  io_trace_traceCommitInfo_blocks_0_bits_tracePipe_ilastsize;
        input  io_trace_traceCommitInfo_blocks_1_valid;
        input  io_trace_traceCommitInfo_blocks_1_bits_ftqIdx_value;
        input  io_trace_traceCommitInfo_blocks_1_bits_ftqOffset;
        input  io_trace_traceCommitInfo_blocks_1_bits_tracePipe_itype;
        input  io_trace_traceCommitInfo_blocks_1_bits_tracePipe_iretire;
        input  io_trace_traceCommitInfo_blocks_1_bits_tracePipe_ilastsize;
        input  io_trace_traceCommitInfo_blocks_2_valid;
        input  io_trace_traceCommitInfo_blocks_2_bits_ftqIdx_value;
        input  io_trace_traceCommitInfo_blocks_2_bits_ftqOffset;
        input  io_trace_traceCommitInfo_blocks_2_bits_tracePipe_itype;
        input  io_trace_traceCommitInfo_blocks_2_bits_tracePipe_iretire;
        input  io_trace_traceCommitInfo_blocks_2_bits_tracePipe_ilastsize;
        input  io_trace_traceCommitInfo_blocks_3_valid;
        input  io_trace_traceCommitInfo_blocks_3_bits_ftqIdx_value;
        input  io_trace_traceCommitInfo_blocks_3_bits_ftqOffset;
        input  io_trace_traceCommitInfo_blocks_3_bits_tracePipe_itype;
        input  io_trace_traceCommitInfo_blocks_3_bits_tracePipe_iretire;
        input  io_trace_traceCommitInfo_blocks_3_bits_tracePipe_ilastsize;
        input  io_trace_traceCommitInfo_blocks_4_valid;
        input  io_trace_traceCommitInfo_blocks_4_bits_ftqIdx_value;
        input  io_trace_traceCommitInfo_blocks_4_bits_ftqOffset;
        input  io_trace_traceCommitInfo_blocks_4_bits_tracePipe_itype;
        input  io_trace_traceCommitInfo_blocks_4_bits_tracePipe_iretire;
        input  io_trace_traceCommitInfo_blocks_4_bits_tracePipe_ilastsize;
        input  io_trace_traceCommitInfo_blocks_5_valid;
        input  io_trace_traceCommitInfo_blocks_5_bits_ftqIdx_value;
        input  io_trace_traceCommitInfo_blocks_5_bits_ftqOffset;
        input  io_trace_traceCommitInfo_blocks_5_bits_tracePipe_itype;
        input  io_trace_traceCommitInfo_blocks_5_bits_tracePipe_iretire;
        input  io_trace_traceCommitInfo_blocks_5_bits_tracePipe_ilastsize;
        input  io_trace_traceCommitInfo_blocks_6_valid;
        input  io_trace_traceCommitInfo_blocks_6_bits_ftqIdx_value;
        input  io_trace_traceCommitInfo_blocks_6_bits_ftqOffset;
        input  io_trace_traceCommitInfo_blocks_6_bits_tracePipe_itype;
        input  io_trace_traceCommitInfo_blocks_6_bits_tracePipe_iretire;
        input  io_trace_traceCommitInfo_blocks_6_bits_tracePipe_ilastsize;
        input  io_trace_traceCommitInfo_blocks_7_valid;
        input  io_trace_traceCommitInfo_blocks_7_bits_ftqIdx_value;
        input  io_trace_traceCommitInfo_blocks_7_bits_ftqOffset;
        input  io_trace_traceCommitInfo_blocks_7_bits_tracePipe_itype;
        input  io_trace_traceCommitInfo_blocks_7_bits_tracePipe_iretire;
        input  io_trace_traceCommitInfo_blocks_7_bits_tracePipe_ilastsize;
        input  io_rabCommits_isCommit;
        input  io_rabCommits_commitValid_0;
        input  io_rabCommits_commitValid_1;
        input  io_rabCommits_commitValid_2;
        input  io_rabCommits_commitValid_3;
        input  io_rabCommits_commitValid_4;
        input  io_rabCommits_commitValid_5;
        input  io_rabCommits_isWalk;
        input  io_rabCommits_walkValid_0;
        input  io_rabCommits_walkValid_1;
        input  io_rabCommits_walkValid_2;
        input  io_rabCommits_walkValid_3;
        input  io_rabCommits_walkValid_4;
        input  io_rabCommits_walkValid_5;
        input  io_rabCommits_info_0_ldest;
        input  io_rabCommits_info_0_pdest;
        input  io_rabCommits_info_0_rfWen;
        input  io_rabCommits_info_0_fpWen;
        input  io_rabCommits_info_0_vecWen;
        input  io_rabCommits_info_0_v0Wen;
        input  io_rabCommits_info_0_vlWen;
        input  io_rabCommits_info_0_isMove;
        input  io_rabCommits_info_1_ldest;
        input  io_rabCommits_info_1_pdest;
        input  io_rabCommits_info_1_rfWen;
        input  io_rabCommits_info_1_fpWen;
        input  io_rabCommits_info_1_vecWen;
        input  io_rabCommits_info_1_v0Wen;
        input  io_rabCommits_info_1_vlWen;
        input  io_rabCommits_info_1_isMove;
        input  io_rabCommits_info_2_ldest;
        input  io_rabCommits_info_2_pdest;
        input  io_rabCommits_info_2_rfWen;
        input  io_rabCommits_info_2_fpWen;
        input  io_rabCommits_info_2_vecWen;
        input  io_rabCommits_info_2_v0Wen;
        input  io_rabCommits_info_2_vlWen;
        input  io_rabCommits_info_2_isMove;
        input  io_rabCommits_info_3_ldest;
        input  io_rabCommits_info_3_pdest;
        input  io_rabCommits_info_3_rfWen;
        input  io_rabCommits_info_3_fpWen;
        input  io_rabCommits_info_3_vecWen;
        input  io_rabCommits_info_3_v0Wen;
        input  io_rabCommits_info_3_vlWen;
        input  io_rabCommits_info_3_isMove;
        input  io_rabCommits_info_4_ldest;
        input  io_rabCommits_info_4_pdest;
        input  io_rabCommits_info_4_rfWen;
        input  io_rabCommits_info_4_fpWen;
        input  io_rabCommits_info_4_vecWen;
        input  io_rabCommits_info_4_v0Wen;
        input  io_rabCommits_info_4_vlWen;
        input  io_rabCommits_info_4_isMove;
        input  io_rabCommits_info_5_ldest;
        input  io_rabCommits_info_5_pdest;
        input  io_rabCommits_info_5_rfWen;
        input  io_rabCommits_info_5_fpWen;
        input  io_rabCommits_info_5_vecWen;
        input  io_rabCommits_info_5_v0Wen;
        input  io_rabCommits_info_5_vlWen;
        input  io_rabCommits_info_5_isMove;
        input  io_diffCommits_commitValid_0;
        input  io_diffCommits_commitValid_1;
        input  io_diffCommits_commitValid_2;
        input  io_diffCommits_commitValid_3;
        input  io_diffCommits_commitValid_4;
        input  io_diffCommits_commitValid_5;
        input  io_diffCommits_commitValid_6;
        input  io_diffCommits_commitValid_7;
        input  io_diffCommits_commitValid_8;
        input  io_diffCommits_commitValid_9;
        input  io_diffCommits_commitValid_10;
        input  io_diffCommits_commitValid_11;
        input  io_diffCommits_commitValid_12;
        input  io_diffCommits_commitValid_13;
        input  io_diffCommits_commitValid_14;
        input  io_diffCommits_commitValid_15;
        input  io_diffCommits_commitValid_16;
        input  io_diffCommits_commitValid_17;
        input  io_diffCommits_commitValid_18;
        input  io_diffCommits_commitValid_19;
        input  io_diffCommits_commitValid_20;
        input  io_diffCommits_commitValid_21;
        input  io_diffCommits_commitValid_22;
        input  io_diffCommits_commitValid_23;
        input  io_diffCommits_commitValid_24;
        input  io_diffCommits_commitValid_25;
        input  io_diffCommits_commitValid_26;
        input  io_diffCommits_commitValid_27;
        input  io_diffCommits_commitValid_28;
        input  io_diffCommits_commitValid_29;
        input  io_diffCommits_commitValid_30;
        input  io_diffCommits_commitValid_31;
        input  io_diffCommits_commitValid_32;
        input  io_diffCommits_commitValid_33;
        input  io_diffCommits_commitValid_34;
        input  io_diffCommits_commitValid_35;
        input  io_diffCommits_commitValid_36;
        input  io_diffCommits_commitValid_37;
        input  io_diffCommits_commitValid_38;
        input  io_diffCommits_commitValid_39;
        input  io_diffCommits_commitValid_40;
        input  io_diffCommits_commitValid_41;
        input  io_diffCommits_commitValid_42;
        input  io_diffCommits_commitValid_43;
        input  io_diffCommits_commitValid_44;
        input  io_diffCommits_commitValid_45;
        input  io_diffCommits_commitValid_46;
        input  io_diffCommits_commitValid_47;
        input  io_diffCommits_commitValid_48;
        input  io_diffCommits_commitValid_49;
        input  io_diffCommits_commitValid_50;
        input  io_diffCommits_commitValid_51;
        input  io_diffCommits_commitValid_52;
        input  io_diffCommits_commitValid_53;
        input  io_diffCommits_commitValid_54;
        input  io_diffCommits_commitValid_55;
        input  io_diffCommits_commitValid_56;
        input  io_diffCommits_commitValid_57;
        input  io_diffCommits_commitValid_58;
        input  io_diffCommits_commitValid_59;
        input  io_diffCommits_commitValid_60;
        input  io_diffCommits_commitValid_61;
        input  io_diffCommits_commitValid_62;
        input  io_diffCommits_commitValid_63;
        input  io_diffCommits_commitValid_64;
        input  io_diffCommits_commitValid_65;
        input  io_diffCommits_commitValid_66;
        input  io_diffCommits_commitValid_67;
        input  io_diffCommits_commitValid_68;
        input  io_diffCommits_commitValid_69;
        input  io_diffCommits_commitValid_70;
        input  io_diffCommits_commitValid_71;
        input  io_diffCommits_commitValid_72;
        input  io_diffCommits_commitValid_73;
        input  io_diffCommits_commitValid_74;
        input  io_diffCommits_commitValid_75;
        input  io_diffCommits_commitValid_76;
        input  io_diffCommits_commitValid_77;
        input  io_diffCommits_commitValid_78;
        input  io_diffCommits_commitValid_79;
        input  io_diffCommits_commitValid_80;
        input  io_diffCommits_commitValid_81;
        input  io_diffCommits_commitValid_82;
        input  io_diffCommits_commitValid_83;
        input  io_diffCommits_commitValid_84;
        input  io_diffCommits_commitValid_85;
        input  io_diffCommits_commitValid_86;
        input  io_diffCommits_commitValid_87;
        input  io_diffCommits_commitValid_88;
        input  io_diffCommits_commitValid_89;
        input  io_diffCommits_commitValid_90;
        input  io_diffCommits_commitValid_91;
        input  io_diffCommits_commitValid_92;
        input  io_diffCommits_commitValid_93;
        input  io_diffCommits_commitValid_94;
        input  io_diffCommits_commitValid_95;
        input  io_diffCommits_commitValid_96;
        input  io_diffCommits_commitValid_97;
        input  io_diffCommits_commitValid_98;
        input  io_diffCommits_commitValid_99;
        input  io_diffCommits_commitValid_100;
        input  io_diffCommits_commitValid_101;
        input  io_diffCommits_commitValid_102;
        input  io_diffCommits_commitValid_103;
        input  io_diffCommits_commitValid_104;
        input  io_diffCommits_commitValid_105;
        input  io_diffCommits_commitValid_106;
        input  io_diffCommits_commitValid_107;
        input  io_diffCommits_commitValid_108;
        input  io_diffCommits_commitValid_109;
        input  io_diffCommits_commitValid_110;
        input  io_diffCommits_commitValid_111;
        input  io_diffCommits_commitValid_112;
        input  io_diffCommits_commitValid_113;
        input  io_diffCommits_commitValid_114;
        input  io_diffCommits_commitValid_115;
        input  io_diffCommits_commitValid_116;
        input  io_diffCommits_commitValid_117;
        input  io_diffCommits_commitValid_118;
        input  io_diffCommits_commitValid_119;
        input  io_diffCommits_commitValid_120;
        input  io_diffCommits_commitValid_121;
        input  io_diffCommits_commitValid_122;
        input  io_diffCommits_commitValid_123;
        input  io_diffCommits_commitValid_124;
        input  io_diffCommits_commitValid_125;
        input  io_diffCommits_commitValid_126;
        input  io_diffCommits_commitValid_127;
        input  io_diffCommits_commitValid_128;
        input  io_diffCommits_commitValid_129;
        input  io_diffCommits_commitValid_130;
        input  io_diffCommits_commitValid_131;
        input  io_diffCommits_commitValid_132;
        input  io_diffCommits_commitValid_133;
        input  io_diffCommits_commitValid_134;
        input  io_diffCommits_commitValid_135;
        input  io_diffCommits_commitValid_136;
        input  io_diffCommits_commitValid_137;
        input  io_diffCommits_commitValid_138;
        input  io_diffCommits_commitValid_139;
        input  io_diffCommits_commitValid_140;
        input  io_diffCommits_commitValid_141;
        input  io_diffCommits_commitValid_142;
        input  io_diffCommits_commitValid_143;
        input  io_diffCommits_commitValid_144;
        input  io_diffCommits_commitValid_145;
        input  io_diffCommits_commitValid_146;
        input  io_diffCommits_commitValid_147;
        input  io_diffCommits_commitValid_148;
        input  io_diffCommits_commitValid_149;
        input  io_diffCommits_commitValid_150;
        input  io_diffCommits_commitValid_151;
        input  io_diffCommits_commitValid_152;
        input  io_diffCommits_commitValid_153;
        input  io_diffCommits_commitValid_154;
        input  io_diffCommits_commitValid_155;
        input  io_diffCommits_commitValid_156;
        input  io_diffCommits_commitValid_157;
        input  io_diffCommits_commitValid_158;
        input  io_diffCommits_commitValid_159;
        input  io_diffCommits_commitValid_160;
        input  io_diffCommits_commitValid_161;
        input  io_diffCommits_commitValid_162;
        input  io_diffCommits_commitValid_163;
        input  io_diffCommits_commitValid_164;
        input  io_diffCommits_commitValid_165;
        input  io_diffCommits_commitValid_166;
        input  io_diffCommits_commitValid_167;
        input  io_diffCommits_commitValid_168;
        input  io_diffCommits_commitValid_169;
        input  io_diffCommits_commitValid_170;
        input  io_diffCommits_commitValid_171;
        input  io_diffCommits_commitValid_172;
        input  io_diffCommits_commitValid_173;
        input  io_diffCommits_commitValid_174;
        input  io_diffCommits_commitValid_175;
        input  io_diffCommits_commitValid_176;
        input  io_diffCommits_commitValid_177;
        input  io_diffCommits_commitValid_178;
        input  io_diffCommits_commitValid_179;
        input  io_diffCommits_commitValid_180;
        input  io_diffCommits_commitValid_181;
        input  io_diffCommits_commitValid_182;
        input  io_diffCommits_commitValid_183;
        input  io_diffCommits_commitValid_184;
        input  io_diffCommits_commitValid_185;
        input  io_diffCommits_commitValid_186;
        input  io_diffCommits_commitValid_187;
        input  io_diffCommits_commitValid_188;
        input  io_diffCommits_commitValid_189;
        input  io_diffCommits_commitValid_190;
        input  io_diffCommits_commitValid_191;
        input  io_diffCommits_commitValid_192;
        input  io_diffCommits_commitValid_193;
        input  io_diffCommits_commitValid_194;
        input  io_diffCommits_commitValid_195;
        input  io_diffCommits_commitValid_196;
        input  io_diffCommits_commitValid_197;
        input  io_diffCommits_commitValid_198;
        input  io_diffCommits_commitValid_199;
        input  io_diffCommits_commitValid_200;
        input  io_diffCommits_commitValid_201;
        input  io_diffCommits_commitValid_202;
        input  io_diffCommits_commitValid_203;
        input  io_diffCommits_commitValid_204;
        input  io_diffCommits_commitValid_205;
        input  io_diffCommits_commitValid_206;
        input  io_diffCommits_commitValid_207;
        input  io_diffCommits_commitValid_208;
        input  io_diffCommits_commitValid_209;
        input  io_diffCommits_commitValid_210;
        input  io_diffCommits_commitValid_211;
        input  io_diffCommits_commitValid_212;
        input  io_diffCommits_commitValid_213;
        input  io_diffCommits_commitValid_214;
        input  io_diffCommits_commitValid_215;
        input  io_diffCommits_commitValid_216;
        input  io_diffCommits_commitValid_217;
        input  io_diffCommits_commitValid_218;
        input  io_diffCommits_commitValid_219;
        input  io_diffCommits_commitValid_220;
        input  io_diffCommits_commitValid_221;
        input  io_diffCommits_commitValid_222;
        input  io_diffCommits_commitValid_223;
        input  io_diffCommits_commitValid_224;
        input  io_diffCommits_commitValid_225;
        input  io_diffCommits_commitValid_226;
        input  io_diffCommits_commitValid_227;
        input  io_diffCommits_commitValid_228;
        input  io_diffCommits_commitValid_229;
        input  io_diffCommits_commitValid_230;
        input  io_diffCommits_commitValid_231;
        input  io_diffCommits_commitValid_232;
        input  io_diffCommits_commitValid_233;
        input  io_diffCommits_commitValid_234;
        input  io_diffCommits_commitValid_235;
        input  io_diffCommits_commitValid_236;
        input  io_diffCommits_commitValid_237;
        input  io_diffCommits_commitValid_238;
        input  io_diffCommits_commitValid_239;
        input  io_diffCommits_commitValid_240;
        input  io_diffCommits_commitValid_241;
        input  io_diffCommits_commitValid_242;
        input  io_diffCommits_commitValid_243;
        input  io_diffCommits_commitValid_244;
        input  io_diffCommits_commitValid_245;
        input  io_diffCommits_commitValid_246;
        input  io_diffCommits_commitValid_247;
        input  io_diffCommits_commitValid_248;
        input  io_diffCommits_commitValid_249;
        input  io_diffCommits_commitValid_250;
        input  io_diffCommits_commitValid_251;
        input  io_diffCommits_commitValid_252;
        input  io_diffCommits_commitValid_253;
        input  io_diffCommits_commitValid_254;
        input  io_diffCommits_info_0_ldest;
        input  io_diffCommits_info_0_pdest;
        input  io_diffCommits_info_0_rfWen;
        input  io_diffCommits_info_0_fpWen;
        input  io_diffCommits_info_0_vecWen;
        input  io_diffCommits_info_0_v0Wen;
        input  io_diffCommits_info_0_vlWen;
        input  io_diffCommits_info_1_ldest;
        input  io_diffCommits_info_1_pdest;
        input  io_diffCommits_info_1_rfWen;
        input  io_diffCommits_info_1_fpWen;
        input  io_diffCommits_info_1_vecWen;
        input  io_diffCommits_info_1_v0Wen;
        input  io_diffCommits_info_1_vlWen;
        input  io_diffCommits_info_2_ldest;
        input  io_diffCommits_info_2_pdest;
        input  io_diffCommits_info_2_rfWen;
        input  io_diffCommits_info_2_fpWen;
        input  io_diffCommits_info_2_vecWen;
        input  io_diffCommits_info_2_v0Wen;
        input  io_diffCommits_info_2_vlWen;
        input  io_diffCommits_info_3_ldest;
        input  io_diffCommits_info_3_pdest;
        input  io_diffCommits_info_3_rfWen;
        input  io_diffCommits_info_3_fpWen;
        input  io_diffCommits_info_3_vecWen;
        input  io_diffCommits_info_3_v0Wen;
        input  io_diffCommits_info_3_vlWen;
        input  io_diffCommits_info_4_ldest;
        input  io_diffCommits_info_4_pdest;
        input  io_diffCommits_info_4_rfWen;
        input  io_diffCommits_info_4_fpWen;
        input  io_diffCommits_info_4_vecWen;
        input  io_diffCommits_info_4_v0Wen;
        input  io_diffCommits_info_4_vlWen;
        input  io_diffCommits_info_5_ldest;
        input  io_diffCommits_info_5_pdest;
        input  io_diffCommits_info_5_rfWen;
        input  io_diffCommits_info_5_fpWen;
        input  io_diffCommits_info_5_vecWen;
        input  io_diffCommits_info_5_v0Wen;
        input  io_diffCommits_info_5_vlWen;
        input  io_diffCommits_info_6_ldest;
        input  io_diffCommits_info_6_pdest;
        input  io_diffCommits_info_6_rfWen;
        input  io_diffCommits_info_6_fpWen;
        input  io_diffCommits_info_6_vecWen;
        input  io_diffCommits_info_6_v0Wen;
        input  io_diffCommits_info_6_vlWen;
        input  io_diffCommits_info_7_ldest;
        input  io_diffCommits_info_7_pdest;
        input  io_diffCommits_info_7_rfWen;
        input  io_diffCommits_info_7_fpWen;
        input  io_diffCommits_info_7_vecWen;
        input  io_diffCommits_info_7_v0Wen;
        input  io_diffCommits_info_7_vlWen;
        input  io_diffCommits_info_8_ldest;
        input  io_diffCommits_info_8_pdest;
        input  io_diffCommits_info_8_rfWen;
        input  io_diffCommits_info_8_fpWen;
        input  io_diffCommits_info_8_vecWen;
        input  io_diffCommits_info_8_v0Wen;
        input  io_diffCommits_info_8_vlWen;
        input  io_diffCommits_info_9_ldest;
        input  io_diffCommits_info_9_pdest;
        input  io_diffCommits_info_9_rfWen;
        input  io_diffCommits_info_9_fpWen;
        input  io_diffCommits_info_9_vecWen;
        input  io_diffCommits_info_9_v0Wen;
        input  io_diffCommits_info_9_vlWen;
        input  io_diffCommits_info_10_ldest;
        input  io_diffCommits_info_10_pdest;
        input  io_diffCommits_info_10_rfWen;
        input  io_diffCommits_info_10_fpWen;
        input  io_diffCommits_info_10_vecWen;
        input  io_diffCommits_info_10_v0Wen;
        input  io_diffCommits_info_10_vlWen;
        input  io_diffCommits_info_11_ldest;
        input  io_diffCommits_info_11_pdest;
        input  io_diffCommits_info_11_rfWen;
        input  io_diffCommits_info_11_fpWen;
        input  io_diffCommits_info_11_vecWen;
        input  io_diffCommits_info_11_v0Wen;
        input  io_diffCommits_info_11_vlWen;
        input  io_diffCommits_info_12_ldest;
        input  io_diffCommits_info_12_pdest;
        input  io_diffCommits_info_12_rfWen;
        input  io_diffCommits_info_12_fpWen;
        input  io_diffCommits_info_12_vecWen;
        input  io_diffCommits_info_12_v0Wen;
        input  io_diffCommits_info_12_vlWen;
        input  io_diffCommits_info_13_ldest;
        input  io_diffCommits_info_13_pdest;
        input  io_diffCommits_info_13_rfWen;
        input  io_diffCommits_info_13_fpWen;
        input  io_diffCommits_info_13_vecWen;
        input  io_diffCommits_info_13_v0Wen;
        input  io_diffCommits_info_13_vlWen;
        input  io_diffCommits_info_14_ldest;
        input  io_diffCommits_info_14_pdest;
        input  io_diffCommits_info_14_rfWen;
        input  io_diffCommits_info_14_fpWen;
        input  io_diffCommits_info_14_vecWen;
        input  io_diffCommits_info_14_v0Wen;
        input  io_diffCommits_info_14_vlWen;
        input  io_diffCommits_info_15_ldest;
        input  io_diffCommits_info_15_pdest;
        input  io_diffCommits_info_15_rfWen;
        input  io_diffCommits_info_15_fpWen;
        input  io_diffCommits_info_15_vecWen;
        input  io_diffCommits_info_15_v0Wen;
        input  io_diffCommits_info_15_vlWen;
        input  io_diffCommits_info_16_ldest;
        input  io_diffCommits_info_16_pdest;
        input  io_diffCommits_info_16_rfWen;
        input  io_diffCommits_info_16_fpWen;
        input  io_diffCommits_info_16_vecWen;
        input  io_diffCommits_info_16_v0Wen;
        input  io_diffCommits_info_16_vlWen;
        input  io_diffCommits_info_17_ldest;
        input  io_diffCommits_info_17_pdest;
        input  io_diffCommits_info_17_rfWen;
        input  io_diffCommits_info_17_fpWen;
        input  io_diffCommits_info_17_vecWen;
        input  io_diffCommits_info_17_v0Wen;
        input  io_diffCommits_info_17_vlWen;
        input  io_diffCommits_info_18_ldest;
        input  io_diffCommits_info_18_pdest;
        input  io_diffCommits_info_18_rfWen;
        input  io_diffCommits_info_18_fpWen;
        input  io_diffCommits_info_18_vecWen;
        input  io_diffCommits_info_18_v0Wen;
        input  io_diffCommits_info_18_vlWen;
        input  io_diffCommits_info_19_ldest;
        input  io_diffCommits_info_19_pdest;
        input  io_diffCommits_info_19_rfWen;
        input  io_diffCommits_info_19_fpWen;
        input  io_diffCommits_info_19_vecWen;
        input  io_diffCommits_info_19_v0Wen;
        input  io_diffCommits_info_19_vlWen;
        input  io_diffCommits_info_20_ldest;
        input  io_diffCommits_info_20_pdest;
        input  io_diffCommits_info_20_rfWen;
        input  io_diffCommits_info_20_fpWen;
        input  io_diffCommits_info_20_vecWen;
        input  io_diffCommits_info_20_v0Wen;
        input  io_diffCommits_info_20_vlWen;
        input  io_diffCommits_info_21_ldest;
        input  io_diffCommits_info_21_pdest;
        input  io_diffCommits_info_21_rfWen;
        input  io_diffCommits_info_21_fpWen;
        input  io_diffCommits_info_21_vecWen;
        input  io_diffCommits_info_21_v0Wen;
        input  io_diffCommits_info_21_vlWen;
        input  io_diffCommits_info_22_ldest;
        input  io_diffCommits_info_22_pdest;
        input  io_diffCommits_info_22_rfWen;
        input  io_diffCommits_info_22_fpWen;
        input  io_diffCommits_info_22_vecWen;
        input  io_diffCommits_info_22_v0Wen;
        input  io_diffCommits_info_22_vlWen;
        input  io_diffCommits_info_23_ldest;
        input  io_diffCommits_info_23_pdest;
        input  io_diffCommits_info_23_rfWen;
        input  io_diffCommits_info_23_fpWen;
        input  io_diffCommits_info_23_vecWen;
        input  io_diffCommits_info_23_v0Wen;
        input  io_diffCommits_info_23_vlWen;
        input  io_diffCommits_info_24_ldest;
        input  io_diffCommits_info_24_pdest;
        input  io_diffCommits_info_24_rfWen;
        input  io_diffCommits_info_24_fpWen;
        input  io_diffCommits_info_24_vecWen;
        input  io_diffCommits_info_24_v0Wen;
        input  io_diffCommits_info_24_vlWen;
        input  io_diffCommits_info_25_ldest;
        input  io_diffCommits_info_25_pdest;
        input  io_diffCommits_info_25_rfWen;
        input  io_diffCommits_info_25_fpWen;
        input  io_diffCommits_info_25_vecWen;
        input  io_diffCommits_info_25_v0Wen;
        input  io_diffCommits_info_25_vlWen;
        input  io_diffCommits_info_26_ldest;
        input  io_diffCommits_info_26_pdest;
        input  io_diffCommits_info_26_rfWen;
        input  io_diffCommits_info_26_fpWen;
        input  io_diffCommits_info_26_vecWen;
        input  io_diffCommits_info_26_v0Wen;
        input  io_diffCommits_info_26_vlWen;
        input  io_diffCommits_info_27_ldest;
        input  io_diffCommits_info_27_pdest;
        input  io_diffCommits_info_27_rfWen;
        input  io_diffCommits_info_27_fpWen;
        input  io_diffCommits_info_27_vecWen;
        input  io_diffCommits_info_27_v0Wen;
        input  io_diffCommits_info_27_vlWen;
        input  io_diffCommits_info_28_ldest;
        input  io_diffCommits_info_28_pdest;
        input  io_diffCommits_info_28_rfWen;
        input  io_diffCommits_info_28_fpWen;
        input  io_diffCommits_info_28_vecWen;
        input  io_diffCommits_info_28_v0Wen;
        input  io_diffCommits_info_28_vlWen;
        input  io_diffCommits_info_29_ldest;
        input  io_diffCommits_info_29_pdest;
        input  io_diffCommits_info_29_rfWen;
        input  io_diffCommits_info_29_fpWen;
        input  io_diffCommits_info_29_vecWen;
        input  io_diffCommits_info_29_v0Wen;
        input  io_diffCommits_info_29_vlWen;
        input  io_diffCommits_info_30_ldest;
        input  io_diffCommits_info_30_pdest;
        input  io_diffCommits_info_30_rfWen;
        input  io_diffCommits_info_30_fpWen;
        input  io_diffCommits_info_30_vecWen;
        input  io_diffCommits_info_30_v0Wen;
        input  io_diffCommits_info_30_vlWen;
        input  io_diffCommits_info_31_ldest;
        input  io_diffCommits_info_31_pdest;
        input  io_diffCommits_info_31_rfWen;
        input  io_diffCommits_info_31_fpWen;
        input  io_diffCommits_info_31_vecWen;
        input  io_diffCommits_info_31_v0Wen;
        input  io_diffCommits_info_31_vlWen;
        input  io_diffCommits_info_32_ldest;
        input  io_diffCommits_info_32_pdest;
        input  io_diffCommits_info_32_rfWen;
        input  io_diffCommits_info_32_fpWen;
        input  io_diffCommits_info_32_vecWen;
        input  io_diffCommits_info_32_v0Wen;
        input  io_diffCommits_info_32_vlWen;
        input  io_diffCommits_info_33_ldest;
        input  io_diffCommits_info_33_pdest;
        input  io_diffCommits_info_33_rfWen;
        input  io_diffCommits_info_33_fpWen;
        input  io_diffCommits_info_33_vecWen;
        input  io_diffCommits_info_33_v0Wen;
        input  io_diffCommits_info_33_vlWen;
        input  io_diffCommits_info_34_ldest;
        input  io_diffCommits_info_34_pdest;
        input  io_diffCommits_info_34_rfWen;
        input  io_diffCommits_info_34_fpWen;
        input  io_diffCommits_info_34_vecWen;
        input  io_diffCommits_info_34_v0Wen;
        input  io_diffCommits_info_34_vlWen;
        input  io_diffCommits_info_35_ldest;
        input  io_diffCommits_info_35_pdest;
        input  io_diffCommits_info_35_rfWen;
        input  io_diffCommits_info_35_fpWen;
        input  io_diffCommits_info_35_vecWen;
        input  io_diffCommits_info_35_v0Wen;
        input  io_diffCommits_info_35_vlWen;
        input  io_diffCommits_info_36_ldest;
        input  io_diffCommits_info_36_pdest;
        input  io_diffCommits_info_36_rfWen;
        input  io_diffCommits_info_36_fpWen;
        input  io_diffCommits_info_36_vecWen;
        input  io_diffCommits_info_36_v0Wen;
        input  io_diffCommits_info_36_vlWen;
        input  io_diffCommits_info_37_ldest;
        input  io_diffCommits_info_37_pdest;
        input  io_diffCommits_info_37_rfWen;
        input  io_diffCommits_info_37_fpWen;
        input  io_diffCommits_info_37_vecWen;
        input  io_diffCommits_info_37_v0Wen;
        input  io_diffCommits_info_37_vlWen;
        input  io_diffCommits_info_38_ldest;
        input  io_diffCommits_info_38_pdest;
        input  io_diffCommits_info_38_rfWen;
        input  io_diffCommits_info_38_fpWen;
        input  io_diffCommits_info_38_vecWen;
        input  io_diffCommits_info_38_v0Wen;
        input  io_diffCommits_info_38_vlWen;
        input  io_diffCommits_info_39_ldest;
        input  io_diffCommits_info_39_pdest;
        input  io_diffCommits_info_39_rfWen;
        input  io_diffCommits_info_39_fpWen;
        input  io_diffCommits_info_39_vecWen;
        input  io_diffCommits_info_39_v0Wen;
        input  io_diffCommits_info_39_vlWen;
        input  io_diffCommits_info_40_ldest;
        input  io_diffCommits_info_40_pdest;
        input  io_diffCommits_info_40_rfWen;
        input  io_diffCommits_info_40_fpWen;
        input  io_diffCommits_info_40_vecWen;
        input  io_diffCommits_info_40_v0Wen;
        input  io_diffCommits_info_40_vlWen;
        input  io_diffCommits_info_41_ldest;
        input  io_diffCommits_info_41_pdest;
        input  io_diffCommits_info_41_rfWen;
        input  io_diffCommits_info_41_fpWen;
        input  io_diffCommits_info_41_vecWen;
        input  io_diffCommits_info_41_v0Wen;
        input  io_diffCommits_info_41_vlWen;
        input  io_diffCommits_info_42_ldest;
        input  io_diffCommits_info_42_pdest;
        input  io_diffCommits_info_42_rfWen;
        input  io_diffCommits_info_42_fpWen;
        input  io_diffCommits_info_42_vecWen;
        input  io_diffCommits_info_42_v0Wen;
        input  io_diffCommits_info_42_vlWen;
        input  io_diffCommits_info_43_ldest;
        input  io_diffCommits_info_43_pdest;
        input  io_diffCommits_info_43_rfWen;
        input  io_diffCommits_info_43_fpWen;
        input  io_diffCommits_info_43_vecWen;
        input  io_diffCommits_info_43_v0Wen;
        input  io_diffCommits_info_43_vlWen;
        input  io_diffCommits_info_44_ldest;
        input  io_diffCommits_info_44_pdest;
        input  io_diffCommits_info_44_rfWen;
        input  io_diffCommits_info_44_fpWen;
        input  io_diffCommits_info_44_vecWen;
        input  io_diffCommits_info_44_v0Wen;
        input  io_diffCommits_info_44_vlWen;
        input  io_diffCommits_info_45_ldest;
        input  io_diffCommits_info_45_pdest;
        input  io_diffCommits_info_45_rfWen;
        input  io_diffCommits_info_45_fpWen;
        input  io_diffCommits_info_45_vecWen;
        input  io_diffCommits_info_45_v0Wen;
        input  io_diffCommits_info_45_vlWen;
        input  io_diffCommits_info_46_ldest;
        input  io_diffCommits_info_46_pdest;
        input  io_diffCommits_info_46_rfWen;
        input  io_diffCommits_info_46_fpWen;
        input  io_diffCommits_info_46_vecWen;
        input  io_diffCommits_info_46_v0Wen;
        input  io_diffCommits_info_46_vlWen;
        input  io_diffCommits_info_47_ldest;
        input  io_diffCommits_info_47_pdest;
        input  io_diffCommits_info_47_rfWen;
        input  io_diffCommits_info_47_fpWen;
        input  io_diffCommits_info_47_vecWen;
        input  io_diffCommits_info_47_v0Wen;
        input  io_diffCommits_info_47_vlWen;
        input  io_diffCommits_info_48_ldest;
        input  io_diffCommits_info_48_pdest;
        input  io_diffCommits_info_48_rfWen;
        input  io_diffCommits_info_48_fpWen;
        input  io_diffCommits_info_48_vecWen;
        input  io_diffCommits_info_48_v0Wen;
        input  io_diffCommits_info_48_vlWen;
        input  io_diffCommits_info_49_ldest;
        input  io_diffCommits_info_49_pdest;
        input  io_diffCommits_info_49_rfWen;
        input  io_diffCommits_info_49_fpWen;
        input  io_diffCommits_info_49_vecWen;
        input  io_diffCommits_info_49_v0Wen;
        input  io_diffCommits_info_49_vlWen;
        input  io_diffCommits_info_50_ldest;
        input  io_diffCommits_info_50_pdest;
        input  io_diffCommits_info_50_rfWen;
        input  io_diffCommits_info_50_fpWen;
        input  io_diffCommits_info_50_vecWen;
        input  io_diffCommits_info_50_v0Wen;
        input  io_diffCommits_info_50_vlWen;
        input  io_diffCommits_info_51_ldest;
        input  io_diffCommits_info_51_pdest;
        input  io_diffCommits_info_51_rfWen;
        input  io_diffCommits_info_51_fpWen;
        input  io_diffCommits_info_51_vecWen;
        input  io_diffCommits_info_51_v0Wen;
        input  io_diffCommits_info_51_vlWen;
        input  io_diffCommits_info_52_ldest;
        input  io_diffCommits_info_52_pdest;
        input  io_diffCommits_info_52_rfWen;
        input  io_diffCommits_info_52_fpWen;
        input  io_diffCommits_info_52_vecWen;
        input  io_diffCommits_info_52_v0Wen;
        input  io_diffCommits_info_52_vlWen;
        input  io_diffCommits_info_53_ldest;
        input  io_diffCommits_info_53_pdest;
        input  io_diffCommits_info_53_rfWen;
        input  io_diffCommits_info_53_fpWen;
        input  io_diffCommits_info_53_vecWen;
        input  io_diffCommits_info_53_v0Wen;
        input  io_diffCommits_info_53_vlWen;
        input  io_diffCommits_info_54_ldest;
        input  io_diffCommits_info_54_pdest;
        input  io_diffCommits_info_54_rfWen;
        input  io_diffCommits_info_54_fpWen;
        input  io_diffCommits_info_54_vecWen;
        input  io_diffCommits_info_54_v0Wen;
        input  io_diffCommits_info_54_vlWen;
        input  io_diffCommits_info_55_ldest;
        input  io_diffCommits_info_55_pdest;
        input  io_diffCommits_info_55_rfWen;
        input  io_diffCommits_info_55_fpWen;
        input  io_diffCommits_info_55_vecWen;
        input  io_diffCommits_info_55_v0Wen;
        input  io_diffCommits_info_55_vlWen;
        input  io_diffCommits_info_56_ldest;
        input  io_diffCommits_info_56_pdest;
        input  io_diffCommits_info_56_rfWen;
        input  io_diffCommits_info_56_fpWen;
        input  io_diffCommits_info_56_vecWen;
        input  io_diffCommits_info_56_v0Wen;
        input  io_diffCommits_info_56_vlWen;
        input  io_diffCommits_info_57_ldest;
        input  io_diffCommits_info_57_pdest;
        input  io_diffCommits_info_57_rfWen;
        input  io_diffCommits_info_57_fpWen;
        input  io_diffCommits_info_57_vecWen;
        input  io_diffCommits_info_57_v0Wen;
        input  io_diffCommits_info_57_vlWen;
        input  io_diffCommits_info_58_ldest;
        input  io_diffCommits_info_58_pdest;
        input  io_diffCommits_info_58_rfWen;
        input  io_diffCommits_info_58_fpWen;
        input  io_diffCommits_info_58_vecWen;
        input  io_diffCommits_info_58_v0Wen;
        input  io_diffCommits_info_58_vlWen;
        input  io_diffCommits_info_59_ldest;
        input  io_diffCommits_info_59_pdest;
        input  io_diffCommits_info_59_rfWen;
        input  io_diffCommits_info_59_fpWen;
        input  io_diffCommits_info_59_vecWen;
        input  io_diffCommits_info_59_v0Wen;
        input  io_diffCommits_info_59_vlWen;
        input  io_diffCommits_info_60_ldest;
        input  io_diffCommits_info_60_pdest;
        input  io_diffCommits_info_60_rfWen;
        input  io_diffCommits_info_60_fpWen;
        input  io_diffCommits_info_60_vecWen;
        input  io_diffCommits_info_60_v0Wen;
        input  io_diffCommits_info_60_vlWen;
        input  io_diffCommits_info_61_ldest;
        input  io_diffCommits_info_61_pdest;
        input  io_diffCommits_info_61_rfWen;
        input  io_diffCommits_info_61_fpWen;
        input  io_diffCommits_info_61_vecWen;
        input  io_diffCommits_info_61_v0Wen;
        input  io_diffCommits_info_61_vlWen;
        input  io_diffCommits_info_62_ldest;
        input  io_diffCommits_info_62_pdest;
        input  io_diffCommits_info_62_rfWen;
        input  io_diffCommits_info_62_fpWen;
        input  io_diffCommits_info_62_vecWen;
        input  io_diffCommits_info_62_v0Wen;
        input  io_diffCommits_info_62_vlWen;
        input  io_diffCommits_info_63_ldest;
        input  io_diffCommits_info_63_pdest;
        input  io_diffCommits_info_63_rfWen;
        input  io_diffCommits_info_63_fpWen;
        input  io_diffCommits_info_63_vecWen;
        input  io_diffCommits_info_63_v0Wen;
        input  io_diffCommits_info_63_vlWen;
        input  io_diffCommits_info_64_ldest;
        input  io_diffCommits_info_64_pdest;
        input  io_diffCommits_info_64_rfWen;
        input  io_diffCommits_info_64_fpWen;
        input  io_diffCommits_info_64_vecWen;
        input  io_diffCommits_info_64_v0Wen;
        input  io_diffCommits_info_64_vlWen;
        input  io_diffCommits_info_65_ldest;
        input  io_diffCommits_info_65_pdest;
        input  io_diffCommits_info_65_rfWen;
        input  io_diffCommits_info_65_fpWen;
        input  io_diffCommits_info_65_vecWen;
        input  io_diffCommits_info_65_v0Wen;
        input  io_diffCommits_info_65_vlWen;
        input  io_diffCommits_info_66_ldest;
        input  io_diffCommits_info_66_pdest;
        input  io_diffCommits_info_66_rfWen;
        input  io_diffCommits_info_66_fpWen;
        input  io_diffCommits_info_66_vecWen;
        input  io_diffCommits_info_66_v0Wen;
        input  io_diffCommits_info_66_vlWen;
        input  io_diffCommits_info_67_ldest;
        input  io_diffCommits_info_67_pdest;
        input  io_diffCommits_info_67_rfWen;
        input  io_diffCommits_info_67_fpWen;
        input  io_diffCommits_info_67_vecWen;
        input  io_diffCommits_info_67_v0Wen;
        input  io_diffCommits_info_67_vlWen;
        input  io_diffCommits_info_68_ldest;
        input  io_diffCommits_info_68_pdest;
        input  io_diffCommits_info_68_rfWen;
        input  io_diffCommits_info_68_fpWen;
        input  io_diffCommits_info_68_vecWen;
        input  io_diffCommits_info_68_v0Wen;
        input  io_diffCommits_info_68_vlWen;
        input  io_diffCommits_info_69_ldest;
        input  io_diffCommits_info_69_pdest;
        input  io_diffCommits_info_69_rfWen;
        input  io_diffCommits_info_69_fpWen;
        input  io_diffCommits_info_69_vecWen;
        input  io_diffCommits_info_69_v0Wen;
        input  io_diffCommits_info_69_vlWen;
        input  io_diffCommits_info_70_ldest;
        input  io_diffCommits_info_70_pdest;
        input  io_diffCommits_info_70_rfWen;
        input  io_diffCommits_info_70_fpWen;
        input  io_diffCommits_info_70_vecWen;
        input  io_diffCommits_info_70_v0Wen;
        input  io_diffCommits_info_70_vlWen;
        input  io_diffCommits_info_71_ldest;
        input  io_diffCommits_info_71_pdest;
        input  io_diffCommits_info_71_rfWen;
        input  io_diffCommits_info_71_fpWen;
        input  io_diffCommits_info_71_vecWen;
        input  io_diffCommits_info_71_v0Wen;
        input  io_diffCommits_info_71_vlWen;
        input  io_diffCommits_info_72_ldest;
        input  io_diffCommits_info_72_pdest;
        input  io_diffCommits_info_72_rfWen;
        input  io_diffCommits_info_72_fpWen;
        input  io_diffCommits_info_72_vecWen;
        input  io_diffCommits_info_72_v0Wen;
        input  io_diffCommits_info_72_vlWen;
        input  io_diffCommits_info_73_ldest;
        input  io_diffCommits_info_73_pdest;
        input  io_diffCommits_info_73_rfWen;
        input  io_diffCommits_info_73_fpWen;
        input  io_diffCommits_info_73_vecWen;
        input  io_diffCommits_info_73_v0Wen;
        input  io_diffCommits_info_73_vlWen;
        input  io_diffCommits_info_74_ldest;
        input  io_diffCommits_info_74_pdest;
        input  io_diffCommits_info_74_rfWen;
        input  io_diffCommits_info_74_fpWen;
        input  io_diffCommits_info_74_vecWen;
        input  io_diffCommits_info_74_v0Wen;
        input  io_diffCommits_info_74_vlWen;
        input  io_diffCommits_info_75_ldest;
        input  io_diffCommits_info_75_pdest;
        input  io_diffCommits_info_75_rfWen;
        input  io_diffCommits_info_75_fpWen;
        input  io_diffCommits_info_75_vecWen;
        input  io_diffCommits_info_75_v0Wen;
        input  io_diffCommits_info_75_vlWen;
        input  io_diffCommits_info_76_ldest;
        input  io_diffCommits_info_76_pdest;
        input  io_diffCommits_info_76_rfWen;
        input  io_diffCommits_info_76_fpWen;
        input  io_diffCommits_info_76_vecWen;
        input  io_diffCommits_info_76_v0Wen;
        input  io_diffCommits_info_76_vlWen;
        input  io_diffCommits_info_77_ldest;
        input  io_diffCommits_info_77_pdest;
        input  io_diffCommits_info_77_rfWen;
        input  io_diffCommits_info_77_fpWen;
        input  io_diffCommits_info_77_vecWen;
        input  io_diffCommits_info_77_v0Wen;
        input  io_diffCommits_info_77_vlWen;
        input  io_diffCommits_info_78_ldest;
        input  io_diffCommits_info_78_pdest;
        input  io_diffCommits_info_78_rfWen;
        input  io_diffCommits_info_78_fpWen;
        input  io_diffCommits_info_78_vecWen;
        input  io_diffCommits_info_78_v0Wen;
        input  io_diffCommits_info_78_vlWen;
        input  io_diffCommits_info_79_ldest;
        input  io_diffCommits_info_79_pdest;
        input  io_diffCommits_info_79_rfWen;
        input  io_diffCommits_info_79_fpWen;
        input  io_diffCommits_info_79_vecWen;
        input  io_diffCommits_info_79_v0Wen;
        input  io_diffCommits_info_79_vlWen;
        input  io_diffCommits_info_80_ldest;
        input  io_diffCommits_info_80_pdest;
        input  io_diffCommits_info_80_rfWen;
        input  io_diffCommits_info_80_fpWen;
        input  io_diffCommits_info_80_vecWen;
        input  io_diffCommits_info_80_v0Wen;
        input  io_diffCommits_info_80_vlWen;
        input  io_diffCommits_info_81_ldest;
        input  io_diffCommits_info_81_pdest;
        input  io_diffCommits_info_81_rfWen;
        input  io_diffCommits_info_81_fpWen;
        input  io_diffCommits_info_81_vecWen;
        input  io_diffCommits_info_81_v0Wen;
        input  io_diffCommits_info_81_vlWen;
        input  io_diffCommits_info_82_ldest;
        input  io_diffCommits_info_82_pdest;
        input  io_diffCommits_info_82_rfWen;
        input  io_diffCommits_info_82_fpWen;
        input  io_diffCommits_info_82_vecWen;
        input  io_diffCommits_info_82_v0Wen;
        input  io_diffCommits_info_82_vlWen;
        input  io_diffCommits_info_83_ldest;
        input  io_diffCommits_info_83_pdest;
        input  io_diffCommits_info_83_rfWen;
        input  io_diffCommits_info_83_fpWen;
        input  io_diffCommits_info_83_vecWen;
        input  io_diffCommits_info_83_v0Wen;
        input  io_diffCommits_info_83_vlWen;
        input  io_diffCommits_info_84_ldest;
        input  io_diffCommits_info_84_pdest;
        input  io_diffCommits_info_84_rfWen;
        input  io_diffCommits_info_84_fpWen;
        input  io_diffCommits_info_84_vecWen;
        input  io_diffCommits_info_84_v0Wen;
        input  io_diffCommits_info_84_vlWen;
        input  io_diffCommits_info_85_ldest;
        input  io_diffCommits_info_85_pdest;
        input  io_diffCommits_info_85_rfWen;
        input  io_diffCommits_info_85_fpWen;
        input  io_diffCommits_info_85_vecWen;
        input  io_diffCommits_info_85_v0Wen;
        input  io_diffCommits_info_85_vlWen;
        input  io_diffCommits_info_86_ldest;
        input  io_diffCommits_info_86_pdest;
        input  io_diffCommits_info_86_rfWen;
        input  io_diffCommits_info_86_fpWen;
        input  io_diffCommits_info_86_vecWen;
        input  io_diffCommits_info_86_v0Wen;
        input  io_diffCommits_info_86_vlWen;
        input  io_diffCommits_info_87_ldest;
        input  io_diffCommits_info_87_pdest;
        input  io_diffCommits_info_87_rfWen;
        input  io_diffCommits_info_87_fpWen;
        input  io_diffCommits_info_87_vecWen;
        input  io_diffCommits_info_87_v0Wen;
        input  io_diffCommits_info_87_vlWen;
        input  io_diffCommits_info_88_ldest;
        input  io_diffCommits_info_88_pdest;
        input  io_diffCommits_info_88_rfWen;
        input  io_diffCommits_info_88_fpWen;
        input  io_diffCommits_info_88_vecWen;
        input  io_diffCommits_info_88_v0Wen;
        input  io_diffCommits_info_88_vlWen;
        input  io_diffCommits_info_89_ldest;
        input  io_diffCommits_info_89_pdest;
        input  io_diffCommits_info_89_rfWen;
        input  io_diffCommits_info_89_fpWen;
        input  io_diffCommits_info_89_vecWen;
        input  io_diffCommits_info_89_v0Wen;
        input  io_diffCommits_info_89_vlWen;
        input  io_diffCommits_info_90_ldest;
        input  io_diffCommits_info_90_pdest;
        input  io_diffCommits_info_90_rfWen;
        input  io_diffCommits_info_90_fpWen;
        input  io_diffCommits_info_90_vecWen;
        input  io_diffCommits_info_90_v0Wen;
        input  io_diffCommits_info_90_vlWen;
        input  io_diffCommits_info_91_ldest;
        input  io_diffCommits_info_91_pdest;
        input  io_diffCommits_info_91_rfWen;
        input  io_diffCommits_info_91_fpWen;
        input  io_diffCommits_info_91_vecWen;
        input  io_diffCommits_info_91_v0Wen;
        input  io_diffCommits_info_91_vlWen;
        input  io_diffCommits_info_92_ldest;
        input  io_diffCommits_info_92_pdest;
        input  io_diffCommits_info_92_rfWen;
        input  io_diffCommits_info_92_fpWen;
        input  io_diffCommits_info_92_vecWen;
        input  io_diffCommits_info_92_v0Wen;
        input  io_diffCommits_info_92_vlWen;
        input  io_diffCommits_info_93_ldest;
        input  io_diffCommits_info_93_pdest;
        input  io_diffCommits_info_93_rfWen;
        input  io_diffCommits_info_93_fpWen;
        input  io_diffCommits_info_93_vecWen;
        input  io_diffCommits_info_93_v0Wen;
        input  io_diffCommits_info_93_vlWen;
        input  io_diffCommits_info_94_ldest;
        input  io_diffCommits_info_94_pdest;
        input  io_diffCommits_info_94_rfWen;
        input  io_diffCommits_info_94_fpWen;
        input  io_diffCommits_info_94_vecWen;
        input  io_diffCommits_info_94_v0Wen;
        input  io_diffCommits_info_94_vlWen;
        input  io_diffCommits_info_95_ldest;
        input  io_diffCommits_info_95_pdest;
        input  io_diffCommits_info_95_rfWen;
        input  io_diffCommits_info_95_fpWen;
        input  io_diffCommits_info_95_vecWen;
        input  io_diffCommits_info_95_v0Wen;
        input  io_diffCommits_info_95_vlWen;
        input  io_diffCommits_info_96_ldest;
        input  io_diffCommits_info_96_pdest;
        input  io_diffCommits_info_96_rfWen;
        input  io_diffCommits_info_96_fpWen;
        input  io_diffCommits_info_96_vecWen;
        input  io_diffCommits_info_96_v0Wen;
        input  io_diffCommits_info_96_vlWen;
        input  io_diffCommits_info_97_ldest;
        input  io_diffCommits_info_97_pdest;
        input  io_diffCommits_info_97_rfWen;
        input  io_diffCommits_info_97_fpWen;
        input  io_diffCommits_info_97_vecWen;
        input  io_diffCommits_info_97_v0Wen;
        input  io_diffCommits_info_97_vlWen;
        input  io_diffCommits_info_98_ldest;
        input  io_diffCommits_info_98_pdest;
        input  io_diffCommits_info_98_rfWen;
        input  io_diffCommits_info_98_fpWen;
        input  io_diffCommits_info_98_vecWen;
        input  io_diffCommits_info_98_v0Wen;
        input  io_diffCommits_info_98_vlWen;
        input  io_diffCommits_info_99_ldest;
        input  io_diffCommits_info_99_pdest;
        input  io_diffCommits_info_99_rfWen;
        input  io_diffCommits_info_99_fpWen;
        input  io_diffCommits_info_99_vecWen;
        input  io_diffCommits_info_99_v0Wen;
        input  io_diffCommits_info_99_vlWen;
        input  io_diffCommits_info_100_ldest;
        input  io_diffCommits_info_100_pdest;
        input  io_diffCommits_info_100_rfWen;
        input  io_diffCommits_info_100_fpWen;
        input  io_diffCommits_info_100_vecWen;
        input  io_diffCommits_info_100_v0Wen;
        input  io_diffCommits_info_100_vlWen;
        input  io_diffCommits_info_101_ldest;
        input  io_diffCommits_info_101_pdest;
        input  io_diffCommits_info_101_rfWen;
        input  io_diffCommits_info_101_fpWen;
        input  io_diffCommits_info_101_vecWen;
        input  io_diffCommits_info_101_v0Wen;
        input  io_diffCommits_info_101_vlWen;
        input  io_diffCommits_info_102_ldest;
        input  io_diffCommits_info_102_pdest;
        input  io_diffCommits_info_102_rfWen;
        input  io_diffCommits_info_102_fpWen;
        input  io_diffCommits_info_102_vecWen;
        input  io_diffCommits_info_102_v0Wen;
        input  io_diffCommits_info_102_vlWen;
        input  io_diffCommits_info_103_ldest;
        input  io_diffCommits_info_103_pdest;
        input  io_diffCommits_info_103_rfWen;
        input  io_diffCommits_info_103_fpWen;
        input  io_diffCommits_info_103_vecWen;
        input  io_diffCommits_info_103_v0Wen;
        input  io_diffCommits_info_103_vlWen;
        input  io_diffCommits_info_104_ldest;
        input  io_diffCommits_info_104_pdest;
        input  io_diffCommits_info_104_rfWen;
        input  io_diffCommits_info_104_fpWen;
        input  io_diffCommits_info_104_vecWen;
        input  io_diffCommits_info_104_v0Wen;
        input  io_diffCommits_info_104_vlWen;
        input  io_diffCommits_info_105_ldest;
        input  io_diffCommits_info_105_pdest;
        input  io_diffCommits_info_105_rfWen;
        input  io_diffCommits_info_105_fpWen;
        input  io_diffCommits_info_105_vecWen;
        input  io_diffCommits_info_105_v0Wen;
        input  io_diffCommits_info_105_vlWen;
        input  io_diffCommits_info_106_ldest;
        input  io_diffCommits_info_106_pdest;
        input  io_diffCommits_info_106_rfWen;
        input  io_diffCommits_info_106_fpWen;
        input  io_diffCommits_info_106_vecWen;
        input  io_diffCommits_info_106_v0Wen;
        input  io_diffCommits_info_106_vlWen;
        input  io_diffCommits_info_107_ldest;
        input  io_diffCommits_info_107_pdest;
        input  io_diffCommits_info_107_rfWen;
        input  io_diffCommits_info_107_fpWen;
        input  io_diffCommits_info_107_vecWen;
        input  io_diffCommits_info_107_v0Wen;
        input  io_diffCommits_info_107_vlWen;
        input  io_diffCommits_info_108_ldest;
        input  io_diffCommits_info_108_pdest;
        input  io_diffCommits_info_108_rfWen;
        input  io_diffCommits_info_108_fpWen;
        input  io_diffCommits_info_108_vecWen;
        input  io_diffCommits_info_108_v0Wen;
        input  io_diffCommits_info_108_vlWen;
        input  io_diffCommits_info_109_ldest;
        input  io_diffCommits_info_109_pdest;
        input  io_diffCommits_info_109_rfWen;
        input  io_diffCommits_info_109_fpWen;
        input  io_diffCommits_info_109_vecWen;
        input  io_diffCommits_info_109_v0Wen;
        input  io_diffCommits_info_109_vlWen;
        input  io_diffCommits_info_110_ldest;
        input  io_diffCommits_info_110_pdest;
        input  io_diffCommits_info_110_rfWen;
        input  io_diffCommits_info_110_fpWen;
        input  io_diffCommits_info_110_vecWen;
        input  io_diffCommits_info_110_v0Wen;
        input  io_diffCommits_info_110_vlWen;
        input  io_diffCommits_info_111_ldest;
        input  io_diffCommits_info_111_pdest;
        input  io_diffCommits_info_111_rfWen;
        input  io_diffCommits_info_111_fpWen;
        input  io_diffCommits_info_111_vecWen;
        input  io_diffCommits_info_111_v0Wen;
        input  io_diffCommits_info_111_vlWen;
        input  io_diffCommits_info_112_ldest;
        input  io_diffCommits_info_112_pdest;
        input  io_diffCommits_info_112_rfWen;
        input  io_diffCommits_info_112_fpWen;
        input  io_diffCommits_info_112_vecWen;
        input  io_diffCommits_info_112_v0Wen;
        input  io_diffCommits_info_112_vlWen;
        input  io_diffCommits_info_113_ldest;
        input  io_diffCommits_info_113_pdest;
        input  io_diffCommits_info_113_rfWen;
        input  io_diffCommits_info_113_fpWen;
        input  io_diffCommits_info_113_vecWen;
        input  io_diffCommits_info_113_v0Wen;
        input  io_diffCommits_info_113_vlWen;
        input  io_diffCommits_info_114_ldest;
        input  io_diffCommits_info_114_pdest;
        input  io_diffCommits_info_114_rfWen;
        input  io_diffCommits_info_114_fpWen;
        input  io_diffCommits_info_114_vecWen;
        input  io_diffCommits_info_114_v0Wen;
        input  io_diffCommits_info_114_vlWen;
        input  io_diffCommits_info_115_ldest;
        input  io_diffCommits_info_115_pdest;
        input  io_diffCommits_info_115_rfWen;
        input  io_diffCommits_info_115_fpWen;
        input  io_diffCommits_info_115_vecWen;
        input  io_diffCommits_info_115_v0Wen;
        input  io_diffCommits_info_115_vlWen;
        input  io_diffCommits_info_116_ldest;
        input  io_diffCommits_info_116_pdest;
        input  io_diffCommits_info_116_rfWen;
        input  io_diffCommits_info_116_fpWen;
        input  io_diffCommits_info_116_vecWen;
        input  io_diffCommits_info_116_v0Wen;
        input  io_diffCommits_info_116_vlWen;
        input  io_diffCommits_info_117_ldest;
        input  io_diffCommits_info_117_pdest;
        input  io_diffCommits_info_117_rfWen;
        input  io_diffCommits_info_117_fpWen;
        input  io_diffCommits_info_117_vecWen;
        input  io_diffCommits_info_117_v0Wen;
        input  io_diffCommits_info_117_vlWen;
        input  io_diffCommits_info_118_ldest;
        input  io_diffCommits_info_118_pdest;
        input  io_diffCommits_info_118_rfWen;
        input  io_diffCommits_info_118_fpWen;
        input  io_diffCommits_info_118_vecWen;
        input  io_diffCommits_info_118_v0Wen;
        input  io_diffCommits_info_118_vlWen;
        input  io_diffCommits_info_119_ldest;
        input  io_diffCommits_info_119_pdest;
        input  io_diffCommits_info_119_rfWen;
        input  io_diffCommits_info_119_fpWen;
        input  io_diffCommits_info_119_vecWen;
        input  io_diffCommits_info_119_v0Wen;
        input  io_diffCommits_info_119_vlWen;
        input  io_diffCommits_info_120_ldest;
        input  io_diffCommits_info_120_pdest;
        input  io_diffCommits_info_120_rfWen;
        input  io_diffCommits_info_120_fpWen;
        input  io_diffCommits_info_120_vecWen;
        input  io_diffCommits_info_120_v0Wen;
        input  io_diffCommits_info_120_vlWen;
        input  io_diffCommits_info_121_ldest;
        input  io_diffCommits_info_121_pdest;
        input  io_diffCommits_info_121_rfWen;
        input  io_diffCommits_info_121_fpWen;
        input  io_diffCommits_info_121_vecWen;
        input  io_diffCommits_info_121_v0Wen;
        input  io_diffCommits_info_121_vlWen;
        input  io_diffCommits_info_122_ldest;
        input  io_diffCommits_info_122_pdest;
        input  io_diffCommits_info_122_rfWen;
        input  io_diffCommits_info_122_fpWen;
        input  io_diffCommits_info_122_vecWen;
        input  io_diffCommits_info_122_v0Wen;
        input  io_diffCommits_info_122_vlWen;
        input  io_diffCommits_info_123_ldest;
        input  io_diffCommits_info_123_pdest;
        input  io_diffCommits_info_123_rfWen;
        input  io_diffCommits_info_123_fpWen;
        input  io_diffCommits_info_123_vecWen;
        input  io_diffCommits_info_123_v0Wen;
        input  io_diffCommits_info_123_vlWen;
        input  io_diffCommits_info_124_ldest;
        input  io_diffCommits_info_124_pdest;
        input  io_diffCommits_info_124_rfWen;
        input  io_diffCommits_info_124_fpWen;
        input  io_diffCommits_info_124_vecWen;
        input  io_diffCommits_info_124_v0Wen;
        input  io_diffCommits_info_124_vlWen;
        input  io_diffCommits_info_125_ldest;
        input  io_diffCommits_info_125_pdest;
        input  io_diffCommits_info_125_rfWen;
        input  io_diffCommits_info_125_fpWen;
        input  io_diffCommits_info_125_vecWen;
        input  io_diffCommits_info_125_v0Wen;
        input  io_diffCommits_info_125_vlWen;
        input  io_diffCommits_info_126_ldest;
        input  io_diffCommits_info_126_pdest;
        input  io_diffCommits_info_126_rfWen;
        input  io_diffCommits_info_126_fpWen;
        input  io_diffCommits_info_126_vecWen;
        input  io_diffCommits_info_126_v0Wen;
        input  io_diffCommits_info_126_vlWen;
        input  io_diffCommits_info_127_ldest;
        input  io_diffCommits_info_127_pdest;
        input  io_diffCommits_info_127_rfWen;
        input  io_diffCommits_info_127_fpWen;
        input  io_diffCommits_info_127_vecWen;
        input  io_diffCommits_info_127_v0Wen;
        input  io_diffCommits_info_127_vlWen;
        input  io_diffCommits_info_128_ldest;
        input  io_diffCommits_info_128_pdest;
        input  io_diffCommits_info_128_rfWen;
        input  io_diffCommits_info_128_fpWen;
        input  io_diffCommits_info_128_vecWen;
        input  io_diffCommits_info_128_v0Wen;
        input  io_diffCommits_info_128_vlWen;
        input  io_diffCommits_info_129_ldest;
        input  io_diffCommits_info_129_pdest;
        input  io_diffCommits_info_129_rfWen;
        input  io_diffCommits_info_129_fpWen;
        input  io_diffCommits_info_129_vecWen;
        input  io_diffCommits_info_129_v0Wen;
        input  io_diffCommits_info_129_vlWen;
        input  io_diffCommits_info_130_ldest;
        input  io_diffCommits_info_130_pdest;
        input  io_diffCommits_info_130_rfWen;
        input  io_diffCommits_info_130_fpWen;
        input  io_diffCommits_info_130_vecWen;
        input  io_diffCommits_info_130_v0Wen;
        input  io_diffCommits_info_130_vlWen;
        input  io_diffCommits_info_131_ldest;
        input  io_diffCommits_info_131_pdest;
        input  io_diffCommits_info_131_rfWen;
        input  io_diffCommits_info_131_fpWen;
        input  io_diffCommits_info_131_vecWen;
        input  io_diffCommits_info_131_v0Wen;
        input  io_diffCommits_info_131_vlWen;
        input  io_diffCommits_info_132_ldest;
        input  io_diffCommits_info_132_pdest;
        input  io_diffCommits_info_132_rfWen;
        input  io_diffCommits_info_132_fpWen;
        input  io_diffCommits_info_132_vecWen;
        input  io_diffCommits_info_132_v0Wen;
        input  io_diffCommits_info_132_vlWen;
        input  io_diffCommits_info_133_ldest;
        input  io_diffCommits_info_133_pdest;
        input  io_diffCommits_info_133_rfWen;
        input  io_diffCommits_info_133_fpWen;
        input  io_diffCommits_info_133_vecWen;
        input  io_diffCommits_info_133_v0Wen;
        input  io_diffCommits_info_133_vlWen;
        input  io_diffCommits_info_134_ldest;
        input  io_diffCommits_info_134_pdest;
        input  io_diffCommits_info_134_rfWen;
        input  io_diffCommits_info_134_fpWen;
        input  io_diffCommits_info_134_vecWen;
        input  io_diffCommits_info_134_v0Wen;
        input  io_diffCommits_info_134_vlWen;
        input  io_diffCommits_info_135_ldest;
        input  io_diffCommits_info_135_pdest;
        input  io_diffCommits_info_135_rfWen;
        input  io_diffCommits_info_135_fpWen;
        input  io_diffCommits_info_135_vecWen;
        input  io_diffCommits_info_135_v0Wen;
        input  io_diffCommits_info_135_vlWen;
        input  io_diffCommits_info_136_ldest;
        input  io_diffCommits_info_136_pdest;
        input  io_diffCommits_info_136_rfWen;
        input  io_diffCommits_info_136_fpWen;
        input  io_diffCommits_info_136_vecWen;
        input  io_diffCommits_info_136_v0Wen;
        input  io_diffCommits_info_136_vlWen;
        input  io_diffCommits_info_137_ldest;
        input  io_diffCommits_info_137_pdest;
        input  io_diffCommits_info_137_rfWen;
        input  io_diffCommits_info_137_fpWen;
        input  io_diffCommits_info_137_vecWen;
        input  io_diffCommits_info_137_v0Wen;
        input  io_diffCommits_info_137_vlWen;
        input  io_diffCommits_info_138_ldest;
        input  io_diffCommits_info_138_pdest;
        input  io_diffCommits_info_138_rfWen;
        input  io_diffCommits_info_138_fpWen;
        input  io_diffCommits_info_138_vecWen;
        input  io_diffCommits_info_138_v0Wen;
        input  io_diffCommits_info_138_vlWen;
        input  io_diffCommits_info_139_ldest;
        input  io_diffCommits_info_139_pdest;
        input  io_diffCommits_info_139_rfWen;
        input  io_diffCommits_info_139_fpWen;
        input  io_diffCommits_info_139_vecWen;
        input  io_diffCommits_info_139_v0Wen;
        input  io_diffCommits_info_139_vlWen;
        input  io_diffCommits_info_140_ldest;
        input  io_diffCommits_info_140_pdest;
        input  io_diffCommits_info_140_rfWen;
        input  io_diffCommits_info_140_fpWen;
        input  io_diffCommits_info_140_vecWen;
        input  io_diffCommits_info_140_v0Wen;
        input  io_diffCommits_info_140_vlWen;
        input  io_diffCommits_info_141_ldest;
        input  io_diffCommits_info_141_pdest;
        input  io_diffCommits_info_141_rfWen;
        input  io_diffCommits_info_141_fpWen;
        input  io_diffCommits_info_141_vecWen;
        input  io_diffCommits_info_141_v0Wen;
        input  io_diffCommits_info_141_vlWen;
        input  io_diffCommits_info_142_ldest;
        input  io_diffCommits_info_142_pdest;
        input  io_diffCommits_info_142_rfWen;
        input  io_diffCommits_info_142_fpWen;
        input  io_diffCommits_info_142_vecWen;
        input  io_diffCommits_info_142_v0Wen;
        input  io_diffCommits_info_142_vlWen;
        input  io_diffCommits_info_143_ldest;
        input  io_diffCommits_info_143_pdest;
        input  io_diffCommits_info_143_rfWen;
        input  io_diffCommits_info_143_fpWen;
        input  io_diffCommits_info_143_vecWen;
        input  io_diffCommits_info_143_v0Wen;
        input  io_diffCommits_info_143_vlWen;
        input  io_diffCommits_info_144_ldest;
        input  io_diffCommits_info_144_pdest;
        input  io_diffCommits_info_144_rfWen;
        input  io_diffCommits_info_144_fpWen;
        input  io_diffCommits_info_144_vecWen;
        input  io_diffCommits_info_144_v0Wen;
        input  io_diffCommits_info_144_vlWen;
        input  io_diffCommits_info_145_ldest;
        input  io_diffCommits_info_145_pdest;
        input  io_diffCommits_info_145_rfWen;
        input  io_diffCommits_info_145_fpWen;
        input  io_diffCommits_info_145_vecWen;
        input  io_diffCommits_info_145_v0Wen;
        input  io_diffCommits_info_145_vlWen;
        input  io_diffCommits_info_146_ldest;
        input  io_diffCommits_info_146_pdest;
        input  io_diffCommits_info_146_rfWen;
        input  io_diffCommits_info_146_fpWen;
        input  io_diffCommits_info_146_vecWen;
        input  io_diffCommits_info_146_v0Wen;
        input  io_diffCommits_info_146_vlWen;
        input  io_diffCommits_info_147_ldest;
        input  io_diffCommits_info_147_pdest;
        input  io_diffCommits_info_147_rfWen;
        input  io_diffCommits_info_147_fpWen;
        input  io_diffCommits_info_147_vecWen;
        input  io_diffCommits_info_147_v0Wen;
        input  io_diffCommits_info_147_vlWen;
        input  io_diffCommits_info_148_ldest;
        input  io_diffCommits_info_148_pdest;
        input  io_diffCommits_info_148_rfWen;
        input  io_diffCommits_info_148_fpWen;
        input  io_diffCommits_info_148_vecWen;
        input  io_diffCommits_info_148_v0Wen;
        input  io_diffCommits_info_148_vlWen;
        input  io_diffCommits_info_149_ldest;
        input  io_diffCommits_info_149_pdest;
        input  io_diffCommits_info_149_rfWen;
        input  io_diffCommits_info_149_fpWen;
        input  io_diffCommits_info_149_vecWen;
        input  io_diffCommits_info_149_v0Wen;
        input  io_diffCommits_info_149_vlWen;
        input  io_diffCommits_info_150_ldest;
        input  io_diffCommits_info_150_pdest;
        input  io_diffCommits_info_150_rfWen;
        input  io_diffCommits_info_150_fpWen;
        input  io_diffCommits_info_150_vecWen;
        input  io_diffCommits_info_150_v0Wen;
        input  io_diffCommits_info_150_vlWen;
        input  io_diffCommits_info_151_ldest;
        input  io_diffCommits_info_151_pdest;
        input  io_diffCommits_info_151_rfWen;
        input  io_diffCommits_info_151_fpWen;
        input  io_diffCommits_info_151_vecWen;
        input  io_diffCommits_info_151_v0Wen;
        input  io_diffCommits_info_151_vlWen;
        input  io_diffCommits_info_152_ldest;
        input  io_diffCommits_info_152_pdest;
        input  io_diffCommits_info_152_rfWen;
        input  io_diffCommits_info_152_fpWen;
        input  io_diffCommits_info_152_vecWen;
        input  io_diffCommits_info_152_v0Wen;
        input  io_diffCommits_info_152_vlWen;
        input  io_diffCommits_info_153_ldest;
        input  io_diffCommits_info_153_pdest;
        input  io_diffCommits_info_153_rfWen;
        input  io_diffCommits_info_153_fpWen;
        input  io_diffCommits_info_153_vecWen;
        input  io_diffCommits_info_153_v0Wen;
        input  io_diffCommits_info_153_vlWen;
        input  io_diffCommits_info_154_ldest;
        input  io_diffCommits_info_154_pdest;
        input  io_diffCommits_info_154_rfWen;
        input  io_diffCommits_info_154_fpWen;
        input  io_diffCommits_info_154_vecWen;
        input  io_diffCommits_info_154_v0Wen;
        input  io_diffCommits_info_154_vlWen;
        input  io_diffCommits_info_155_ldest;
        input  io_diffCommits_info_155_pdest;
        input  io_diffCommits_info_155_rfWen;
        input  io_diffCommits_info_155_fpWen;
        input  io_diffCommits_info_155_vecWen;
        input  io_diffCommits_info_155_v0Wen;
        input  io_diffCommits_info_155_vlWen;
        input  io_diffCommits_info_156_ldest;
        input  io_diffCommits_info_156_pdest;
        input  io_diffCommits_info_156_rfWen;
        input  io_diffCommits_info_156_fpWen;
        input  io_diffCommits_info_156_vecWen;
        input  io_diffCommits_info_156_v0Wen;
        input  io_diffCommits_info_156_vlWen;
        input  io_diffCommits_info_157_ldest;
        input  io_diffCommits_info_157_pdest;
        input  io_diffCommits_info_157_rfWen;
        input  io_diffCommits_info_157_fpWen;
        input  io_diffCommits_info_157_vecWen;
        input  io_diffCommits_info_157_v0Wen;
        input  io_diffCommits_info_157_vlWen;
        input  io_diffCommits_info_158_ldest;
        input  io_diffCommits_info_158_pdest;
        input  io_diffCommits_info_158_rfWen;
        input  io_diffCommits_info_158_fpWen;
        input  io_diffCommits_info_158_vecWen;
        input  io_diffCommits_info_158_v0Wen;
        input  io_diffCommits_info_158_vlWen;
        input  io_diffCommits_info_159_ldest;
        input  io_diffCommits_info_159_pdest;
        input  io_diffCommits_info_159_rfWen;
        input  io_diffCommits_info_159_fpWen;
        input  io_diffCommits_info_159_vecWen;
        input  io_diffCommits_info_159_v0Wen;
        input  io_diffCommits_info_159_vlWen;
        input  io_diffCommits_info_160_ldest;
        input  io_diffCommits_info_160_pdest;
        input  io_diffCommits_info_160_rfWen;
        input  io_diffCommits_info_160_fpWen;
        input  io_diffCommits_info_160_vecWen;
        input  io_diffCommits_info_160_v0Wen;
        input  io_diffCommits_info_160_vlWen;
        input  io_diffCommits_info_161_ldest;
        input  io_diffCommits_info_161_pdest;
        input  io_diffCommits_info_161_rfWen;
        input  io_diffCommits_info_161_fpWen;
        input  io_diffCommits_info_161_vecWen;
        input  io_diffCommits_info_161_v0Wen;
        input  io_diffCommits_info_161_vlWen;
        input  io_diffCommits_info_162_ldest;
        input  io_diffCommits_info_162_pdest;
        input  io_diffCommits_info_162_rfWen;
        input  io_diffCommits_info_162_fpWen;
        input  io_diffCommits_info_162_vecWen;
        input  io_diffCommits_info_162_v0Wen;
        input  io_diffCommits_info_162_vlWen;
        input  io_diffCommits_info_163_ldest;
        input  io_diffCommits_info_163_pdest;
        input  io_diffCommits_info_163_rfWen;
        input  io_diffCommits_info_163_fpWen;
        input  io_diffCommits_info_163_vecWen;
        input  io_diffCommits_info_163_v0Wen;
        input  io_diffCommits_info_163_vlWen;
        input  io_diffCommits_info_164_ldest;
        input  io_diffCommits_info_164_pdest;
        input  io_diffCommits_info_164_rfWen;
        input  io_diffCommits_info_164_fpWen;
        input  io_diffCommits_info_164_vecWen;
        input  io_diffCommits_info_164_v0Wen;
        input  io_diffCommits_info_164_vlWen;
        input  io_diffCommits_info_165_ldest;
        input  io_diffCommits_info_165_pdest;
        input  io_diffCommits_info_165_rfWen;
        input  io_diffCommits_info_165_fpWen;
        input  io_diffCommits_info_165_vecWen;
        input  io_diffCommits_info_165_v0Wen;
        input  io_diffCommits_info_165_vlWen;
        input  io_diffCommits_info_166_ldest;
        input  io_diffCommits_info_166_pdest;
        input  io_diffCommits_info_166_rfWen;
        input  io_diffCommits_info_166_fpWen;
        input  io_diffCommits_info_166_vecWen;
        input  io_diffCommits_info_166_v0Wen;
        input  io_diffCommits_info_166_vlWen;
        input  io_diffCommits_info_167_ldest;
        input  io_diffCommits_info_167_pdest;
        input  io_diffCommits_info_167_rfWen;
        input  io_diffCommits_info_167_fpWen;
        input  io_diffCommits_info_167_vecWen;
        input  io_diffCommits_info_167_v0Wen;
        input  io_diffCommits_info_167_vlWen;
        input  io_diffCommits_info_168_ldest;
        input  io_diffCommits_info_168_pdest;
        input  io_diffCommits_info_168_rfWen;
        input  io_diffCommits_info_168_fpWen;
        input  io_diffCommits_info_168_vecWen;
        input  io_diffCommits_info_168_v0Wen;
        input  io_diffCommits_info_168_vlWen;
        input  io_diffCommits_info_169_ldest;
        input  io_diffCommits_info_169_pdest;
        input  io_diffCommits_info_169_rfWen;
        input  io_diffCommits_info_169_fpWen;
        input  io_diffCommits_info_169_vecWen;
        input  io_diffCommits_info_169_v0Wen;
        input  io_diffCommits_info_169_vlWen;
        input  io_diffCommits_info_170_ldest;
        input  io_diffCommits_info_170_pdest;
        input  io_diffCommits_info_170_rfWen;
        input  io_diffCommits_info_170_fpWen;
        input  io_diffCommits_info_170_vecWen;
        input  io_diffCommits_info_170_v0Wen;
        input  io_diffCommits_info_170_vlWen;
        input  io_diffCommits_info_171_ldest;
        input  io_diffCommits_info_171_pdest;
        input  io_diffCommits_info_171_rfWen;
        input  io_diffCommits_info_171_fpWen;
        input  io_diffCommits_info_171_vecWen;
        input  io_diffCommits_info_171_v0Wen;
        input  io_diffCommits_info_171_vlWen;
        input  io_diffCommits_info_172_ldest;
        input  io_diffCommits_info_172_pdest;
        input  io_diffCommits_info_172_rfWen;
        input  io_diffCommits_info_172_fpWen;
        input  io_diffCommits_info_172_vecWen;
        input  io_diffCommits_info_172_v0Wen;
        input  io_diffCommits_info_172_vlWen;
        input  io_diffCommits_info_173_ldest;
        input  io_diffCommits_info_173_pdest;
        input  io_diffCommits_info_173_rfWen;
        input  io_diffCommits_info_173_fpWen;
        input  io_diffCommits_info_173_vecWen;
        input  io_diffCommits_info_173_v0Wen;
        input  io_diffCommits_info_173_vlWen;
        input  io_diffCommits_info_174_ldest;
        input  io_diffCommits_info_174_pdest;
        input  io_diffCommits_info_174_rfWen;
        input  io_diffCommits_info_174_fpWen;
        input  io_diffCommits_info_174_vecWen;
        input  io_diffCommits_info_174_v0Wen;
        input  io_diffCommits_info_174_vlWen;
        input  io_diffCommits_info_175_ldest;
        input  io_diffCommits_info_175_pdest;
        input  io_diffCommits_info_175_rfWen;
        input  io_diffCommits_info_175_fpWen;
        input  io_diffCommits_info_175_vecWen;
        input  io_diffCommits_info_175_v0Wen;
        input  io_diffCommits_info_175_vlWen;
        input  io_diffCommits_info_176_ldest;
        input  io_diffCommits_info_176_pdest;
        input  io_diffCommits_info_176_rfWen;
        input  io_diffCommits_info_176_fpWen;
        input  io_diffCommits_info_176_vecWen;
        input  io_diffCommits_info_176_v0Wen;
        input  io_diffCommits_info_176_vlWen;
        input  io_diffCommits_info_177_ldest;
        input  io_diffCommits_info_177_pdest;
        input  io_diffCommits_info_177_rfWen;
        input  io_diffCommits_info_177_fpWen;
        input  io_diffCommits_info_177_vecWen;
        input  io_diffCommits_info_177_v0Wen;
        input  io_diffCommits_info_177_vlWen;
        input  io_diffCommits_info_178_ldest;
        input  io_diffCommits_info_178_pdest;
        input  io_diffCommits_info_178_rfWen;
        input  io_diffCommits_info_178_fpWen;
        input  io_diffCommits_info_178_vecWen;
        input  io_diffCommits_info_178_v0Wen;
        input  io_diffCommits_info_178_vlWen;
        input  io_diffCommits_info_179_ldest;
        input  io_diffCommits_info_179_pdest;
        input  io_diffCommits_info_179_rfWen;
        input  io_diffCommits_info_179_fpWen;
        input  io_diffCommits_info_179_vecWen;
        input  io_diffCommits_info_179_v0Wen;
        input  io_diffCommits_info_179_vlWen;
        input  io_diffCommits_info_180_ldest;
        input  io_diffCommits_info_180_pdest;
        input  io_diffCommits_info_180_rfWen;
        input  io_diffCommits_info_180_fpWen;
        input  io_diffCommits_info_180_vecWen;
        input  io_diffCommits_info_180_v0Wen;
        input  io_diffCommits_info_180_vlWen;
        input  io_diffCommits_info_181_ldest;
        input  io_diffCommits_info_181_pdest;
        input  io_diffCommits_info_181_rfWen;
        input  io_diffCommits_info_181_fpWen;
        input  io_diffCommits_info_181_vecWen;
        input  io_diffCommits_info_181_v0Wen;
        input  io_diffCommits_info_181_vlWen;
        input  io_diffCommits_info_182_ldest;
        input  io_diffCommits_info_182_pdest;
        input  io_diffCommits_info_182_rfWen;
        input  io_diffCommits_info_182_fpWen;
        input  io_diffCommits_info_182_vecWen;
        input  io_diffCommits_info_182_v0Wen;
        input  io_diffCommits_info_182_vlWen;
        input  io_diffCommits_info_183_ldest;
        input  io_diffCommits_info_183_pdest;
        input  io_diffCommits_info_183_rfWen;
        input  io_diffCommits_info_183_fpWen;
        input  io_diffCommits_info_183_vecWen;
        input  io_diffCommits_info_183_v0Wen;
        input  io_diffCommits_info_183_vlWen;
        input  io_diffCommits_info_184_ldest;
        input  io_diffCommits_info_184_pdest;
        input  io_diffCommits_info_184_rfWen;
        input  io_diffCommits_info_184_fpWen;
        input  io_diffCommits_info_184_vecWen;
        input  io_diffCommits_info_184_v0Wen;
        input  io_diffCommits_info_184_vlWen;
        input  io_diffCommits_info_185_ldest;
        input  io_diffCommits_info_185_pdest;
        input  io_diffCommits_info_185_rfWen;
        input  io_diffCommits_info_185_fpWen;
        input  io_diffCommits_info_185_vecWen;
        input  io_diffCommits_info_185_v0Wen;
        input  io_diffCommits_info_185_vlWen;
        input  io_diffCommits_info_186_ldest;
        input  io_diffCommits_info_186_pdest;
        input  io_diffCommits_info_186_rfWen;
        input  io_diffCommits_info_186_fpWen;
        input  io_diffCommits_info_186_vecWen;
        input  io_diffCommits_info_186_v0Wen;
        input  io_diffCommits_info_186_vlWen;
        input  io_diffCommits_info_187_ldest;
        input  io_diffCommits_info_187_pdest;
        input  io_diffCommits_info_187_rfWen;
        input  io_diffCommits_info_187_fpWen;
        input  io_diffCommits_info_187_vecWen;
        input  io_diffCommits_info_187_v0Wen;
        input  io_diffCommits_info_187_vlWen;
        input  io_diffCommits_info_188_ldest;
        input  io_diffCommits_info_188_pdest;
        input  io_diffCommits_info_188_rfWen;
        input  io_diffCommits_info_188_fpWen;
        input  io_diffCommits_info_188_vecWen;
        input  io_diffCommits_info_188_v0Wen;
        input  io_diffCommits_info_188_vlWen;
        input  io_diffCommits_info_189_ldest;
        input  io_diffCommits_info_189_pdest;
        input  io_diffCommits_info_189_rfWen;
        input  io_diffCommits_info_189_fpWen;
        input  io_diffCommits_info_189_vecWen;
        input  io_diffCommits_info_189_v0Wen;
        input  io_diffCommits_info_189_vlWen;
        input  io_diffCommits_info_190_ldest;
        input  io_diffCommits_info_190_pdest;
        input  io_diffCommits_info_190_rfWen;
        input  io_diffCommits_info_190_fpWen;
        input  io_diffCommits_info_190_vecWen;
        input  io_diffCommits_info_190_v0Wen;
        input  io_diffCommits_info_190_vlWen;
        input  io_diffCommits_info_191_ldest;
        input  io_diffCommits_info_191_pdest;
        input  io_diffCommits_info_191_rfWen;
        input  io_diffCommits_info_191_fpWen;
        input  io_diffCommits_info_191_vecWen;
        input  io_diffCommits_info_191_v0Wen;
        input  io_diffCommits_info_191_vlWen;
        input  io_diffCommits_info_192_ldest;
        input  io_diffCommits_info_192_pdest;
        input  io_diffCommits_info_192_rfWen;
        input  io_diffCommits_info_192_fpWen;
        input  io_diffCommits_info_192_vecWen;
        input  io_diffCommits_info_192_v0Wen;
        input  io_diffCommits_info_192_vlWen;
        input  io_diffCommits_info_193_ldest;
        input  io_diffCommits_info_193_pdest;
        input  io_diffCommits_info_193_rfWen;
        input  io_diffCommits_info_193_fpWen;
        input  io_diffCommits_info_193_vecWen;
        input  io_diffCommits_info_193_v0Wen;
        input  io_diffCommits_info_193_vlWen;
        input  io_diffCommits_info_194_ldest;
        input  io_diffCommits_info_194_pdest;
        input  io_diffCommits_info_194_rfWen;
        input  io_diffCommits_info_194_fpWen;
        input  io_diffCommits_info_194_vecWen;
        input  io_diffCommits_info_194_v0Wen;
        input  io_diffCommits_info_194_vlWen;
        input  io_diffCommits_info_195_ldest;
        input  io_diffCommits_info_195_pdest;
        input  io_diffCommits_info_195_rfWen;
        input  io_diffCommits_info_195_fpWen;
        input  io_diffCommits_info_195_vecWen;
        input  io_diffCommits_info_195_v0Wen;
        input  io_diffCommits_info_195_vlWen;
        input  io_diffCommits_info_196_ldest;
        input  io_diffCommits_info_196_pdest;
        input  io_diffCommits_info_196_rfWen;
        input  io_diffCommits_info_196_fpWen;
        input  io_diffCommits_info_196_vecWen;
        input  io_diffCommits_info_196_v0Wen;
        input  io_diffCommits_info_196_vlWen;
        input  io_diffCommits_info_197_ldest;
        input  io_diffCommits_info_197_pdest;
        input  io_diffCommits_info_197_rfWen;
        input  io_diffCommits_info_197_fpWen;
        input  io_diffCommits_info_197_vecWen;
        input  io_diffCommits_info_197_v0Wen;
        input  io_diffCommits_info_197_vlWen;
        input  io_diffCommits_info_198_ldest;
        input  io_diffCommits_info_198_pdest;
        input  io_diffCommits_info_198_rfWen;
        input  io_diffCommits_info_198_fpWen;
        input  io_diffCommits_info_198_vecWen;
        input  io_diffCommits_info_198_v0Wen;
        input  io_diffCommits_info_198_vlWen;
        input  io_diffCommits_info_199_ldest;
        input  io_diffCommits_info_199_pdest;
        input  io_diffCommits_info_199_rfWen;
        input  io_diffCommits_info_199_fpWen;
        input  io_diffCommits_info_199_vecWen;
        input  io_diffCommits_info_199_v0Wen;
        input  io_diffCommits_info_199_vlWen;
        input  io_diffCommits_info_200_ldest;
        input  io_diffCommits_info_200_pdest;
        input  io_diffCommits_info_200_rfWen;
        input  io_diffCommits_info_200_fpWen;
        input  io_diffCommits_info_200_vecWen;
        input  io_diffCommits_info_200_v0Wen;
        input  io_diffCommits_info_200_vlWen;
        input  io_diffCommits_info_201_ldest;
        input  io_diffCommits_info_201_pdest;
        input  io_diffCommits_info_201_rfWen;
        input  io_diffCommits_info_201_fpWen;
        input  io_diffCommits_info_201_vecWen;
        input  io_diffCommits_info_201_v0Wen;
        input  io_diffCommits_info_201_vlWen;
        input  io_diffCommits_info_202_ldest;
        input  io_diffCommits_info_202_pdest;
        input  io_diffCommits_info_202_rfWen;
        input  io_diffCommits_info_202_fpWen;
        input  io_diffCommits_info_202_vecWen;
        input  io_diffCommits_info_202_v0Wen;
        input  io_diffCommits_info_202_vlWen;
        input  io_diffCommits_info_203_ldest;
        input  io_diffCommits_info_203_pdest;
        input  io_diffCommits_info_203_rfWen;
        input  io_diffCommits_info_203_fpWen;
        input  io_diffCommits_info_203_vecWen;
        input  io_diffCommits_info_203_v0Wen;
        input  io_diffCommits_info_203_vlWen;
        input  io_diffCommits_info_204_ldest;
        input  io_diffCommits_info_204_pdest;
        input  io_diffCommits_info_204_rfWen;
        input  io_diffCommits_info_204_fpWen;
        input  io_diffCommits_info_204_vecWen;
        input  io_diffCommits_info_204_v0Wen;
        input  io_diffCommits_info_204_vlWen;
        input  io_diffCommits_info_205_ldest;
        input  io_diffCommits_info_205_pdest;
        input  io_diffCommits_info_205_rfWen;
        input  io_diffCommits_info_205_fpWen;
        input  io_diffCommits_info_205_vecWen;
        input  io_diffCommits_info_205_v0Wen;
        input  io_diffCommits_info_205_vlWen;
        input  io_diffCommits_info_206_ldest;
        input  io_diffCommits_info_206_pdest;
        input  io_diffCommits_info_206_rfWen;
        input  io_diffCommits_info_206_fpWen;
        input  io_diffCommits_info_206_vecWen;
        input  io_diffCommits_info_206_v0Wen;
        input  io_diffCommits_info_206_vlWen;
        input  io_diffCommits_info_207_ldest;
        input  io_diffCommits_info_207_pdest;
        input  io_diffCommits_info_207_rfWen;
        input  io_diffCommits_info_207_fpWen;
        input  io_diffCommits_info_207_vecWen;
        input  io_diffCommits_info_207_v0Wen;
        input  io_diffCommits_info_207_vlWen;
        input  io_diffCommits_info_208_ldest;
        input  io_diffCommits_info_208_pdest;
        input  io_diffCommits_info_208_rfWen;
        input  io_diffCommits_info_208_fpWen;
        input  io_diffCommits_info_208_vecWen;
        input  io_diffCommits_info_208_v0Wen;
        input  io_diffCommits_info_208_vlWen;
        input  io_diffCommits_info_209_ldest;
        input  io_diffCommits_info_209_pdest;
        input  io_diffCommits_info_209_rfWen;
        input  io_diffCommits_info_209_fpWen;
        input  io_diffCommits_info_209_vecWen;
        input  io_diffCommits_info_209_v0Wen;
        input  io_diffCommits_info_209_vlWen;
        input  io_diffCommits_info_210_ldest;
        input  io_diffCommits_info_210_pdest;
        input  io_diffCommits_info_210_rfWen;
        input  io_diffCommits_info_210_fpWen;
        input  io_diffCommits_info_210_vecWen;
        input  io_diffCommits_info_210_v0Wen;
        input  io_diffCommits_info_210_vlWen;
        input  io_diffCommits_info_211_ldest;
        input  io_diffCommits_info_211_pdest;
        input  io_diffCommits_info_211_rfWen;
        input  io_diffCommits_info_211_fpWen;
        input  io_diffCommits_info_211_vecWen;
        input  io_diffCommits_info_211_v0Wen;
        input  io_diffCommits_info_211_vlWen;
        input  io_diffCommits_info_212_ldest;
        input  io_diffCommits_info_212_pdest;
        input  io_diffCommits_info_212_rfWen;
        input  io_diffCommits_info_212_fpWen;
        input  io_diffCommits_info_212_vecWen;
        input  io_diffCommits_info_212_v0Wen;
        input  io_diffCommits_info_212_vlWen;
        input  io_diffCommits_info_213_ldest;
        input  io_diffCommits_info_213_pdest;
        input  io_diffCommits_info_213_rfWen;
        input  io_diffCommits_info_213_fpWen;
        input  io_diffCommits_info_213_vecWen;
        input  io_diffCommits_info_213_v0Wen;
        input  io_diffCommits_info_213_vlWen;
        input  io_diffCommits_info_214_ldest;
        input  io_diffCommits_info_214_pdest;
        input  io_diffCommits_info_214_rfWen;
        input  io_diffCommits_info_214_fpWen;
        input  io_diffCommits_info_214_vecWen;
        input  io_diffCommits_info_214_v0Wen;
        input  io_diffCommits_info_214_vlWen;
        input  io_diffCommits_info_215_ldest;
        input  io_diffCommits_info_215_pdest;
        input  io_diffCommits_info_215_rfWen;
        input  io_diffCommits_info_215_fpWen;
        input  io_diffCommits_info_215_vecWen;
        input  io_diffCommits_info_215_v0Wen;
        input  io_diffCommits_info_215_vlWen;
        input  io_diffCommits_info_216_ldest;
        input  io_diffCommits_info_216_pdest;
        input  io_diffCommits_info_216_rfWen;
        input  io_diffCommits_info_216_fpWen;
        input  io_diffCommits_info_216_vecWen;
        input  io_diffCommits_info_216_v0Wen;
        input  io_diffCommits_info_216_vlWen;
        input  io_diffCommits_info_217_ldest;
        input  io_diffCommits_info_217_pdest;
        input  io_diffCommits_info_217_rfWen;
        input  io_diffCommits_info_217_fpWen;
        input  io_diffCommits_info_217_vecWen;
        input  io_diffCommits_info_217_v0Wen;
        input  io_diffCommits_info_217_vlWen;
        input  io_diffCommits_info_218_ldest;
        input  io_diffCommits_info_218_pdest;
        input  io_diffCommits_info_218_rfWen;
        input  io_diffCommits_info_218_fpWen;
        input  io_diffCommits_info_218_vecWen;
        input  io_diffCommits_info_218_v0Wen;
        input  io_diffCommits_info_218_vlWen;
        input  io_diffCommits_info_219_ldest;
        input  io_diffCommits_info_219_pdest;
        input  io_diffCommits_info_219_rfWen;
        input  io_diffCommits_info_219_fpWen;
        input  io_diffCommits_info_219_vecWen;
        input  io_diffCommits_info_219_v0Wen;
        input  io_diffCommits_info_219_vlWen;
        input  io_diffCommits_info_220_ldest;
        input  io_diffCommits_info_220_pdest;
        input  io_diffCommits_info_220_rfWen;
        input  io_diffCommits_info_220_fpWen;
        input  io_diffCommits_info_220_vecWen;
        input  io_diffCommits_info_220_v0Wen;
        input  io_diffCommits_info_220_vlWen;
        input  io_diffCommits_info_221_ldest;
        input  io_diffCommits_info_221_pdest;
        input  io_diffCommits_info_221_rfWen;
        input  io_diffCommits_info_221_fpWen;
        input  io_diffCommits_info_221_vecWen;
        input  io_diffCommits_info_221_v0Wen;
        input  io_diffCommits_info_221_vlWen;
        input  io_diffCommits_info_222_ldest;
        input  io_diffCommits_info_222_pdest;
        input  io_diffCommits_info_222_rfWen;
        input  io_diffCommits_info_222_fpWen;
        input  io_diffCommits_info_222_vecWen;
        input  io_diffCommits_info_222_v0Wen;
        input  io_diffCommits_info_222_vlWen;
        input  io_diffCommits_info_223_ldest;
        input  io_diffCommits_info_223_pdest;
        input  io_diffCommits_info_223_rfWen;
        input  io_diffCommits_info_223_fpWen;
        input  io_diffCommits_info_223_vecWen;
        input  io_diffCommits_info_223_v0Wen;
        input  io_diffCommits_info_223_vlWen;
        input  io_diffCommits_info_224_ldest;
        input  io_diffCommits_info_224_pdest;
        input  io_diffCommits_info_224_rfWen;
        input  io_diffCommits_info_224_fpWen;
        input  io_diffCommits_info_224_vecWen;
        input  io_diffCommits_info_224_v0Wen;
        input  io_diffCommits_info_224_vlWen;
        input  io_diffCommits_info_225_ldest;
        input  io_diffCommits_info_225_pdest;
        input  io_diffCommits_info_225_rfWen;
        input  io_diffCommits_info_225_fpWen;
        input  io_diffCommits_info_225_vecWen;
        input  io_diffCommits_info_225_v0Wen;
        input  io_diffCommits_info_225_vlWen;
        input  io_diffCommits_info_226_ldest;
        input  io_diffCommits_info_226_pdest;
        input  io_diffCommits_info_226_rfWen;
        input  io_diffCommits_info_226_fpWen;
        input  io_diffCommits_info_226_vecWen;
        input  io_diffCommits_info_226_v0Wen;
        input  io_diffCommits_info_226_vlWen;
        input  io_diffCommits_info_227_ldest;
        input  io_diffCommits_info_227_pdest;
        input  io_diffCommits_info_227_rfWen;
        input  io_diffCommits_info_227_fpWen;
        input  io_diffCommits_info_227_vecWen;
        input  io_diffCommits_info_227_v0Wen;
        input  io_diffCommits_info_227_vlWen;
        input  io_diffCommits_info_228_ldest;
        input  io_diffCommits_info_228_pdest;
        input  io_diffCommits_info_228_rfWen;
        input  io_diffCommits_info_228_fpWen;
        input  io_diffCommits_info_228_vecWen;
        input  io_diffCommits_info_228_v0Wen;
        input  io_diffCommits_info_228_vlWen;
        input  io_diffCommits_info_229_ldest;
        input  io_diffCommits_info_229_pdest;
        input  io_diffCommits_info_229_rfWen;
        input  io_diffCommits_info_229_fpWen;
        input  io_diffCommits_info_229_vecWen;
        input  io_diffCommits_info_229_v0Wen;
        input  io_diffCommits_info_229_vlWen;
        input  io_diffCommits_info_230_ldest;
        input  io_diffCommits_info_230_pdest;
        input  io_diffCommits_info_230_rfWen;
        input  io_diffCommits_info_230_fpWen;
        input  io_diffCommits_info_230_vecWen;
        input  io_diffCommits_info_230_v0Wen;
        input  io_diffCommits_info_230_vlWen;
        input  io_diffCommits_info_231_ldest;
        input  io_diffCommits_info_231_pdest;
        input  io_diffCommits_info_231_rfWen;
        input  io_diffCommits_info_231_fpWen;
        input  io_diffCommits_info_231_vecWen;
        input  io_diffCommits_info_231_v0Wen;
        input  io_diffCommits_info_231_vlWen;
        input  io_diffCommits_info_232_ldest;
        input  io_diffCommits_info_232_pdest;
        input  io_diffCommits_info_232_rfWen;
        input  io_diffCommits_info_232_fpWen;
        input  io_diffCommits_info_232_vecWen;
        input  io_diffCommits_info_232_v0Wen;
        input  io_diffCommits_info_232_vlWen;
        input  io_diffCommits_info_233_ldest;
        input  io_diffCommits_info_233_pdest;
        input  io_diffCommits_info_233_rfWen;
        input  io_diffCommits_info_233_fpWen;
        input  io_diffCommits_info_233_vecWen;
        input  io_diffCommits_info_233_v0Wen;
        input  io_diffCommits_info_233_vlWen;
        input  io_diffCommits_info_234_ldest;
        input  io_diffCommits_info_234_pdest;
        input  io_diffCommits_info_234_rfWen;
        input  io_diffCommits_info_234_fpWen;
        input  io_diffCommits_info_234_vecWen;
        input  io_diffCommits_info_234_v0Wen;
        input  io_diffCommits_info_234_vlWen;
        input  io_diffCommits_info_235_ldest;
        input  io_diffCommits_info_235_pdest;
        input  io_diffCommits_info_235_rfWen;
        input  io_diffCommits_info_235_fpWen;
        input  io_diffCommits_info_235_vecWen;
        input  io_diffCommits_info_235_v0Wen;
        input  io_diffCommits_info_235_vlWen;
        input  io_diffCommits_info_236_ldest;
        input  io_diffCommits_info_236_pdest;
        input  io_diffCommits_info_236_rfWen;
        input  io_diffCommits_info_236_fpWen;
        input  io_diffCommits_info_236_vecWen;
        input  io_diffCommits_info_236_v0Wen;
        input  io_diffCommits_info_236_vlWen;
        input  io_diffCommits_info_237_ldest;
        input  io_diffCommits_info_237_pdest;
        input  io_diffCommits_info_237_rfWen;
        input  io_diffCommits_info_237_fpWen;
        input  io_diffCommits_info_237_vecWen;
        input  io_diffCommits_info_237_v0Wen;
        input  io_diffCommits_info_237_vlWen;
        input  io_diffCommits_info_238_ldest;
        input  io_diffCommits_info_238_pdest;
        input  io_diffCommits_info_238_rfWen;
        input  io_diffCommits_info_238_fpWen;
        input  io_diffCommits_info_238_vecWen;
        input  io_diffCommits_info_238_v0Wen;
        input  io_diffCommits_info_238_vlWen;
        input  io_diffCommits_info_239_ldest;
        input  io_diffCommits_info_239_pdest;
        input  io_diffCommits_info_239_rfWen;
        input  io_diffCommits_info_239_fpWen;
        input  io_diffCommits_info_239_vecWen;
        input  io_diffCommits_info_239_v0Wen;
        input  io_diffCommits_info_239_vlWen;
        input  io_diffCommits_info_240_ldest;
        input  io_diffCommits_info_240_pdest;
        input  io_diffCommits_info_240_rfWen;
        input  io_diffCommits_info_240_fpWen;
        input  io_diffCommits_info_240_vecWen;
        input  io_diffCommits_info_240_v0Wen;
        input  io_diffCommits_info_240_vlWen;
        input  io_diffCommits_info_241_ldest;
        input  io_diffCommits_info_241_pdest;
        input  io_diffCommits_info_241_rfWen;
        input  io_diffCommits_info_241_fpWen;
        input  io_diffCommits_info_241_vecWen;
        input  io_diffCommits_info_241_v0Wen;
        input  io_diffCommits_info_241_vlWen;
        input  io_diffCommits_info_242_ldest;
        input  io_diffCommits_info_242_pdest;
        input  io_diffCommits_info_242_rfWen;
        input  io_diffCommits_info_242_fpWen;
        input  io_diffCommits_info_242_vecWen;
        input  io_diffCommits_info_242_v0Wen;
        input  io_diffCommits_info_242_vlWen;
        input  io_diffCommits_info_243_ldest;
        input  io_diffCommits_info_243_pdest;
        input  io_diffCommits_info_243_rfWen;
        input  io_diffCommits_info_243_fpWen;
        input  io_diffCommits_info_243_vecWen;
        input  io_diffCommits_info_243_v0Wen;
        input  io_diffCommits_info_243_vlWen;
        input  io_diffCommits_info_244_ldest;
        input  io_diffCommits_info_244_pdest;
        input  io_diffCommits_info_244_rfWen;
        input  io_diffCommits_info_244_fpWen;
        input  io_diffCommits_info_244_vecWen;
        input  io_diffCommits_info_244_v0Wen;
        input  io_diffCommits_info_244_vlWen;
        input  io_diffCommits_info_245_ldest;
        input  io_diffCommits_info_245_pdest;
        input  io_diffCommits_info_245_rfWen;
        input  io_diffCommits_info_245_fpWen;
        input  io_diffCommits_info_245_vecWen;
        input  io_diffCommits_info_245_v0Wen;
        input  io_diffCommits_info_245_vlWen;
        input  io_diffCommits_info_246_ldest;
        input  io_diffCommits_info_246_pdest;
        input  io_diffCommits_info_246_rfWen;
        input  io_diffCommits_info_246_fpWen;
        input  io_diffCommits_info_246_vecWen;
        input  io_diffCommits_info_246_v0Wen;
        input  io_diffCommits_info_246_vlWen;
        input  io_diffCommits_info_247_ldest;
        input  io_diffCommits_info_247_pdest;
        input  io_diffCommits_info_247_rfWen;
        input  io_diffCommits_info_247_fpWen;
        input  io_diffCommits_info_247_vecWen;
        input  io_diffCommits_info_247_v0Wen;
        input  io_diffCommits_info_247_vlWen;
        input  io_diffCommits_info_248_ldest;
        input  io_diffCommits_info_248_pdest;
        input  io_diffCommits_info_248_rfWen;
        input  io_diffCommits_info_248_fpWen;
        input  io_diffCommits_info_248_vecWen;
        input  io_diffCommits_info_248_v0Wen;
        input  io_diffCommits_info_248_vlWen;
        input  io_diffCommits_info_249_ldest;
        input  io_diffCommits_info_249_pdest;
        input  io_diffCommits_info_249_rfWen;
        input  io_diffCommits_info_249_fpWen;
        input  io_diffCommits_info_249_vecWen;
        input  io_diffCommits_info_249_v0Wen;
        input  io_diffCommits_info_249_vlWen;
        input  io_diffCommits_info_250_ldest;
        input  io_diffCommits_info_250_pdest;
        input  io_diffCommits_info_250_rfWen;
        input  io_diffCommits_info_250_fpWen;
        input  io_diffCommits_info_250_vecWen;
        input  io_diffCommits_info_250_v0Wen;
        input  io_diffCommits_info_250_vlWen;
        input  io_diffCommits_info_251_ldest;
        input  io_diffCommits_info_251_pdest;
        input  io_diffCommits_info_251_rfWen;
        input  io_diffCommits_info_251_fpWen;
        input  io_diffCommits_info_251_vecWen;
        input  io_diffCommits_info_251_v0Wen;
        input  io_diffCommits_info_251_vlWen;
        input  io_diffCommits_info_252_ldest;
        input  io_diffCommits_info_252_pdest;
        input  io_diffCommits_info_252_rfWen;
        input  io_diffCommits_info_252_fpWen;
        input  io_diffCommits_info_252_vecWen;
        input  io_diffCommits_info_252_v0Wen;
        input  io_diffCommits_info_252_vlWen;
        input  io_diffCommits_info_253_ldest;
        input  io_diffCommits_info_253_pdest;
        input  io_diffCommits_info_253_rfWen;
        input  io_diffCommits_info_253_fpWen;
        input  io_diffCommits_info_253_vecWen;
        input  io_diffCommits_info_253_v0Wen;
        input  io_diffCommits_info_253_vlWen;
        input  io_diffCommits_info_254_ldest;
        input  io_diffCommits_info_254_pdest;
        input  io_diffCommits_info_254_rfWen;
        input  io_diffCommits_info_254_fpWen;
        input  io_diffCommits_info_254_vecWen;
        input  io_diffCommits_info_254_v0Wen;
        input  io_diffCommits_info_254_vlWen;
        input  io_diffCommits_info_255_ldest;
        input  io_diffCommits_info_255_pdest;
        input  io_diffCommits_info_256_ldest;
        input  io_diffCommits_info_256_pdest;
        input  io_diffCommits_info_257_ldest;
        input  io_diffCommits_info_257_pdest;
        input  io_diffCommits_info_258_ldest;
        input  io_diffCommits_info_258_pdest;
        input  io_diffCommits_info_259_ldest;
        input  io_diffCommits_info_259_pdest;
        input  io_diffCommits_info_260_ldest;
        input  io_diffCommits_info_260_pdest;
        input  io_diffCommits_info_261_ldest;
        input  io_diffCommits_info_261_pdest;
        input  io_diffCommits_info_262_ldest;
        input  io_diffCommits_info_262_pdest;
        input  io_diffCommits_info_263_ldest;
        input  io_diffCommits_info_263_pdest;
        input  io_diffCommits_info_264_ldest;
        input  io_diffCommits_info_264_pdest;
        input  io_diffCommits_info_265_ldest;
        input  io_diffCommits_info_265_pdest;
        input  io_diffCommits_info_266_ldest;
        input  io_diffCommits_info_266_pdest;
        input  io_diffCommits_info_267_ldest;
        input  io_diffCommits_info_267_pdest;
        input  io_diffCommits_info_268_ldest;
        input  io_diffCommits_info_268_pdest;
        input  io_diffCommits_info_269_ldest;
        input  io_diffCommits_info_269_pdest;
        input  io_diffCommits_info_270_ldest;
        input  io_diffCommits_info_270_pdest;
        input  io_diffCommits_info_271_ldest;
        input  io_diffCommits_info_271_pdest;
        input  io_diffCommits_info_272_ldest;
        input  io_diffCommits_info_272_pdest;
        input  io_diffCommits_info_273_ldest;
        input  io_diffCommits_info_273_pdest;
        input  io_diffCommits_info_274_ldest;
        input  io_diffCommits_info_274_pdest;
        input  io_diffCommits_info_275_ldest;
        input  io_diffCommits_info_275_pdest;
        input  io_diffCommits_info_276_ldest;
        input  io_diffCommits_info_276_pdest;
        input  io_diffCommits_info_277_ldest;
        input  io_diffCommits_info_277_pdest;
        input  io_diffCommits_info_278_ldest;
        input  io_diffCommits_info_278_pdest;
        input  io_diffCommits_info_279_ldest;
        input  io_diffCommits_info_279_pdest;
        input  io_diffCommits_info_280_ldest;
        input  io_diffCommits_info_280_pdest;
        input  io_diffCommits_info_281_ldest;
        input  io_diffCommits_info_281_pdest;
        input  io_diffCommits_info_282_ldest;
        input  io_diffCommits_info_282_pdest;
        input  io_diffCommits_info_283_ldest;
        input  io_diffCommits_info_283_pdest;
        input  io_diffCommits_info_284_ldest;
        input  io_diffCommits_info_284_pdest;
        input  io_diffCommits_info_285_ldest;
        input  io_diffCommits_info_285_pdest;
        input  io_diffCommits_info_286_ldest;
        input  io_diffCommits_info_286_pdest;
        input  io_diffCommits_info_287_ldest;
        input  io_diffCommits_info_287_pdest;
        input  io_diffCommits_info_288_ldest;
        input  io_diffCommits_info_288_pdest;
        input  io_diffCommits_info_289_ldest;
        input  io_diffCommits_info_289_pdest;
        input  io_diffCommits_info_290_ldest;
        input  io_diffCommits_info_290_pdest;
        input  io_diffCommits_info_291_ldest;
        input  io_diffCommits_info_291_pdest;
        input  io_diffCommits_info_292_ldest;
        input  io_diffCommits_info_292_pdest;
        input  io_diffCommits_info_293_ldest;
        input  io_diffCommits_info_293_pdest;
        input  io_diffCommits_info_294_ldest;
        input  io_diffCommits_info_294_pdest;
        input  io_diffCommits_info_295_ldest;
        input  io_diffCommits_info_295_pdest;
        input  io_diffCommits_info_296_ldest;
        input  io_diffCommits_info_296_pdest;
        input  io_diffCommits_info_297_ldest;
        input  io_diffCommits_info_297_pdest;
        input  io_diffCommits_info_298_ldest;
        input  io_diffCommits_info_298_pdest;
        input  io_diffCommits_info_299_ldest;
        input  io_diffCommits_info_299_pdest;
        input  io_diffCommits_info_300_ldest;
        input  io_diffCommits_info_300_pdest;
        input  io_diffCommits_info_301_ldest;
        input  io_diffCommits_info_301_pdest;
        input  io_diffCommits_info_302_ldest;
        input  io_diffCommits_info_302_pdest;
        input  io_diffCommits_info_303_ldest;
        input  io_diffCommits_info_303_pdest;
        input  io_diffCommits_info_304_ldest;
        input  io_diffCommits_info_304_pdest;
        input  io_diffCommits_info_305_ldest;
        input  io_diffCommits_info_305_pdest;
        input  io_diffCommits_info_306_ldest;
        input  io_diffCommits_info_306_pdest;
        input  io_diffCommits_info_307_ldest;
        input  io_diffCommits_info_307_pdest;
        input  io_diffCommits_info_308_ldest;
        input  io_diffCommits_info_308_pdest;
        input  io_diffCommits_info_309_ldest;
        input  io_diffCommits_info_309_pdest;
        input  io_diffCommits_info_310_ldest;
        input  io_diffCommits_info_310_pdest;
        input  io_diffCommits_info_311_ldest;
        input  io_diffCommits_info_311_pdest;
        input  io_diffCommits_info_312_ldest;
        input  io_diffCommits_info_312_pdest;
        input  io_diffCommits_info_313_ldest;
        input  io_diffCommits_info_313_pdest;
        input  io_diffCommits_info_314_ldest;
        input  io_diffCommits_info_314_pdest;
        input  io_diffCommits_info_315_ldest;
        input  io_diffCommits_info_315_pdest;
        input  io_diffCommits_info_316_ldest;
        input  io_diffCommits_info_316_pdest;
        input  io_diffCommits_info_317_ldest;
        input  io_diffCommits_info_317_pdest;
        input  io_diffCommits_info_318_ldest;
        input  io_diffCommits_info_318_pdest;
        input  io_diffCommits_info_319_ldest;
        input  io_diffCommits_info_319_pdest;
        input  io_diffCommits_info_320_ldest;
        input  io_diffCommits_info_320_pdest;
        input  io_diffCommits_info_321_ldest;
        input  io_diffCommits_info_321_pdest;
        input  io_diffCommits_info_322_ldest;
        input  io_diffCommits_info_322_pdest;
        input  io_diffCommits_info_323_ldest;
        input  io_diffCommits_info_323_pdest;
        input  io_diffCommits_info_324_ldest;
        input  io_diffCommits_info_324_pdest;
        input  io_diffCommits_info_325_ldest;
        input  io_diffCommits_info_325_pdest;
        input  io_diffCommits_info_326_ldest;
        input  io_diffCommits_info_326_pdest;
        input  io_diffCommits_info_327_ldest;
        input  io_diffCommits_info_327_pdest;
        input  io_diffCommits_info_328_ldest;
        input  io_diffCommits_info_328_pdest;
        input  io_diffCommits_info_329_ldest;
        input  io_diffCommits_info_329_pdest;
        input  io_diffCommits_info_330_ldest;
        input  io_diffCommits_info_330_pdest;
        input  io_diffCommits_info_331_ldest;
        input  io_diffCommits_info_331_pdest;
        input  io_diffCommits_info_332_ldest;
        input  io_diffCommits_info_332_pdest;
        input  io_diffCommits_info_333_ldest;
        input  io_diffCommits_info_333_pdest;
        input  io_diffCommits_info_334_ldest;
        input  io_diffCommits_info_334_pdest;
        input  io_diffCommits_info_335_ldest;
        input  io_diffCommits_info_335_pdest;
        input  io_diffCommits_info_336_ldest;
        input  io_diffCommits_info_336_pdest;
        input  io_diffCommits_info_337_ldest;
        input  io_diffCommits_info_337_pdest;
        input  io_diffCommits_info_338_ldest;
        input  io_diffCommits_info_338_pdest;
        input  io_diffCommits_info_339_ldest;
        input  io_diffCommits_info_339_pdest;
        input  io_diffCommits_info_340_ldest;
        input  io_diffCommits_info_340_pdest;
        input  io_diffCommits_info_341_ldest;
        input  io_diffCommits_info_341_pdest;
        input  io_diffCommits_info_342_ldest;
        input  io_diffCommits_info_342_pdest;
        input  io_diffCommits_info_343_ldest;
        input  io_diffCommits_info_343_pdest;
        input  io_diffCommits_info_344_ldest;
        input  io_diffCommits_info_344_pdest;
        input  io_diffCommits_info_345_ldest;
        input  io_diffCommits_info_345_pdest;
        input  io_diffCommits_info_346_ldest;
        input  io_diffCommits_info_346_pdest;
        input  io_diffCommits_info_347_ldest;
        input  io_diffCommits_info_347_pdest;
        input  io_diffCommits_info_348_ldest;
        input  io_diffCommits_info_348_pdest;
        input  io_diffCommits_info_349_ldest;
        input  io_diffCommits_info_349_pdest;
        input  io_diffCommits_info_350_ldest;
        input  io_diffCommits_info_350_pdest;
        input  io_diffCommits_info_351_ldest;
        input  io_diffCommits_info_351_pdest;
        input  io_diffCommits_info_352_ldest;
        input  io_diffCommits_info_352_pdest;
        input  io_diffCommits_info_353_ldest;
        input  io_diffCommits_info_353_pdest;
        input  io_diffCommits_info_354_ldest;
        input  io_diffCommits_info_354_pdest;
        input  io_diffCommits_info_355_ldest;
        input  io_diffCommits_info_355_pdest;
        input  io_diffCommits_info_356_ldest;
        input  io_diffCommits_info_356_pdest;
        input  io_diffCommits_info_357_ldest;
        input  io_diffCommits_info_357_pdest;
        input  io_diffCommits_info_358_ldest;
        input  io_diffCommits_info_358_pdest;
        input  io_diffCommits_info_359_ldest;
        input  io_diffCommits_info_359_pdest;
        input  io_diffCommits_info_360_ldest;
        input  io_diffCommits_info_360_pdest;
        input  io_diffCommits_info_361_ldest;
        input  io_diffCommits_info_361_pdest;
        input  io_diffCommits_info_362_ldest;
        input  io_diffCommits_info_362_pdest;
        input  io_diffCommits_info_363_ldest;
        input  io_diffCommits_info_363_pdest;
        input  io_diffCommits_info_364_ldest;
        input  io_diffCommits_info_364_pdest;
        input  io_diffCommits_info_365_ldest;
        input  io_diffCommits_info_365_pdest;
        input  io_diffCommits_info_366_ldest;
        input  io_diffCommits_info_366_pdest;
        input  io_diffCommits_info_367_ldest;
        input  io_diffCommits_info_367_pdest;
        input  io_diffCommits_info_368_ldest;
        input  io_diffCommits_info_368_pdest;
        input  io_diffCommits_info_369_ldest;
        input  io_diffCommits_info_369_pdest;
        input  io_diffCommits_info_370_ldest;
        input  io_diffCommits_info_370_pdest;
        input  io_diffCommits_info_371_ldest;
        input  io_diffCommits_info_371_pdest;
        input  io_diffCommits_info_372_ldest;
        input  io_diffCommits_info_372_pdest;
        input  io_diffCommits_info_373_ldest;
        input  io_diffCommits_info_373_pdest;
        input  io_diffCommits_info_374_ldest;
        input  io_diffCommits_info_374_pdest;
        input  io_diffCommits_info_375_ldest;
        input  io_diffCommits_info_375_pdest;
        input  io_diffCommits_info_376_ldest;
        input  io_diffCommits_info_376_pdest;
        input  io_diffCommits_info_377_ldest;
        input  io_diffCommits_info_377_pdest;
        input  io_diffCommits_info_378_ldest;
        input  io_diffCommits_info_378_pdest;
        input  io_diffCommits_info_379_ldest;
        input  io_diffCommits_info_379_pdest;
        input  io_diffCommits_info_380_ldest;
        input  io_diffCommits_info_380_pdest;
        input  io_diffCommits_info_381_ldest;
        input  io_diffCommits_info_381_pdest;
        input  io_diffCommits_info_382_ldest;
        input  io_diffCommits_info_382_pdest;
        input  io_diffCommits_info_383_ldest;
        input  io_diffCommits_info_383_pdest;
        input  io_diffCommits_info_384_ldest;
        input  io_diffCommits_info_384_pdest;
        input  io_diffCommits_info_385_ldest;
        input  io_diffCommits_info_385_pdest;
        input  io_diffCommits_info_386_ldest;
        input  io_diffCommits_info_386_pdest;
        input  io_diffCommits_info_387_ldest;
        input  io_diffCommits_info_387_pdest;
        input  io_diffCommits_info_388_ldest;
        input  io_diffCommits_info_388_pdest;
        input  io_diffCommits_info_389_ldest;
        input  io_diffCommits_info_389_pdest;
        input  io_lsq_scommit;
        input  io_lsq_pendingMMIOld;
        input  io_lsq_pendingst;
        input  io_lsq_pendingPtr_flag;
        input  io_lsq_pendingPtr_value;
        input  io_robDeqPtr_flag;
        input  io_robDeqPtr_value;
        input  io_csr_fflags_valid;
        input  io_csr_fflags_bits;
        input  io_csr_vxsat_valid;
        input  io_csr_vxsat_bits;
        input  io_csr_vstart_valid;
        input  io_csr_vstart_bits;
        input  io_csr_dirty_fs;
        input  io_csr_dirty_vs;
        input  io_csr_perfinfo_retiredInstr;
        input  io_cpu_halt;
        input  io_wfi_wfiReq;
        input  io_toDecode_isResumeVType;
        input  io_toDecode_walkToArchVType;
        input  io_toDecode_walkVType_valid;
        input  io_toDecode_walkVType_bits_illegal;
        input  io_toDecode_walkVType_bits_vma;
        input  io_toDecode_walkVType_bits_vta;
        input  io_toDecode_walkVType_bits_vsew;
        input  io_toDecode_walkVType_bits_vlmul;
        input  io_toDecode_commitVType_vtype_valid;
        input  io_toDecode_commitVType_vtype_bits_illegal;
        input  io_toDecode_commitVType_vtype_bits_vma;
        input  io_toDecode_commitVType_vtype_bits_vta;
        input  io_toDecode_commitVType_vtype_bits_vsew;
        input  io_toDecode_commitVType_vtype_bits_vlmul;
        input  io_toDecode_commitVType_hasVsetvl;
        input  io_readGPAMemAddr_valid;
        input  io_readGPAMemAddr_bits_ftqPtr_value;
        input  io_readGPAMemAddr_bits_ftqOffset;
        input  io_toVecExcpMod_logicPhyRegMap_0_valid;
        input  io_toVecExcpMod_logicPhyRegMap_0_bits_lreg;
        input  io_toVecExcpMod_logicPhyRegMap_0_bits_preg;
        input  io_toVecExcpMod_logicPhyRegMap_1_valid;
        input  io_toVecExcpMod_logicPhyRegMap_1_bits_lreg;
        input  io_toVecExcpMod_logicPhyRegMap_1_bits_preg;
        input  io_toVecExcpMod_logicPhyRegMap_2_valid;
        input  io_toVecExcpMod_logicPhyRegMap_2_bits_lreg;
        input  io_toVecExcpMod_logicPhyRegMap_2_bits_preg;
        input  io_toVecExcpMod_logicPhyRegMap_3_valid;
        input  io_toVecExcpMod_logicPhyRegMap_3_bits_lreg;
        input  io_toVecExcpMod_logicPhyRegMap_3_bits_preg;
        input  io_toVecExcpMod_logicPhyRegMap_4_valid;
        input  io_toVecExcpMod_logicPhyRegMap_4_bits_lreg;
        input  io_toVecExcpMod_logicPhyRegMap_4_bits_preg;
        input  io_toVecExcpMod_logicPhyRegMap_5_valid;
        input  io_toVecExcpMod_logicPhyRegMap_5_bits_lreg;
        input  io_toVecExcpMod_logicPhyRegMap_5_bits_preg;
        input  io_toVecExcpMod_excpInfo_valid;
        input  io_toVecExcpMod_excpInfo_bits_vstart;
        input  io_toVecExcpMod_excpInfo_bits_vsew;
        input  io_toVecExcpMod_excpInfo_bits_veew;
        input  io_toVecExcpMod_excpInfo_bits_vlmul;
        input  io_toVecExcpMod_excpInfo_bits_nf;
        input  io_toVecExcpMod_excpInfo_bits_isStride;
        input  io_toVecExcpMod_excpInfo_bits_isIndexed;
        input  io_toVecExcpMod_excpInfo_bits_isWhole;
        input  io_toVecExcpMod_excpInfo_bits_isVlm;
        input  io_storeDebugInfo_1_pc;
        input  io_perf_0_value;
        input  io_perf_1_value;
        input  io_perf_2_value;
        input  io_perf_3_value;
        input  io_perf_4_value;
        input  io_perf_5_value;
        input  io_perf_6_value;
        input  io_perf_7_value;
        input  io_perf_8_value;
        input  io_perf_9_value;
        input  io_perf_10_value;
        input  io_perf_11_value;
        input  io_perf_12_value;
        input  io_perf_13_value;
        input  io_perf_14_value;
        input  io_perf_15_value;
        input  io_perf_16_value;
        input  io_perf_17_value;
        input  io_error_0;

    endclocking:mon_cb

    modport drv_mp (clocking drv_cb);
    modport mon_mp (clocking mon_cb);

endinterface:Rob_output_agent_interface

`endif


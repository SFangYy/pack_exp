//=========================================================
//File name    : WriteBack_in_connect.sv
//Author       : nanyunhao
//Module name  : WriteBack_in_connect
//Discribution : WriteBack_in_connect : WriteBack_in Interface connection macro
//Date         : 2026-01-22
//=========================================================
`ifndef WRITEBACK_IN_CONNECT__SV
`define WRITEBACK_IN_CONNECT__SV

`define ROB__WRITEBACK_IN_CONNECT(U_IF_NAME,AGENT_PATH,RTL_PATH) \
    WriteBack_in_agent_interface  U_IF_NAME (clk,tc_if.rst_n); \
    initial begin \
        uvm_config_db#(virtual WriteBack_in_agent_interface)::set(null,`"*AGENT_PATH*`", "vif", U_IF_NAME); \
    end \
    `ifdef ROB_UT \
    initial begin \
        force RTL_PATH.io_writeback_24_valid = U_IF_NAME.io_writeback_24_valid; \
        force RTL_PATH.io_writeback_24_bits_data_0 = U_IF_NAME.io_writeback_24_bits_data_0; \
        force RTL_PATH.io_writeback_24_bits_pdest = U_IF_NAME.io_writeback_24_bits_pdest; \
        force RTL_PATH.io_writeback_24_bits_robIdx_flag = U_IF_NAME.io_writeback_24_bits_robIdx_flag; \
        force RTL_PATH.io_writeback_24_bits_robIdx_value = U_IF_NAME.io_writeback_24_bits_robIdx_value; \
        force RTL_PATH.io_writeback_24_bits_vecWen = U_IF_NAME.io_writeback_24_bits_vecWen; \
        force RTL_PATH.io_writeback_24_bits_v0Wen = U_IF_NAME.io_writeback_24_bits_v0Wen; \
        force RTL_PATH.io_writeback_24_bits_vlWen = U_IF_NAME.io_writeback_24_bits_vlWen; \
        force RTL_PATH.io_writeback_24_bits_exceptionVec_0 = U_IF_NAME.io_writeback_24_bits_exceptionVec_0; \
        force RTL_PATH.io_writeback_24_bits_exceptionVec_1 = U_IF_NAME.io_writeback_24_bits_exceptionVec_1; \
        force RTL_PATH.io_writeback_24_bits_exceptionVec_2 = U_IF_NAME.io_writeback_24_bits_exceptionVec_2; \
        force RTL_PATH.io_writeback_24_bits_exceptionVec_3 = U_IF_NAME.io_writeback_24_bits_exceptionVec_3; \
        force RTL_PATH.io_writeback_24_bits_exceptionVec_4 = U_IF_NAME.io_writeback_24_bits_exceptionVec_4; \
        force RTL_PATH.io_writeback_24_bits_exceptionVec_5 = U_IF_NAME.io_writeback_24_bits_exceptionVec_5; \
        force RTL_PATH.io_writeback_24_bits_exceptionVec_6 = U_IF_NAME.io_writeback_24_bits_exceptionVec_6; \
        force RTL_PATH.io_writeback_24_bits_exceptionVec_7 = U_IF_NAME.io_writeback_24_bits_exceptionVec_7; \
        force RTL_PATH.io_writeback_24_bits_exceptionVec_8 = U_IF_NAME.io_writeback_24_bits_exceptionVec_8; \
        force RTL_PATH.io_writeback_24_bits_exceptionVec_9 = U_IF_NAME.io_writeback_24_bits_exceptionVec_9; \
        force RTL_PATH.io_writeback_24_bits_exceptionVec_10 = U_IF_NAME.io_writeback_24_bits_exceptionVec_10; \
        force RTL_PATH.io_writeback_24_bits_exceptionVec_11 = U_IF_NAME.io_writeback_24_bits_exceptionVec_11; \
        force RTL_PATH.io_writeback_24_bits_exceptionVec_12 = U_IF_NAME.io_writeback_24_bits_exceptionVec_12; \
        force RTL_PATH.io_writeback_24_bits_exceptionVec_13 = U_IF_NAME.io_writeback_24_bits_exceptionVec_13; \
        force RTL_PATH.io_writeback_24_bits_exceptionVec_14 = U_IF_NAME.io_writeback_24_bits_exceptionVec_14; \
        force RTL_PATH.io_writeback_24_bits_exceptionVec_15 = U_IF_NAME.io_writeback_24_bits_exceptionVec_15; \
        force RTL_PATH.io_writeback_24_bits_exceptionVec_16 = U_IF_NAME.io_writeback_24_bits_exceptionVec_16; \
        force RTL_PATH.io_writeback_24_bits_exceptionVec_17 = U_IF_NAME.io_writeback_24_bits_exceptionVec_17; \
        force RTL_PATH.io_writeback_24_bits_exceptionVec_18 = U_IF_NAME.io_writeback_24_bits_exceptionVec_18; \
        force RTL_PATH.io_writeback_24_bits_exceptionVec_19 = U_IF_NAME.io_writeback_24_bits_exceptionVec_19; \
        force RTL_PATH.io_writeback_24_bits_exceptionVec_20 = U_IF_NAME.io_writeback_24_bits_exceptionVec_20; \
        force RTL_PATH.io_writeback_24_bits_exceptionVec_21 = U_IF_NAME.io_writeback_24_bits_exceptionVec_21; \
        force RTL_PATH.io_writeback_24_bits_exceptionVec_22 = U_IF_NAME.io_writeback_24_bits_exceptionVec_22; \
        force RTL_PATH.io_writeback_24_bits_exceptionVec_23 = U_IF_NAME.io_writeback_24_bits_exceptionVec_23; \
        force RTL_PATH.io_writeback_24_bits_flushPipe = U_IF_NAME.io_writeback_24_bits_flushPipe; \
        force RTL_PATH.io_writeback_24_bits_replay = U_IF_NAME.io_writeback_24_bits_replay; \
        force RTL_PATH.io_writeback_24_bits_trigger = U_IF_NAME.io_writeback_24_bits_trigger; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_vill = U_IF_NAME.io_writeback_24_bits_vls_vpu_vill; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_vma = U_IF_NAME.io_writeback_24_bits_vls_vpu_vma; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_vta = U_IF_NAME.io_writeback_24_bits_vls_vpu_vta; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_vsew = U_IF_NAME.io_writeback_24_bits_vls_vpu_vsew; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_vlmul = U_IF_NAME.io_writeback_24_bits_vls_vpu_vlmul; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_specVill = U_IF_NAME.io_writeback_24_bits_vls_vpu_specVill; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_specVma = U_IF_NAME.io_writeback_24_bits_vls_vpu_specVma; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_specVta = U_IF_NAME.io_writeback_24_bits_vls_vpu_specVta; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_specVsew = U_IF_NAME.io_writeback_24_bits_vls_vpu_specVsew; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_specVlmul = U_IF_NAME.io_writeback_24_bits_vls_vpu_specVlmul; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_vm = U_IF_NAME.io_writeback_24_bits_vls_vpu_vm; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_vstart = U_IF_NAME.io_writeback_24_bits_vls_vpu_vstart; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_frm = U_IF_NAME.io_writeback_24_bits_vls_vpu_frm; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst = U_IF_NAME.io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_fpu_isFP32Instr = U_IF_NAME.io_writeback_24_bits_vls_vpu_fpu_isFP32Instr; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_fpu_isFP64Instr = U_IF_NAME.io_writeback_24_bits_vls_vpu_fpu_isFP64Instr; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_fpu_isReduction = U_IF_NAME.io_writeback_24_bits_vls_vpu_fpu_isReduction; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2 = U_IF_NAME.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4 = U_IF_NAME.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8 = U_IF_NAME.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_vxrm = U_IF_NAME.io_writeback_24_bits_vls_vpu_vxrm; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_vuopIdx = U_IF_NAME.io_writeback_24_bits_vls_vpu_vuopIdx; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_lastUop = U_IF_NAME.io_writeback_24_bits_vls_vpu_lastUop; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_vmask = U_IF_NAME.io_writeback_24_bits_vls_vpu_vmask; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_vl = U_IF_NAME.io_writeback_24_bits_vls_vpu_vl; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_nf = U_IF_NAME.io_writeback_24_bits_vls_vpu_nf; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_veew = U_IF_NAME.io_writeback_24_bits_vls_vpu_veew; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_isReverse = U_IF_NAME.io_writeback_24_bits_vls_vpu_isReverse; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_isExt = U_IF_NAME.io_writeback_24_bits_vls_vpu_isExt; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_isNarrow = U_IF_NAME.io_writeback_24_bits_vls_vpu_isNarrow; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_isDstMask = U_IF_NAME.io_writeback_24_bits_vls_vpu_isDstMask; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_isOpMask = U_IF_NAME.io_writeback_24_bits_vls_vpu_isOpMask; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_isMove = U_IF_NAME.io_writeback_24_bits_vls_vpu_isMove; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_isDependOldVd = U_IF_NAME.io_writeback_24_bits_vls_vpu_isDependOldVd; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_isWritePartVd = U_IF_NAME.io_writeback_24_bits_vls_vpu_isWritePartVd; \
        force RTL_PATH.io_writeback_24_bits_vls_vpu_isVleff = U_IF_NAME.io_writeback_24_bits_vls_vpu_isVleff; \
        force RTL_PATH.io_writeback_24_bits_vls_oldVdPsrc = U_IF_NAME.io_writeback_24_bits_vls_oldVdPsrc; \
        force RTL_PATH.io_writeback_24_bits_vls_vdIdx = U_IF_NAME.io_writeback_24_bits_vls_vdIdx; \
        force RTL_PATH.io_writeback_24_bits_vls_vdIdxInField = U_IF_NAME.io_writeback_24_bits_vls_vdIdxInField; \
        force RTL_PATH.io_writeback_24_bits_vls_isIndexed = U_IF_NAME.io_writeback_24_bits_vls_isIndexed; \
        force RTL_PATH.io_writeback_24_bits_vls_isMasked = U_IF_NAME.io_writeback_24_bits_vls_isMasked; \
        force RTL_PATH.io_writeback_24_bits_vls_isStrided = U_IF_NAME.io_writeback_24_bits_vls_isStrided; \
        force RTL_PATH.io_writeback_24_bits_vls_isWhole = U_IF_NAME.io_writeback_24_bits_vls_isWhole; \
        force RTL_PATH.io_writeback_24_bits_vls_isVecLoad = U_IF_NAME.io_writeback_24_bits_vls_isVecLoad; \
        force RTL_PATH.io_writeback_24_bits_vls_isVlm = U_IF_NAME.io_writeback_24_bits_vls_isVlm; \
        force RTL_PATH.io_writeback_24_bits_debug_isMMIO = U_IF_NAME.io_writeback_24_bits_debug_isMMIO; \
        force RTL_PATH.io_writeback_24_bits_debug_isNCIO = U_IF_NAME.io_writeback_24_bits_debug_isNCIO; \
        force RTL_PATH.io_writeback_24_bits_debug_isPerfCnt = U_IF_NAME.io_writeback_24_bits_debug_isPerfCnt; \
        force RTL_PATH.io_writeback_24_bits_debug_paddr = U_IF_NAME.io_writeback_24_bits_debug_paddr; \
        force RTL_PATH.io_writeback_24_bits_debug_vaddr = U_IF_NAME.io_writeback_24_bits_debug_vaddr; \
        force RTL_PATH.io_writeback_24_bits_debugInfo_eliminatedMove = U_IF_NAME.io_writeback_24_bits_debugInfo_eliminatedMove; \
        force RTL_PATH.io_writeback_24_bits_debugInfo_renameTime = U_IF_NAME.io_writeback_24_bits_debugInfo_renameTime; \
        force RTL_PATH.io_writeback_24_bits_debugInfo_dispatchTime = U_IF_NAME.io_writeback_24_bits_debugInfo_dispatchTime; \
        force RTL_PATH.io_writeback_24_bits_debugInfo_enqRsTime = U_IF_NAME.io_writeback_24_bits_debugInfo_enqRsTime; \
        force RTL_PATH.io_writeback_24_bits_debugInfo_selectTime = U_IF_NAME.io_writeback_24_bits_debugInfo_selectTime; \
        force RTL_PATH.io_writeback_24_bits_debugInfo_issueTime = U_IF_NAME.io_writeback_24_bits_debugInfo_issueTime; \
        force RTL_PATH.io_writeback_24_bits_debugInfo_writebackTime = U_IF_NAME.io_writeback_24_bits_debugInfo_writebackTime; \
        force RTL_PATH.io_writeback_24_bits_debugInfo_runahead_checkpoint_id = U_IF_NAME.io_writeback_24_bits_debugInfo_runahead_checkpoint_id; \
        force RTL_PATH.io_writeback_24_bits_debugInfo_tlbFirstReqTime = U_IF_NAME.io_writeback_24_bits_debugInfo_tlbFirstReqTime; \
        force RTL_PATH.io_writeback_24_bits_debugInfo_tlbRespTime = U_IF_NAME.io_writeback_24_bits_debugInfo_tlbRespTime; \
        force RTL_PATH.io_writeback_24_bits_debug_seqNum = U_IF_NAME.io_writeback_24_bits_debug_seqNum; \
        force RTL_PATH.io_writeback_23_valid = U_IF_NAME.io_writeback_23_valid; \
        force RTL_PATH.io_writeback_23_bits_data_0 = U_IF_NAME.io_writeback_23_bits_data_0; \
        force RTL_PATH.io_writeback_23_bits_pdest = U_IF_NAME.io_writeback_23_bits_pdest; \
        force RTL_PATH.io_writeback_23_bits_robIdx_flag = U_IF_NAME.io_writeback_23_bits_robIdx_flag; \
        force RTL_PATH.io_writeback_23_bits_robIdx_value = U_IF_NAME.io_writeback_23_bits_robIdx_value; \
        force RTL_PATH.io_writeback_23_bits_vecWen = U_IF_NAME.io_writeback_23_bits_vecWen; \
        force RTL_PATH.io_writeback_23_bits_v0Wen = U_IF_NAME.io_writeback_23_bits_v0Wen; \
        force RTL_PATH.io_writeback_23_bits_vlWen = U_IF_NAME.io_writeback_23_bits_vlWen; \
        force RTL_PATH.io_writeback_23_bits_exceptionVec_0 = U_IF_NAME.io_writeback_23_bits_exceptionVec_0; \
        force RTL_PATH.io_writeback_23_bits_exceptionVec_1 = U_IF_NAME.io_writeback_23_bits_exceptionVec_1; \
        force RTL_PATH.io_writeback_23_bits_exceptionVec_2 = U_IF_NAME.io_writeback_23_bits_exceptionVec_2; \
        force RTL_PATH.io_writeback_23_bits_exceptionVec_3 = U_IF_NAME.io_writeback_23_bits_exceptionVec_3; \
        force RTL_PATH.io_writeback_23_bits_exceptionVec_4 = U_IF_NAME.io_writeback_23_bits_exceptionVec_4; \
        force RTL_PATH.io_writeback_23_bits_exceptionVec_5 = U_IF_NAME.io_writeback_23_bits_exceptionVec_5; \
        force RTL_PATH.io_writeback_23_bits_exceptionVec_6 = U_IF_NAME.io_writeback_23_bits_exceptionVec_6; \
        force RTL_PATH.io_writeback_23_bits_exceptionVec_7 = U_IF_NAME.io_writeback_23_bits_exceptionVec_7; \
        force RTL_PATH.io_writeback_23_bits_exceptionVec_8 = U_IF_NAME.io_writeback_23_bits_exceptionVec_8; \
        force RTL_PATH.io_writeback_23_bits_exceptionVec_9 = U_IF_NAME.io_writeback_23_bits_exceptionVec_9; \
        force RTL_PATH.io_writeback_23_bits_exceptionVec_10 = U_IF_NAME.io_writeback_23_bits_exceptionVec_10; \
        force RTL_PATH.io_writeback_23_bits_exceptionVec_11 = U_IF_NAME.io_writeback_23_bits_exceptionVec_11; \
        force RTL_PATH.io_writeback_23_bits_exceptionVec_12 = U_IF_NAME.io_writeback_23_bits_exceptionVec_12; \
        force RTL_PATH.io_writeback_23_bits_exceptionVec_13 = U_IF_NAME.io_writeback_23_bits_exceptionVec_13; \
        force RTL_PATH.io_writeback_23_bits_exceptionVec_14 = U_IF_NAME.io_writeback_23_bits_exceptionVec_14; \
        force RTL_PATH.io_writeback_23_bits_exceptionVec_15 = U_IF_NAME.io_writeback_23_bits_exceptionVec_15; \
        force RTL_PATH.io_writeback_23_bits_exceptionVec_16 = U_IF_NAME.io_writeback_23_bits_exceptionVec_16; \
        force RTL_PATH.io_writeback_23_bits_exceptionVec_17 = U_IF_NAME.io_writeback_23_bits_exceptionVec_17; \
        force RTL_PATH.io_writeback_23_bits_exceptionVec_18 = U_IF_NAME.io_writeback_23_bits_exceptionVec_18; \
        force RTL_PATH.io_writeback_23_bits_exceptionVec_19 = U_IF_NAME.io_writeback_23_bits_exceptionVec_19; \
        force RTL_PATH.io_writeback_23_bits_exceptionVec_20 = U_IF_NAME.io_writeback_23_bits_exceptionVec_20; \
        force RTL_PATH.io_writeback_23_bits_exceptionVec_21 = U_IF_NAME.io_writeback_23_bits_exceptionVec_21; \
        force RTL_PATH.io_writeback_23_bits_exceptionVec_22 = U_IF_NAME.io_writeback_23_bits_exceptionVec_22; \
        force RTL_PATH.io_writeback_23_bits_exceptionVec_23 = U_IF_NAME.io_writeback_23_bits_exceptionVec_23; \
        force RTL_PATH.io_writeback_23_bits_flushPipe = U_IF_NAME.io_writeback_23_bits_flushPipe; \
        force RTL_PATH.io_writeback_23_bits_replay = U_IF_NAME.io_writeback_23_bits_replay; \
        force RTL_PATH.io_writeback_23_bits_trigger = U_IF_NAME.io_writeback_23_bits_trigger; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_vill = U_IF_NAME.io_writeback_23_bits_vls_vpu_vill; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_vma = U_IF_NAME.io_writeback_23_bits_vls_vpu_vma; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_vta = U_IF_NAME.io_writeback_23_bits_vls_vpu_vta; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_vsew = U_IF_NAME.io_writeback_23_bits_vls_vpu_vsew; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_vlmul = U_IF_NAME.io_writeback_23_bits_vls_vpu_vlmul; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_specVill = U_IF_NAME.io_writeback_23_bits_vls_vpu_specVill; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_specVma = U_IF_NAME.io_writeback_23_bits_vls_vpu_specVma; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_specVta = U_IF_NAME.io_writeback_23_bits_vls_vpu_specVta; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_specVsew = U_IF_NAME.io_writeback_23_bits_vls_vpu_specVsew; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_specVlmul = U_IF_NAME.io_writeback_23_bits_vls_vpu_specVlmul; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_vm = U_IF_NAME.io_writeback_23_bits_vls_vpu_vm; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_vstart = U_IF_NAME.io_writeback_23_bits_vls_vpu_vstart; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_frm = U_IF_NAME.io_writeback_23_bits_vls_vpu_frm; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst = U_IF_NAME.io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_fpu_isFP32Instr = U_IF_NAME.io_writeback_23_bits_vls_vpu_fpu_isFP32Instr; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_fpu_isFP64Instr = U_IF_NAME.io_writeback_23_bits_vls_vpu_fpu_isFP64Instr; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_fpu_isReduction = U_IF_NAME.io_writeback_23_bits_vls_vpu_fpu_isReduction; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2 = U_IF_NAME.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4 = U_IF_NAME.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8 = U_IF_NAME.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_vxrm = U_IF_NAME.io_writeback_23_bits_vls_vpu_vxrm; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_vuopIdx = U_IF_NAME.io_writeback_23_bits_vls_vpu_vuopIdx; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_lastUop = U_IF_NAME.io_writeback_23_bits_vls_vpu_lastUop; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_vmask = U_IF_NAME.io_writeback_23_bits_vls_vpu_vmask; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_vl = U_IF_NAME.io_writeback_23_bits_vls_vpu_vl; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_nf = U_IF_NAME.io_writeback_23_bits_vls_vpu_nf; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_veew = U_IF_NAME.io_writeback_23_bits_vls_vpu_veew; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_isReverse = U_IF_NAME.io_writeback_23_bits_vls_vpu_isReverse; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_isExt = U_IF_NAME.io_writeback_23_bits_vls_vpu_isExt; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_isNarrow = U_IF_NAME.io_writeback_23_bits_vls_vpu_isNarrow; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_isDstMask = U_IF_NAME.io_writeback_23_bits_vls_vpu_isDstMask; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_isOpMask = U_IF_NAME.io_writeback_23_bits_vls_vpu_isOpMask; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_isMove = U_IF_NAME.io_writeback_23_bits_vls_vpu_isMove; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_isDependOldVd = U_IF_NAME.io_writeback_23_bits_vls_vpu_isDependOldVd; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_isWritePartVd = U_IF_NAME.io_writeback_23_bits_vls_vpu_isWritePartVd; \
        force RTL_PATH.io_writeback_23_bits_vls_vpu_isVleff = U_IF_NAME.io_writeback_23_bits_vls_vpu_isVleff; \
        force RTL_PATH.io_writeback_23_bits_vls_oldVdPsrc = U_IF_NAME.io_writeback_23_bits_vls_oldVdPsrc; \
        force RTL_PATH.io_writeback_23_bits_vls_vdIdx = U_IF_NAME.io_writeback_23_bits_vls_vdIdx; \
        force RTL_PATH.io_writeback_23_bits_vls_vdIdxInField = U_IF_NAME.io_writeback_23_bits_vls_vdIdxInField; \
        force RTL_PATH.io_writeback_23_bits_vls_isIndexed = U_IF_NAME.io_writeback_23_bits_vls_isIndexed; \
        force RTL_PATH.io_writeback_23_bits_vls_isMasked = U_IF_NAME.io_writeback_23_bits_vls_isMasked; \
        force RTL_PATH.io_writeback_23_bits_vls_isStrided = U_IF_NAME.io_writeback_23_bits_vls_isStrided; \
        force RTL_PATH.io_writeback_23_bits_vls_isWhole = U_IF_NAME.io_writeback_23_bits_vls_isWhole; \
        force RTL_PATH.io_writeback_23_bits_vls_isVecLoad = U_IF_NAME.io_writeback_23_bits_vls_isVecLoad; \
        force RTL_PATH.io_writeback_23_bits_vls_isVlm = U_IF_NAME.io_writeback_23_bits_vls_isVlm; \
        force RTL_PATH.io_writeback_23_bits_debug_isMMIO = U_IF_NAME.io_writeback_23_bits_debug_isMMIO; \
        force RTL_PATH.io_writeback_23_bits_debug_isNCIO = U_IF_NAME.io_writeback_23_bits_debug_isNCIO; \
        force RTL_PATH.io_writeback_23_bits_debug_isPerfCnt = U_IF_NAME.io_writeback_23_bits_debug_isPerfCnt; \
        force RTL_PATH.io_writeback_23_bits_debug_paddr = U_IF_NAME.io_writeback_23_bits_debug_paddr; \
        force RTL_PATH.io_writeback_23_bits_debug_vaddr = U_IF_NAME.io_writeback_23_bits_debug_vaddr; \
        force RTL_PATH.io_writeback_23_bits_debugInfo_eliminatedMove = U_IF_NAME.io_writeback_23_bits_debugInfo_eliminatedMove; \
        force RTL_PATH.io_writeback_23_bits_debugInfo_renameTime = U_IF_NAME.io_writeback_23_bits_debugInfo_renameTime; \
        force RTL_PATH.io_writeback_23_bits_debugInfo_dispatchTime = U_IF_NAME.io_writeback_23_bits_debugInfo_dispatchTime; \
        force RTL_PATH.io_writeback_23_bits_debugInfo_enqRsTime = U_IF_NAME.io_writeback_23_bits_debugInfo_enqRsTime; \
        force RTL_PATH.io_writeback_23_bits_debugInfo_selectTime = U_IF_NAME.io_writeback_23_bits_debugInfo_selectTime; \
        force RTL_PATH.io_writeback_23_bits_debugInfo_issueTime = U_IF_NAME.io_writeback_23_bits_debugInfo_issueTime; \
        force RTL_PATH.io_writeback_23_bits_debugInfo_writebackTime = U_IF_NAME.io_writeback_23_bits_debugInfo_writebackTime; \
        force RTL_PATH.io_writeback_23_bits_debugInfo_runahead_checkpoint_id = U_IF_NAME.io_writeback_23_bits_debugInfo_runahead_checkpoint_id; \
        force RTL_PATH.io_writeback_23_bits_debugInfo_tlbFirstReqTime = U_IF_NAME.io_writeback_23_bits_debugInfo_tlbFirstReqTime; \
        force RTL_PATH.io_writeback_23_bits_debugInfo_tlbRespTime = U_IF_NAME.io_writeback_23_bits_debugInfo_tlbRespTime; \
        force RTL_PATH.io_writeback_23_bits_debug_seqNum = U_IF_NAME.io_writeback_23_bits_debug_seqNum; \
        force RTL_PATH.io_writeback_22_valid = U_IF_NAME.io_writeback_22_valid; \
        force RTL_PATH.io_writeback_22_bits_data_0 = U_IF_NAME.io_writeback_22_bits_data_0; \
        force RTL_PATH.io_writeback_22_bits_pdest = U_IF_NAME.io_writeback_22_bits_pdest; \
        force RTL_PATH.io_writeback_22_bits_robIdx_flag = U_IF_NAME.io_writeback_22_bits_robIdx_flag; \
        force RTL_PATH.io_writeback_22_bits_robIdx_value = U_IF_NAME.io_writeback_22_bits_robIdx_value; \
        force RTL_PATH.io_writeback_22_bits_intWen = U_IF_NAME.io_writeback_22_bits_intWen; \
        force RTL_PATH.io_writeback_22_bits_fpWen = U_IF_NAME.io_writeback_22_bits_fpWen; \
        force RTL_PATH.io_writeback_22_bits_exceptionVec_0 = U_IF_NAME.io_writeback_22_bits_exceptionVec_0; \
        force RTL_PATH.io_writeback_22_bits_exceptionVec_1 = U_IF_NAME.io_writeback_22_bits_exceptionVec_1; \
        force RTL_PATH.io_writeback_22_bits_exceptionVec_2 = U_IF_NAME.io_writeback_22_bits_exceptionVec_2; \
        force RTL_PATH.io_writeback_22_bits_exceptionVec_3 = U_IF_NAME.io_writeback_22_bits_exceptionVec_3; \
        force RTL_PATH.io_writeback_22_bits_exceptionVec_4 = U_IF_NAME.io_writeback_22_bits_exceptionVec_4; \
        force RTL_PATH.io_writeback_22_bits_exceptionVec_5 = U_IF_NAME.io_writeback_22_bits_exceptionVec_5; \
        force RTL_PATH.io_writeback_22_bits_exceptionVec_6 = U_IF_NAME.io_writeback_22_bits_exceptionVec_6; \
        force RTL_PATH.io_writeback_22_bits_exceptionVec_7 = U_IF_NAME.io_writeback_22_bits_exceptionVec_7; \
        force RTL_PATH.io_writeback_22_bits_exceptionVec_8 = U_IF_NAME.io_writeback_22_bits_exceptionVec_8; \
        force RTL_PATH.io_writeback_22_bits_exceptionVec_9 = U_IF_NAME.io_writeback_22_bits_exceptionVec_9; \
        force RTL_PATH.io_writeback_22_bits_exceptionVec_10 = U_IF_NAME.io_writeback_22_bits_exceptionVec_10; \
        force RTL_PATH.io_writeback_22_bits_exceptionVec_11 = U_IF_NAME.io_writeback_22_bits_exceptionVec_11; \
        force RTL_PATH.io_writeback_22_bits_exceptionVec_12 = U_IF_NAME.io_writeback_22_bits_exceptionVec_12; \
        force RTL_PATH.io_writeback_22_bits_exceptionVec_13 = U_IF_NAME.io_writeback_22_bits_exceptionVec_13; \
        force RTL_PATH.io_writeback_22_bits_exceptionVec_14 = U_IF_NAME.io_writeback_22_bits_exceptionVec_14; \
        force RTL_PATH.io_writeback_22_bits_exceptionVec_15 = U_IF_NAME.io_writeback_22_bits_exceptionVec_15; \
        force RTL_PATH.io_writeback_22_bits_exceptionVec_16 = U_IF_NAME.io_writeback_22_bits_exceptionVec_16; \
        force RTL_PATH.io_writeback_22_bits_exceptionVec_17 = U_IF_NAME.io_writeback_22_bits_exceptionVec_17; \
        force RTL_PATH.io_writeback_22_bits_exceptionVec_18 = U_IF_NAME.io_writeback_22_bits_exceptionVec_18; \
        force RTL_PATH.io_writeback_22_bits_exceptionVec_19 = U_IF_NAME.io_writeback_22_bits_exceptionVec_19; \
        force RTL_PATH.io_writeback_22_bits_exceptionVec_20 = U_IF_NAME.io_writeback_22_bits_exceptionVec_20; \
        force RTL_PATH.io_writeback_22_bits_exceptionVec_21 = U_IF_NAME.io_writeback_22_bits_exceptionVec_21; \
        force RTL_PATH.io_writeback_22_bits_exceptionVec_22 = U_IF_NAME.io_writeback_22_bits_exceptionVec_22; \
        force RTL_PATH.io_writeback_22_bits_exceptionVec_23 = U_IF_NAME.io_writeback_22_bits_exceptionVec_23; \
        force RTL_PATH.io_writeback_22_bits_flushPipe = U_IF_NAME.io_writeback_22_bits_flushPipe; \
        force RTL_PATH.io_writeback_22_bits_replay = U_IF_NAME.io_writeback_22_bits_replay; \
        force RTL_PATH.io_writeback_22_bits_lqIdx_flag = U_IF_NAME.io_writeback_22_bits_lqIdx_flag; \
        force RTL_PATH.io_writeback_22_bits_lqIdx_value = U_IF_NAME.io_writeback_22_bits_lqIdx_value; \
        force RTL_PATH.io_writeback_22_bits_trigger = U_IF_NAME.io_writeback_22_bits_trigger; \
        force RTL_PATH.io_writeback_22_bits_predecodeInfo_valid = U_IF_NAME.io_writeback_22_bits_predecodeInfo_valid; \
        force RTL_PATH.io_writeback_22_bits_predecodeInfo_isRVC = U_IF_NAME.io_writeback_22_bits_predecodeInfo_isRVC; \
        force RTL_PATH.io_writeback_22_bits_predecodeInfo_brType = U_IF_NAME.io_writeback_22_bits_predecodeInfo_brType; \
        force RTL_PATH.io_writeback_22_bits_predecodeInfo_isCall = U_IF_NAME.io_writeback_22_bits_predecodeInfo_isCall; \
        force RTL_PATH.io_writeback_22_bits_predecodeInfo_isRet = U_IF_NAME.io_writeback_22_bits_predecodeInfo_isRet; \
        force RTL_PATH.io_writeback_22_bits_debug_isMMIO = U_IF_NAME.io_writeback_22_bits_debug_isMMIO; \
        force RTL_PATH.io_writeback_22_bits_debug_isNCIO = U_IF_NAME.io_writeback_22_bits_debug_isNCIO; \
        force RTL_PATH.io_writeback_22_bits_debug_isPerfCnt = U_IF_NAME.io_writeback_22_bits_debug_isPerfCnt; \
        force RTL_PATH.io_writeback_22_bits_debug_paddr = U_IF_NAME.io_writeback_22_bits_debug_paddr; \
        force RTL_PATH.io_writeback_22_bits_debug_vaddr = U_IF_NAME.io_writeback_22_bits_debug_vaddr; \
        force RTL_PATH.io_writeback_22_bits_debugInfo_eliminatedMove = U_IF_NAME.io_writeback_22_bits_debugInfo_eliminatedMove; \
        force RTL_PATH.io_writeback_22_bits_debugInfo_renameTime = U_IF_NAME.io_writeback_22_bits_debugInfo_renameTime; \
        force RTL_PATH.io_writeback_22_bits_debugInfo_dispatchTime = U_IF_NAME.io_writeback_22_bits_debugInfo_dispatchTime; \
        force RTL_PATH.io_writeback_22_bits_debugInfo_enqRsTime = U_IF_NAME.io_writeback_22_bits_debugInfo_enqRsTime; \
        force RTL_PATH.io_writeback_22_bits_debugInfo_selectTime = U_IF_NAME.io_writeback_22_bits_debugInfo_selectTime; \
        force RTL_PATH.io_writeback_22_bits_debugInfo_issueTime = U_IF_NAME.io_writeback_22_bits_debugInfo_issueTime; \
        force RTL_PATH.io_writeback_22_bits_debugInfo_writebackTime = U_IF_NAME.io_writeback_22_bits_debugInfo_writebackTime; \
        force RTL_PATH.io_writeback_22_bits_debugInfo_runahead_checkpoint_id = U_IF_NAME.io_writeback_22_bits_debugInfo_runahead_checkpoint_id; \
        force RTL_PATH.io_writeback_22_bits_debugInfo_tlbFirstReqTime = U_IF_NAME.io_writeback_22_bits_debugInfo_tlbFirstReqTime; \
        force RTL_PATH.io_writeback_22_bits_debugInfo_tlbRespTime = U_IF_NAME.io_writeback_22_bits_debugInfo_tlbRespTime; \
        force RTL_PATH.io_writeback_22_bits_debug_seqNum = U_IF_NAME.io_writeback_22_bits_debug_seqNum; \
        force RTL_PATH.io_writeback_21_valid = U_IF_NAME.io_writeback_21_valid; \
        force RTL_PATH.io_writeback_21_bits_data_0 = U_IF_NAME.io_writeback_21_bits_data_0; \
        force RTL_PATH.io_writeback_21_bits_pdest = U_IF_NAME.io_writeback_21_bits_pdest; \
        force RTL_PATH.io_writeback_21_bits_robIdx_flag = U_IF_NAME.io_writeback_21_bits_robIdx_flag; \
        force RTL_PATH.io_writeback_21_bits_robIdx_value = U_IF_NAME.io_writeback_21_bits_robIdx_value; \
        force RTL_PATH.io_writeback_21_bits_intWen = U_IF_NAME.io_writeback_21_bits_intWen; \
        force RTL_PATH.io_writeback_21_bits_fpWen = U_IF_NAME.io_writeback_21_bits_fpWen; \
        force RTL_PATH.io_writeback_21_bits_exceptionVec_0 = U_IF_NAME.io_writeback_21_bits_exceptionVec_0; \
        force RTL_PATH.io_writeback_21_bits_exceptionVec_1 = U_IF_NAME.io_writeback_21_bits_exceptionVec_1; \
        force RTL_PATH.io_writeback_21_bits_exceptionVec_2 = U_IF_NAME.io_writeback_21_bits_exceptionVec_2; \
        force RTL_PATH.io_writeback_21_bits_exceptionVec_3 = U_IF_NAME.io_writeback_21_bits_exceptionVec_3; \
        force RTL_PATH.io_writeback_21_bits_exceptionVec_4 = U_IF_NAME.io_writeback_21_bits_exceptionVec_4; \
        force RTL_PATH.io_writeback_21_bits_exceptionVec_5 = U_IF_NAME.io_writeback_21_bits_exceptionVec_5; \
        force RTL_PATH.io_writeback_21_bits_exceptionVec_6 = U_IF_NAME.io_writeback_21_bits_exceptionVec_6; \
        force RTL_PATH.io_writeback_21_bits_exceptionVec_7 = U_IF_NAME.io_writeback_21_bits_exceptionVec_7; \
        force RTL_PATH.io_writeback_21_bits_exceptionVec_8 = U_IF_NAME.io_writeback_21_bits_exceptionVec_8; \
        force RTL_PATH.io_writeback_21_bits_exceptionVec_9 = U_IF_NAME.io_writeback_21_bits_exceptionVec_9; \
        force RTL_PATH.io_writeback_21_bits_exceptionVec_10 = U_IF_NAME.io_writeback_21_bits_exceptionVec_10; \
        force RTL_PATH.io_writeback_21_bits_exceptionVec_11 = U_IF_NAME.io_writeback_21_bits_exceptionVec_11; \
        force RTL_PATH.io_writeback_21_bits_exceptionVec_12 = U_IF_NAME.io_writeback_21_bits_exceptionVec_12; \
        force RTL_PATH.io_writeback_21_bits_exceptionVec_13 = U_IF_NAME.io_writeback_21_bits_exceptionVec_13; \
        force RTL_PATH.io_writeback_21_bits_exceptionVec_14 = U_IF_NAME.io_writeback_21_bits_exceptionVec_14; \
        force RTL_PATH.io_writeback_21_bits_exceptionVec_15 = U_IF_NAME.io_writeback_21_bits_exceptionVec_15; \
        force RTL_PATH.io_writeback_21_bits_exceptionVec_16 = U_IF_NAME.io_writeback_21_bits_exceptionVec_16; \
        force RTL_PATH.io_writeback_21_bits_exceptionVec_17 = U_IF_NAME.io_writeback_21_bits_exceptionVec_17; \
        force RTL_PATH.io_writeback_21_bits_exceptionVec_18 = U_IF_NAME.io_writeback_21_bits_exceptionVec_18; \
        force RTL_PATH.io_writeback_21_bits_exceptionVec_19 = U_IF_NAME.io_writeback_21_bits_exceptionVec_19; \
        force RTL_PATH.io_writeback_21_bits_exceptionVec_20 = U_IF_NAME.io_writeback_21_bits_exceptionVec_20; \
        force RTL_PATH.io_writeback_21_bits_exceptionVec_21 = U_IF_NAME.io_writeback_21_bits_exceptionVec_21; \
        force RTL_PATH.io_writeback_21_bits_exceptionVec_22 = U_IF_NAME.io_writeback_21_bits_exceptionVec_22; \
        force RTL_PATH.io_writeback_21_bits_exceptionVec_23 = U_IF_NAME.io_writeback_21_bits_exceptionVec_23; \
        force RTL_PATH.io_writeback_21_bits_flushPipe = U_IF_NAME.io_writeback_21_bits_flushPipe; \
        force RTL_PATH.io_writeback_21_bits_replay = U_IF_NAME.io_writeback_21_bits_replay; \
        force RTL_PATH.io_writeback_21_bits_lqIdx_flag = U_IF_NAME.io_writeback_21_bits_lqIdx_flag; \
        force RTL_PATH.io_writeback_21_bits_lqIdx_value = U_IF_NAME.io_writeback_21_bits_lqIdx_value; \
        force RTL_PATH.io_writeback_21_bits_trigger = U_IF_NAME.io_writeback_21_bits_trigger; \
        force RTL_PATH.io_writeback_21_bits_predecodeInfo_valid = U_IF_NAME.io_writeback_21_bits_predecodeInfo_valid; \
        force RTL_PATH.io_writeback_21_bits_predecodeInfo_isRVC = U_IF_NAME.io_writeback_21_bits_predecodeInfo_isRVC; \
        force RTL_PATH.io_writeback_21_bits_predecodeInfo_brType = U_IF_NAME.io_writeback_21_bits_predecodeInfo_brType; \
        force RTL_PATH.io_writeback_21_bits_predecodeInfo_isCall = U_IF_NAME.io_writeback_21_bits_predecodeInfo_isCall; \
        force RTL_PATH.io_writeback_21_bits_predecodeInfo_isRet = U_IF_NAME.io_writeback_21_bits_predecodeInfo_isRet; \
        force RTL_PATH.io_writeback_21_bits_debug_isMMIO = U_IF_NAME.io_writeback_21_bits_debug_isMMIO; \
        force RTL_PATH.io_writeback_21_bits_debug_isNCIO = U_IF_NAME.io_writeback_21_bits_debug_isNCIO; \
        force RTL_PATH.io_writeback_21_bits_debug_isPerfCnt = U_IF_NAME.io_writeback_21_bits_debug_isPerfCnt; \
        force RTL_PATH.io_writeback_21_bits_debug_paddr = U_IF_NAME.io_writeback_21_bits_debug_paddr; \
        force RTL_PATH.io_writeback_21_bits_debug_vaddr = U_IF_NAME.io_writeback_21_bits_debug_vaddr; \
        force RTL_PATH.io_writeback_21_bits_debugInfo_eliminatedMove = U_IF_NAME.io_writeback_21_bits_debugInfo_eliminatedMove; \
        force RTL_PATH.io_writeback_21_bits_debugInfo_renameTime = U_IF_NAME.io_writeback_21_bits_debugInfo_renameTime; \
        force RTL_PATH.io_writeback_21_bits_debugInfo_dispatchTime = U_IF_NAME.io_writeback_21_bits_debugInfo_dispatchTime; \
        force RTL_PATH.io_writeback_21_bits_debugInfo_enqRsTime = U_IF_NAME.io_writeback_21_bits_debugInfo_enqRsTime; \
        force RTL_PATH.io_writeback_21_bits_debugInfo_selectTime = U_IF_NAME.io_writeback_21_bits_debugInfo_selectTime; \
        force RTL_PATH.io_writeback_21_bits_debugInfo_issueTime = U_IF_NAME.io_writeback_21_bits_debugInfo_issueTime; \
        force RTL_PATH.io_writeback_21_bits_debugInfo_writebackTime = U_IF_NAME.io_writeback_21_bits_debugInfo_writebackTime; \
        force RTL_PATH.io_writeback_21_bits_debugInfo_runahead_checkpoint_id = U_IF_NAME.io_writeback_21_bits_debugInfo_runahead_checkpoint_id; \
        force RTL_PATH.io_writeback_21_bits_debugInfo_tlbFirstReqTime = U_IF_NAME.io_writeback_21_bits_debugInfo_tlbFirstReqTime; \
        force RTL_PATH.io_writeback_21_bits_debugInfo_tlbRespTime = U_IF_NAME.io_writeback_21_bits_debugInfo_tlbRespTime; \
        force RTL_PATH.io_writeback_21_bits_debug_seqNum = U_IF_NAME.io_writeback_21_bits_debug_seqNum; \
        force RTL_PATH.io_writeback_20_valid = U_IF_NAME.io_writeback_20_valid; \
        force RTL_PATH.io_writeback_20_bits_data_0 = U_IF_NAME.io_writeback_20_bits_data_0; \
        force RTL_PATH.io_writeback_20_bits_pdest = U_IF_NAME.io_writeback_20_bits_pdest; \
        force RTL_PATH.io_writeback_20_bits_robIdx_flag = U_IF_NAME.io_writeback_20_bits_robIdx_flag; \
        force RTL_PATH.io_writeback_20_bits_robIdx_value = U_IF_NAME.io_writeback_20_bits_robIdx_value; \
        force RTL_PATH.io_writeback_20_bits_intWen = U_IF_NAME.io_writeback_20_bits_intWen; \
        force RTL_PATH.io_writeback_20_bits_fpWen = U_IF_NAME.io_writeback_20_bits_fpWen; \
        force RTL_PATH.io_writeback_20_bits_exceptionVec_0 = U_IF_NAME.io_writeback_20_bits_exceptionVec_0; \
        force RTL_PATH.io_writeback_20_bits_exceptionVec_1 = U_IF_NAME.io_writeback_20_bits_exceptionVec_1; \
        force RTL_PATH.io_writeback_20_bits_exceptionVec_2 = U_IF_NAME.io_writeback_20_bits_exceptionVec_2; \
        force RTL_PATH.io_writeback_20_bits_exceptionVec_3 = U_IF_NAME.io_writeback_20_bits_exceptionVec_3; \
        force RTL_PATH.io_writeback_20_bits_exceptionVec_4 = U_IF_NAME.io_writeback_20_bits_exceptionVec_4; \
        force RTL_PATH.io_writeback_20_bits_exceptionVec_5 = U_IF_NAME.io_writeback_20_bits_exceptionVec_5; \
        force RTL_PATH.io_writeback_20_bits_exceptionVec_6 = U_IF_NAME.io_writeback_20_bits_exceptionVec_6; \
        force RTL_PATH.io_writeback_20_bits_exceptionVec_7 = U_IF_NAME.io_writeback_20_bits_exceptionVec_7; \
        force RTL_PATH.io_writeback_20_bits_exceptionVec_8 = U_IF_NAME.io_writeback_20_bits_exceptionVec_8; \
        force RTL_PATH.io_writeback_20_bits_exceptionVec_9 = U_IF_NAME.io_writeback_20_bits_exceptionVec_9; \
        force RTL_PATH.io_writeback_20_bits_exceptionVec_10 = U_IF_NAME.io_writeback_20_bits_exceptionVec_10; \
        force RTL_PATH.io_writeback_20_bits_exceptionVec_11 = U_IF_NAME.io_writeback_20_bits_exceptionVec_11; \
        force RTL_PATH.io_writeback_20_bits_exceptionVec_12 = U_IF_NAME.io_writeback_20_bits_exceptionVec_12; \
        force RTL_PATH.io_writeback_20_bits_exceptionVec_13 = U_IF_NAME.io_writeback_20_bits_exceptionVec_13; \
        force RTL_PATH.io_writeback_20_bits_exceptionVec_14 = U_IF_NAME.io_writeback_20_bits_exceptionVec_14; \
        force RTL_PATH.io_writeback_20_bits_exceptionVec_15 = U_IF_NAME.io_writeback_20_bits_exceptionVec_15; \
        force RTL_PATH.io_writeback_20_bits_exceptionVec_16 = U_IF_NAME.io_writeback_20_bits_exceptionVec_16; \
        force RTL_PATH.io_writeback_20_bits_exceptionVec_17 = U_IF_NAME.io_writeback_20_bits_exceptionVec_17; \
        force RTL_PATH.io_writeback_20_bits_exceptionVec_18 = U_IF_NAME.io_writeback_20_bits_exceptionVec_18; \
        force RTL_PATH.io_writeback_20_bits_exceptionVec_19 = U_IF_NAME.io_writeback_20_bits_exceptionVec_19; \
        force RTL_PATH.io_writeback_20_bits_exceptionVec_20 = U_IF_NAME.io_writeback_20_bits_exceptionVec_20; \
        force RTL_PATH.io_writeback_20_bits_exceptionVec_21 = U_IF_NAME.io_writeback_20_bits_exceptionVec_21; \
        force RTL_PATH.io_writeback_20_bits_exceptionVec_22 = U_IF_NAME.io_writeback_20_bits_exceptionVec_22; \
        force RTL_PATH.io_writeback_20_bits_exceptionVec_23 = U_IF_NAME.io_writeback_20_bits_exceptionVec_23; \
        force RTL_PATH.io_writeback_20_bits_flushPipe = U_IF_NAME.io_writeback_20_bits_flushPipe; \
        force RTL_PATH.io_writeback_20_bits_replay = U_IF_NAME.io_writeback_20_bits_replay; \
        force RTL_PATH.io_writeback_20_bits_lqIdx_flag = U_IF_NAME.io_writeback_20_bits_lqIdx_flag; \
        force RTL_PATH.io_writeback_20_bits_lqIdx_value = U_IF_NAME.io_writeback_20_bits_lqIdx_value; \
        force RTL_PATH.io_writeback_20_bits_trigger = U_IF_NAME.io_writeback_20_bits_trigger; \
        force RTL_PATH.io_writeback_20_bits_predecodeInfo_valid = U_IF_NAME.io_writeback_20_bits_predecodeInfo_valid; \
        force RTL_PATH.io_writeback_20_bits_predecodeInfo_isRVC = U_IF_NAME.io_writeback_20_bits_predecodeInfo_isRVC; \
        force RTL_PATH.io_writeback_20_bits_predecodeInfo_brType = U_IF_NAME.io_writeback_20_bits_predecodeInfo_brType; \
        force RTL_PATH.io_writeback_20_bits_predecodeInfo_isCall = U_IF_NAME.io_writeback_20_bits_predecodeInfo_isCall; \
        force RTL_PATH.io_writeback_20_bits_predecodeInfo_isRet = U_IF_NAME.io_writeback_20_bits_predecodeInfo_isRet; \
        force RTL_PATH.io_writeback_20_bits_debug_isMMIO = U_IF_NAME.io_writeback_20_bits_debug_isMMIO; \
        force RTL_PATH.io_writeback_20_bits_debug_isNCIO = U_IF_NAME.io_writeback_20_bits_debug_isNCIO; \
        force RTL_PATH.io_writeback_20_bits_debug_isPerfCnt = U_IF_NAME.io_writeback_20_bits_debug_isPerfCnt; \
        force RTL_PATH.io_writeback_20_bits_debug_paddr = U_IF_NAME.io_writeback_20_bits_debug_paddr; \
        force RTL_PATH.io_writeback_20_bits_debug_vaddr = U_IF_NAME.io_writeback_20_bits_debug_vaddr; \
        force RTL_PATH.io_writeback_20_bits_debugInfo_eliminatedMove = U_IF_NAME.io_writeback_20_bits_debugInfo_eliminatedMove; \
        force RTL_PATH.io_writeback_20_bits_debugInfo_renameTime = U_IF_NAME.io_writeback_20_bits_debugInfo_renameTime; \
        force RTL_PATH.io_writeback_20_bits_debugInfo_dispatchTime = U_IF_NAME.io_writeback_20_bits_debugInfo_dispatchTime; \
        force RTL_PATH.io_writeback_20_bits_debugInfo_enqRsTime = U_IF_NAME.io_writeback_20_bits_debugInfo_enqRsTime; \
        force RTL_PATH.io_writeback_20_bits_debugInfo_selectTime = U_IF_NAME.io_writeback_20_bits_debugInfo_selectTime; \
        force RTL_PATH.io_writeback_20_bits_debugInfo_issueTime = U_IF_NAME.io_writeback_20_bits_debugInfo_issueTime; \
        force RTL_PATH.io_writeback_20_bits_debugInfo_writebackTime = U_IF_NAME.io_writeback_20_bits_debugInfo_writebackTime; \
        force RTL_PATH.io_writeback_20_bits_debugInfo_runahead_checkpoint_id = U_IF_NAME.io_writeback_20_bits_debugInfo_runahead_checkpoint_id; \
        force RTL_PATH.io_writeback_20_bits_debugInfo_tlbFirstReqTime = U_IF_NAME.io_writeback_20_bits_debugInfo_tlbFirstReqTime; \
        force RTL_PATH.io_writeback_20_bits_debugInfo_tlbRespTime = U_IF_NAME.io_writeback_20_bits_debugInfo_tlbRespTime; \
        force RTL_PATH.io_writeback_20_bits_debug_seqNum = U_IF_NAME.io_writeback_20_bits_debug_seqNum; \
        force RTL_PATH.io_writeback_19_valid = U_IF_NAME.io_writeback_19_valid; \
        force RTL_PATH.io_writeback_19_bits_data_0 = U_IF_NAME.io_writeback_19_bits_data_0; \
        force RTL_PATH.io_writeback_19_bits_pdest = U_IF_NAME.io_writeback_19_bits_pdest; \
        force RTL_PATH.io_writeback_19_bits_robIdx_flag = U_IF_NAME.io_writeback_19_bits_robIdx_flag; \
        force RTL_PATH.io_writeback_19_bits_robIdx_value = U_IF_NAME.io_writeback_19_bits_robIdx_value; \
        force RTL_PATH.io_writeback_19_bits_intWen = U_IF_NAME.io_writeback_19_bits_intWen; \
        force RTL_PATH.io_writeback_19_bits_exceptionVec_0 = U_IF_NAME.io_writeback_19_bits_exceptionVec_0; \
        force RTL_PATH.io_writeback_19_bits_exceptionVec_1 = U_IF_NAME.io_writeback_19_bits_exceptionVec_1; \
        force RTL_PATH.io_writeback_19_bits_exceptionVec_2 = U_IF_NAME.io_writeback_19_bits_exceptionVec_2; \
        force RTL_PATH.io_writeback_19_bits_exceptionVec_3 = U_IF_NAME.io_writeback_19_bits_exceptionVec_3; \
        force RTL_PATH.io_writeback_19_bits_exceptionVec_4 = U_IF_NAME.io_writeback_19_bits_exceptionVec_4; \
        force RTL_PATH.io_writeback_19_bits_exceptionVec_5 = U_IF_NAME.io_writeback_19_bits_exceptionVec_5; \
        force RTL_PATH.io_writeback_19_bits_exceptionVec_6 = U_IF_NAME.io_writeback_19_bits_exceptionVec_6; \
        force RTL_PATH.io_writeback_19_bits_exceptionVec_7 = U_IF_NAME.io_writeback_19_bits_exceptionVec_7; \
        force RTL_PATH.io_writeback_19_bits_exceptionVec_8 = U_IF_NAME.io_writeback_19_bits_exceptionVec_8; \
        force RTL_PATH.io_writeback_19_bits_exceptionVec_9 = U_IF_NAME.io_writeback_19_bits_exceptionVec_9; \
        force RTL_PATH.io_writeback_19_bits_exceptionVec_10 = U_IF_NAME.io_writeback_19_bits_exceptionVec_10; \
        force RTL_PATH.io_writeback_19_bits_exceptionVec_11 = U_IF_NAME.io_writeback_19_bits_exceptionVec_11; \
        force RTL_PATH.io_writeback_19_bits_exceptionVec_12 = U_IF_NAME.io_writeback_19_bits_exceptionVec_12; \
        force RTL_PATH.io_writeback_19_bits_exceptionVec_13 = U_IF_NAME.io_writeback_19_bits_exceptionVec_13; \
        force RTL_PATH.io_writeback_19_bits_exceptionVec_14 = U_IF_NAME.io_writeback_19_bits_exceptionVec_14; \
        force RTL_PATH.io_writeback_19_bits_exceptionVec_15 = U_IF_NAME.io_writeback_19_bits_exceptionVec_15; \
        force RTL_PATH.io_writeback_19_bits_exceptionVec_16 = U_IF_NAME.io_writeback_19_bits_exceptionVec_16; \
        force RTL_PATH.io_writeback_19_bits_exceptionVec_17 = U_IF_NAME.io_writeback_19_bits_exceptionVec_17; \
        force RTL_PATH.io_writeback_19_bits_exceptionVec_18 = U_IF_NAME.io_writeback_19_bits_exceptionVec_18; \
        force RTL_PATH.io_writeback_19_bits_exceptionVec_19 = U_IF_NAME.io_writeback_19_bits_exceptionVec_19; \
        force RTL_PATH.io_writeback_19_bits_exceptionVec_20 = U_IF_NAME.io_writeback_19_bits_exceptionVec_20; \
        force RTL_PATH.io_writeback_19_bits_exceptionVec_21 = U_IF_NAME.io_writeback_19_bits_exceptionVec_21; \
        force RTL_PATH.io_writeback_19_bits_exceptionVec_22 = U_IF_NAME.io_writeback_19_bits_exceptionVec_22; \
        force RTL_PATH.io_writeback_19_bits_exceptionVec_23 = U_IF_NAME.io_writeback_19_bits_exceptionVec_23; \
        force RTL_PATH.io_writeback_19_bits_flushPipe = U_IF_NAME.io_writeback_19_bits_flushPipe; \
        force RTL_PATH.io_writeback_19_bits_sqIdx_flag = U_IF_NAME.io_writeback_19_bits_sqIdx_flag; \
        force RTL_PATH.io_writeback_19_bits_sqIdx_value = U_IF_NAME.io_writeback_19_bits_sqIdx_value; \
        force RTL_PATH.io_writeback_19_bits_trigger = U_IF_NAME.io_writeback_19_bits_trigger; \
        force RTL_PATH.io_writeback_19_bits_debug_isMMIO = U_IF_NAME.io_writeback_19_bits_debug_isMMIO; \
        force RTL_PATH.io_writeback_19_bits_debug_isNCIO = U_IF_NAME.io_writeback_19_bits_debug_isNCIO; \
        force RTL_PATH.io_writeback_19_bits_debug_isPerfCnt = U_IF_NAME.io_writeback_19_bits_debug_isPerfCnt; \
        force RTL_PATH.io_writeback_19_bits_debug_paddr = U_IF_NAME.io_writeback_19_bits_debug_paddr; \
        force RTL_PATH.io_writeback_19_bits_debug_vaddr = U_IF_NAME.io_writeback_19_bits_debug_vaddr; \
        force RTL_PATH.io_writeback_19_bits_debugInfo_eliminatedMove = U_IF_NAME.io_writeback_19_bits_debugInfo_eliminatedMove; \
        force RTL_PATH.io_writeback_19_bits_debugInfo_renameTime = U_IF_NAME.io_writeback_19_bits_debugInfo_renameTime; \
        force RTL_PATH.io_writeback_19_bits_debugInfo_dispatchTime = U_IF_NAME.io_writeback_19_bits_debugInfo_dispatchTime; \
        force RTL_PATH.io_writeback_19_bits_debugInfo_enqRsTime = U_IF_NAME.io_writeback_19_bits_debugInfo_enqRsTime; \
        force RTL_PATH.io_writeback_19_bits_debugInfo_selectTime = U_IF_NAME.io_writeback_19_bits_debugInfo_selectTime; \
        force RTL_PATH.io_writeback_19_bits_debugInfo_issueTime = U_IF_NAME.io_writeback_19_bits_debugInfo_issueTime; \
        force RTL_PATH.io_writeback_19_bits_debugInfo_writebackTime = U_IF_NAME.io_writeback_19_bits_debugInfo_writebackTime; \
        force RTL_PATH.io_writeback_19_bits_debugInfo_runahead_checkpoint_id = U_IF_NAME.io_writeback_19_bits_debugInfo_runahead_checkpoint_id; \
        force RTL_PATH.io_writeback_19_bits_debugInfo_tlbFirstReqTime = U_IF_NAME.io_writeback_19_bits_debugInfo_tlbFirstReqTime; \
        force RTL_PATH.io_writeback_19_bits_debugInfo_tlbRespTime = U_IF_NAME.io_writeback_19_bits_debugInfo_tlbRespTime; \
        force RTL_PATH.io_writeback_19_bits_debug_seqNum = U_IF_NAME.io_writeback_19_bits_debug_seqNum; \
        force RTL_PATH.io_writeback_18_valid = U_IF_NAME.io_writeback_18_valid; \
        force RTL_PATH.io_writeback_18_bits_data_0 = U_IF_NAME.io_writeback_18_bits_data_0; \
        force RTL_PATH.io_writeback_18_bits_pdest = U_IF_NAME.io_writeback_18_bits_pdest; \
        force RTL_PATH.io_writeback_18_bits_robIdx_flag = U_IF_NAME.io_writeback_18_bits_robIdx_flag; \
        force RTL_PATH.io_writeback_18_bits_robIdx_value = U_IF_NAME.io_writeback_18_bits_robIdx_value; \
        force RTL_PATH.io_writeback_18_bits_intWen = U_IF_NAME.io_writeback_18_bits_intWen; \
        force RTL_PATH.io_writeback_18_bits_exceptionVec_0 = U_IF_NAME.io_writeback_18_bits_exceptionVec_0; \
        force RTL_PATH.io_writeback_18_bits_exceptionVec_1 = U_IF_NAME.io_writeback_18_bits_exceptionVec_1; \
        force RTL_PATH.io_writeback_18_bits_exceptionVec_2 = U_IF_NAME.io_writeback_18_bits_exceptionVec_2; \
        force RTL_PATH.io_writeback_18_bits_exceptionVec_3 = U_IF_NAME.io_writeback_18_bits_exceptionVec_3; \
        force RTL_PATH.io_writeback_18_bits_exceptionVec_4 = U_IF_NAME.io_writeback_18_bits_exceptionVec_4; \
        force RTL_PATH.io_writeback_18_bits_exceptionVec_5 = U_IF_NAME.io_writeback_18_bits_exceptionVec_5; \
        force RTL_PATH.io_writeback_18_bits_exceptionVec_6 = U_IF_NAME.io_writeback_18_bits_exceptionVec_6; \
        force RTL_PATH.io_writeback_18_bits_exceptionVec_7 = U_IF_NAME.io_writeback_18_bits_exceptionVec_7; \
        force RTL_PATH.io_writeback_18_bits_exceptionVec_8 = U_IF_NAME.io_writeback_18_bits_exceptionVec_8; \
        force RTL_PATH.io_writeback_18_bits_exceptionVec_9 = U_IF_NAME.io_writeback_18_bits_exceptionVec_9; \
        force RTL_PATH.io_writeback_18_bits_exceptionVec_10 = U_IF_NAME.io_writeback_18_bits_exceptionVec_10; \
        force RTL_PATH.io_writeback_18_bits_exceptionVec_11 = U_IF_NAME.io_writeback_18_bits_exceptionVec_11; \
        force RTL_PATH.io_writeback_18_bits_exceptionVec_12 = U_IF_NAME.io_writeback_18_bits_exceptionVec_12; \
        force RTL_PATH.io_writeback_18_bits_exceptionVec_13 = U_IF_NAME.io_writeback_18_bits_exceptionVec_13; \
        force RTL_PATH.io_writeback_18_bits_exceptionVec_14 = U_IF_NAME.io_writeback_18_bits_exceptionVec_14; \
        force RTL_PATH.io_writeback_18_bits_exceptionVec_15 = U_IF_NAME.io_writeback_18_bits_exceptionVec_15; \
        force RTL_PATH.io_writeback_18_bits_exceptionVec_16 = U_IF_NAME.io_writeback_18_bits_exceptionVec_16; \
        force RTL_PATH.io_writeback_18_bits_exceptionVec_17 = U_IF_NAME.io_writeback_18_bits_exceptionVec_17; \
        force RTL_PATH.io_writeback_18_bits_exceptionVec_18 = U_IF_NAME.io_writeback_18_bits_exceptionVec_18; \
        force RTL_PATH.io_writeback_18_bits_exceptionVec_19 = U_IF_NAME.io_writeback_18_bits_exceptionVec_19; \
        force RTL_PATH.io_writeback_18_bits_exceptionVec_20 = U_IF_NAME.io_writeback_18_bits_exceptionVec_20; \
        force RTL_PATH.io_writeback_18_bits_exceptionVec_21 = U_IF_NAME.io_writeback_18_bits_exceptionVec_21; \
        force RTL_PATH.io_writeback_18_bits_exceptionVec_22 = U_IF_NAME.io_writeback_18_bits_exceptionVec_22; \
        force RTL_PATH.io_writeback_18_bits_exceptionVec_23 = U_IF_NAME.io_writeback_18_bits_exceptionVec_23; \
        force RTL_PATH.io_writeback_18_bits_flushPipe = U_IF_NAME.io_writeback_18_bits_flushPipe; \
        force RTL_PATH.io_writeback_18_bits_sqIdx_flag = U_IF_NAME.io_writeback_18_bits_sqIdx_flag; \
        force RTL_PATH.io_writeback_18_bits_sqIdx_value = U_IF_NAME.io_writeback_18_bits_sqIdx_value; \
        force RTL_PATH.io_writeback_18_bits_trigger = U_IF_NAME.io_writeback_18_bits_trigger; \
        force RTL_PATH.io_writeback_18_bits_debug_isMMIO = U_IF_NAME.io_writeback_18_bits_debug_isMMIO; \
        force RTL_PATH.io_writeback_18_bits_debug_isNCIO = U_IF_NAME.io_writeback_18_bits_debug_isNCIO; \
        force RTL_PATH.io_writeback_18_bits_debug_isPerfCnt = U_IF_NAME.io_writeback_18_bits_debug_isPerfCnt; \
        force RTL_PATH.io_writeback_18_bits_debug_paddr = U_IF_NAME.io_writeback_18_bits_debug_paddr; \
        force RTL_PATH.io_writeback_18_bits_debug_vaddr = U_IF_NAME.io_writeback_18_bits_debug_vaddr; \
        force RTL_PATH.io_writeback_18_bits_debugInfo_eliminatedMove = U_IF_NAME.io_writeback_18_bits_debugInfo_eliminatedMove; \
        force RTL_PATH.io_writeback_18_bits_debugInfo_renameTime = U_IF_NAME.io_writeback_18_bits_debugInfo_renameTime; \
        force RTL_PATH.io_writeback_18_bits_debugInfo_dispatchTime = U_IF_NAME.io_writeback_18_bits_debugInfo_dispatchTime; \
        force RTL_PATH.io_writeback_18_bits_debugInfo_enqRsTime = U_IF_NAME.io_writeback_18_bits_debugInfo_enqRsTime; \
        force RTL_PATH.io_writeback_18_bits_debugInfo_selectTime = U_IF_NAME.io_writeback_18_bits_debugInfo_selectTime; \
        force RTL_PATH.io_writeback_18_bits_debugInfo_issueTime = U_IF_NAME.io_writeback_18_bits_debugInfo_issueTime; \
        force RTL_PATH.io_writeback_18_bits_debugInfo_writebackTime = U_IF_NAME.io_writeback_18_bits_debugInfo_writebackTime; \
        force RTL_PATH.io_writeback_18_bits_debugInfo_runahead_checkpoint_id = U_IF_NAME.io_writeback_18_bits_debugInfo_runahead_checkpoint_id; \
        force RTL_PATH.io_writeback_18_bits_debugInfo_tlbFirstReqTime = U_IF_NAME.io_writeback_18_bits_debugInfo_tlbFirstReqTime; \
        force RTL_PATH.io_writeback_18_bits_debugInfo_tlbRespTime = U_IF_NAME.io_writeback_18_bits_debugInfo_tlbRespTime; \
        force RTL_PATH.io_writeback_18_bits_debug_seqNum = U_IF_NAME.io_writeback_18_bits_debug_seqNum; \
        force RTL_PATH.io_writeback_17_valid = U_IF_NAME.io_writeback_17_valid; \
        force RTL_PATH.io_writeback_17_bits_data_0 = U_IF_NAME.io_writeback_17_bits_data_0; \
        force RTL_PATH.io_writeback_17_bits_data_1 = U_IF_NAME.io_writeback_17_bits_data_1; \
        force RTL_PATH.io_writeback_17_bits_data_2 = U_IF_NAME.io_writeback_17_bits_data_2; \
        force RTL_PATH.io_writeback_17_bits_pdest = U_IF_NAME.io_writeback_17_bits_pdest; \
        force RTL_PATH.io_writeback_17_bits_robIdx_flag = U_IF_NAME.io_writeback_17_bits_robIdx_flag; \
        force RTL_PATH.io_writeback_17_bits_robIdx_value = U_IF_NAME.io_writeback_17_bits_robIdx_value; \
        force RTL_PATH.io_writeback_17_bits_vecWen = U_IF_NAME.io_writeback_17_bits_vecWen; \
        force RTL_PATH.io_writeback_17_bits_v0Wen = U_IF_NAME.io_writeback_17_bits_v0Wen; \
        force RTL_PATH.io_writeback_17_bits_fflags = U_IF_NAME.io_writeback_17_bits_fflags; \
        force RTL_PATH.io_writeback_17_bits_wflags = U_IF_NAME.io_writeback_17_bits_wflags; \
        force RTL_PATH.io_writeback_17_bits_debugInfo_eliminatedMove = U_IF_NAME.io_writeback_17_bits_debugInfo_eliminatedMove; \
        force RTL_PATH.io_writeback_17_bits_debugInfo_renameTime = U_IF_NAME.io_writeback_17_bits_debugInfo_renameTime; \
        force RTL_PATH.io_writeback_17_bits_debugInfo_dispatchTime = U_IF_NAME.io_writeback_17_bits_debugInfo_dispatchTime; \
        force RTL_PATH.io_writeback_17_bits_debugInfo_enqRsTime = U_IF_NAME.io_writeback_17_bits_debugInfo_enqRsTime; \
        force RTL_PATH.io_writeback_17_bits_debugInfo_selectTime = U_IF_NAME.io_writeback_17_bits_debugInfo_selectTime; \
        force RTL_PATH.io_writeback_17_bits_debugInfo_issueTime = U_IF_NAME.io_writeback_17_bits_debugInfo_issueTime; \
        force RTL_PATH.io_writeback_17_bits_debugInfo_writebackTime = U_IF_NAME.io_writeback_17_bits_debugInfo_writebackTime; \
        force RTL_PATH.io_writeback_17_bits_debugInfo_runahead_checkpoint_id = U_IF_NAME.io_writeback_17_bits_debugInfo_runahead_checkpoint_id; \
        force RTL_PATH.io_writeback_17_bits_debugInfo_tlbFirstReqTime = U_IF_NAME.io_writeback_17_bits_debugInfo_tlbFirstReqTime; \
        force RTL_PATH.io_writeback_17_bits_debugInfo_tlbRespTime = U_IF_NAME.io_writeback_17_bits_debugInfo_tlbRespTime; \
        force RTL_PATH.io_writeback_17_bits_debug_seqNum = U_IF_NAME.io_writeback_17_bits_debug_seqNum; \
        force RTL_PATH.io_writeback_16_valid = U_IF_NAME.io_writeback_16_valid; \
        force RTL_PATH.io_writeback_16_bits_data_0 = U_IF_NAME.io_writeback_16_bits_data_0; \
        force RTL_PATH.io_writeback_16_bits_data_1 = U_IF_NAME.io_writeback_16_bits_data_1; \
        force RTL_PATH.io_writeback_16_bits_data_2 = U_IF_NAME.io_writeback_16_bits_data_2; \
        force RTL_PATH.io_writeback_16_bits_data_3 = U_IF_NAME.io_writeback_16_bits_data_3; \
        force RTL_PATH.io_writeback_16_bits_pdest = U_IF_NAME.io_writeback_16_bits_pdest; \
        force RTL_PATH.io_writeback_16_bits_robIdx_flag = U_IF_NAME.io_writeback_16_bits_robIdx_flag; \
        force RTL_PATH.io_writeback_16_bits_robIdx_value = U_IF_NAME.io_writeback_16_bits_robIdx_value; \
        force RTL_PATH.io_writeback_16_bits_fpWen = U_IF_NAME.io_writeback_16_bits_fpWen; \
        force RTL_PATH.io_writeback_16_bits_vecWen = U_IF_NAME.io_writeback_16_bits_vecWen; \
        force RTL_PATH.io_writeback_16_bits_v0Wen = U_IF_NAME.io_writeback_16_bits_v0Wen; \
        force RTL_PATH.io_writeback_16_bits_fflags = U_IF_NAME.io_writeback_16_bits_fflags; \
        force RTL_PATH.io_writeback_16_bits_wflags = U_IF_NAME.io_writeback_16_bits_wflags; \
        force RTL_PATH.io_writeback_16_bits_debugInfo_eliminatedMove = U_IF_NAME.io_writeback_16_bits_debugInfo_eliminatedMove; \
        force RTL_PATH.io_writeback_16_bits_debugInfo_renameTime = U_IF_NAME.io_writeback_16_bits_debugInfo_renameTime; \
        force RTL_PATH.io_writeback_16_bits_debugInfo_dispatchTime = U_IF_NAME.io_writeback_16_bits_debugInfo_dispatchTime; \
        force RTL_PATH.io_writeback_16_bits_debugInfo_enqRsTime = U_IF_NAME.io_writeback_16_bits_debugInfo_enqRsTime; \
        force RTL_PATH.io_writeback_16_bits_debugInfo_selectTime = U_IF_NAME.io_writeback_16_bits_debugInfo_selectTime; \
        force RTL_PATH.io_writeback_16_bits_debugInfo_issueTime = U_IF_NAME.io_writeback_16_bits_debugInfo_issueTime; \
        force RTL_PATH.io_writeback_16_bits_debugInfo_writebackTime = U_IF_NAME.io_writeback_16_bits_debugInfo_writebackTime; \
        force RTL_PATH.io_writeback_16_bits_debugInfo_runahead_checkpoint_id = U_IF_NAME.io_writeback_16_bits_debugInfo_runahead_checkpoint_id; \
        force RTL_PATH.io_writeback_16_bits_debugInfo_tlbFirstReqTime = U_IF_NAME.io_writeback_16_bits_debugInfo_tlbFirstReqTime; \
        force RTL_PATH.io_writeback_16_bits_debugInfo_tlbRespTime = U_IF_NAME.io_writeback_16_bits_debugInfo_tlbRespTime; \
        force RTL_PATH.io_writeback_16_bits_debug_seqNum = U_IF_NAME.io_writeback_16_bits_debug_seqNum; \
        force RTL_PATH.io_writeback_15_valid = U_IF_NAME.io_writeback_15_valid; \
        force RTL_PATH.io_writeback_15_bits_data_0 = U_IF_NAME.io_writeback_15_bits_data_0; \
        force RTL_PATH.io_writeback_15_bits_data_1 = U_IF_NAME.io_writeback_15_bits_data_1; \
        force RTL_PATH.io_writeback_15_bits_data_2 = U_IF_NAME.io_writeback_15_bits_data_2; \
        force RTL_PATH.io_writeback_15_bits_pdest = U_IF_NAME.io_writeback_15_bits_pdest; \
        force RTL_PATH.io_writeback_15_bits_robIdx_flag = U_IF_NAME.io_writeback_15_bits_robIdx_flag; \
        force RTL_PATH.io_writeback_15_bits_robIdx_value = U_IF_NAME.io_writeback_15_bits_robIdx_value; \
        force RTL_PATH.io_writeback_15_bits_vecWen = U_IF_NAME.io_writeback_15_bits_vecWen; \
        force RTL_PATH.io_writeback_15_bits_v0Wen = U_IF_NAME.io_writeback_15_bits_v0Wen; \
        force RTL_PATH.io_writeback_15_bits_fflags = U_IF_NAME.io_writeback_15_bits_fflags; \
        force RTL_PATH.io_writeback_15_bits_wflags = U_IF_NAME.io_writeback_15_bits_wflags; \
        force RTL_PATH.io_writeback_15_bits_vxsat = U_IF_NAME.io_writeback_15_bits_vxsat; \
        force RTL_PATH.io_writeback_15_bits_debugInfo_eliminatedMove = U_IF_NAME.io_writeback_15_bits_debugInfo_eliminatedMove; \
        force RTL_PATH.io_writeback_15_bits_debugInfo_renameTime = U_IF_NAME.io_writeback_15_bits_debugInfo_renameTime; \
        force RTL_PATH.io_writeback_15_bits_debugInfo_dispatchTime = U_IF_NAME.io_writeback_15_bits_debugInfo_dispatchTime; \
        force RTL_PATH.io_writeback_15_bits_debugInfo_enqRsTime = U_IF_NAME.io_writeback_15_bits_debugInfo_enqRsTime; \
        force RTL_PATH.io_writeback_15_bits_debugInfo_selectTime = U_IF_NAME.io_writeback_15_bits_debugInfo_selectTime; \
        force RTL_PATH.io_writeback_15_bits_debugInfo_issueTime = U_IF_NAME.io_writeback_15_bits_debugInfo_issueTime; \
        force RTL_PATH.io_writeback_15_bits_debugInfo_writebackTime = U_IF_NAME.io_writeback_15_bits_debugInfo_writebackTime; \
        force RTL_PATH.io_writeback_15_bits_debugInfo_runahead_checkpoint_id = U_IF_NAME.io_writeback_15_bits_debugInfo_runahead_checkpoint_id; \
        force RTL_PATH.io_writeback_15_bits_debugInfo_tlbFirstReqTime = U_IF_NAME.io_writeback_15_bits_debugInfo_tlbFirstReqTime; \
        force RTL_PATH.io_writeback_15_bits_debugInfo_tlbRespTime = U_IF_NAME.io_writeback_15_bits_debugInfo_tlbRespTime; \
        force RTL_PATH.io_writeback_15_bits_debug_seqNum = U_IF_NAME.io_writeback_15_bits_debug_seqNum; \
        force RTL_PATH.io_writeback_14_valid = U_IF_NAME.io_writeback_14_valid; \
        force RTL_PATH.io_writeback_14_bits_data_0 = U_IF_NAME.io_writeback_14_bits_data_0; \
        force RTL_PATH.io_writeback_14_bits_data_1 = U_IF_NAME.io_writeback_14_bits_data_1; \
        force RTL_PATH.io_writeback_14_bits_data_2 = U_IF_NAME.io_writeback_14_bits_data_2; \
        force RTL_PATH.io_writeback_14_bits_data_3 = U_IF_NAME.io_writeback_14_bits_data_3; \
        force RTL_PATH.io_writeback_14_bits_data_4 = U_IF_NAME.io_writeback_14_bits_data_4; \
        force RTL_PATH.io_writeback_14_bits_data_5 = U_IF_NAME.io_writeback_14_bits_data_5; \
        force RTL_PATH.io_writeback_14_bits_pdest = U_IF_NAME.io_writeback_14_bits_pdest; \
        force RTL_PATH.io_writeback_14_bits_robIdx_flag = U_IF_NAME.io_writeback_14_bits_robIdx_flag; \
        force RTL_PATH.io_writeback_14_bits_robIdx_value = U_IF_NAME.io_writeback_14_bits_robIdx_value; \
        force RTL_PATH.io_writeback_14_bits_intWen = U_IF_NAME.io_writeback_14_bits_intWen; \
        force RTL_PATH.io_writeback_14_bits_fpWen = U_IF_NAME.io_writeback_14_bits_fpWen; \
        force RTL_PATH.io_writeback_14_bits_vecWen = U_IF_NAME.io_writeback_14_bits_vecWen; \
        force RTL_PATH.io_writeback_14_bits_v0Wen = U_IF_NAME.io_writeback_14_bits_v0Wen; \
        force RTL_PATH.io_writeback_14_bits_vlWen = U_IF_NAME.io_writeback_14_bits_vlWen; \
        force RTL_PATH.io_writeback_14_bits_fflags = U_IF_NAME.io_writeback_14_bits_fflags; \
        force RTL_PATH.io_writeback_14_bits_wflags = U_IF_NAME.io_writeback_14_bits_wflags; \
        force RTL_PATH.io_writeback_14_bits_exceptionVec_2 = U_IF_NAME.io_writeback_14_bits_exceptionVec_2; \
        force RTL_PATH.io_writeback_14_bits_debugInfo_eliminatedMove = U_IF_NAME.io_writeback_14_bits_debugInfo_eliminatedMove; \
        force RTL_PATH.io_writeback_14_bits_debugInfo_renameTime = U_IF_NAME.io_writeback_14_bits_debugInfo_renameTime; \
        force RTL_PATH.io_writeback_14_bits_debugInfo_dispatchTime = U_IF_NAME.io_writeback_14_bits_debugInfo_dispatchTime; \
        force RTL_PATH.io_writeback_14_bits_debugInfo_enqRsTime = U_IF_NAME.io_writeback_14_bits_debugInfo_enqRsTime; \
        force RTL_PATH.io_writeback_14_bits_debugInfo_selectTime = U_IF_NAME.io_writeback_14_bits_debugInfo_selectTime; \
        force RTL_PATH.io_writeback_14_bits_debugInfo_issueTime = U_IF_NAME.io_writeback_14_bits_debugInfo_issueTime; \
        force RTL_PATH.io_writeback_14_bits_debugInfo_writebackTime = U_IF_NAME.io_writeback_14_bits_debugInfo_writebackTime; \
        force RTL_PATH.io_writeback_14_bits_debugInfo_runahead_checkpoint_id = U_IF_NAME.io_writeback_14_bits_debugInfo_runahead_checkpoint_id; \
        force RTL_PATH.io_writeback_14_bits_debugInfo_tlbFirstReqTime = U_IF_NAME.io_writeback_14_bits_debugInfo_tlbFirstReqTime; \
        force RTL_PATH.io_writeback_14_bits_debugInfo_tlbRespTime = U_IF_NAME.io_writeback_14_bits_debugInfo_tlbRespTime; \
        force RTL_PATH.io_writeback_14_bits_debug_seqNum = U_IF_NAME.io_writeback_14_bits_debug_seqNum; \
        force RTL_PATH.io_writeback_13_valid = U_IF_NAME.io_writeback_13_valid; \
        force RTL_PATH.io_writeback_13_bits_data_0 = U_IF_NAME.io_writeback_13_bits_data_0; \
        force RTL_PATH.io_writeback_13_bits_data_1 = U_IF_NAME.io_writeback_13_bits_data_1; \
        force RTL_PATH.io_writeback_13_bits_data_2 = U_IF_NAME.io_writeback_13_bits_data_2; \
        force RTL_PATH.io_writeback_13_bits_pdest = U_IF_NAME.io_writeback_13_bits_pdest; \
        force RTL_PATH.io_writeback_13_bits_robIdx_flag = U_IF_NAME.io_writeback_13_bits_robIdx_flag; \
        force RTL_PATH.io_writeback_13_bits_robIdx_value = U_IF_NAME.io_writeback_13_bits_robIdx_value; \
        force RTL_PATH.io_writeback_13_bits_vecWen = U_IF_NAME.io_writeback_13_bits_vecWen; \
        force RTL_PATH.io_writeback_13_bits_v0Wen = U_IF_NAME.io_writeback_13_bits_v0Wen; \
        force RTL_PATH.io_writeback_13_bits_fflags = U_IF_NAME.io_writeback_13_bits_fflags; \
        force RTL_PATH.io_writeback_13_bits_wflags = U_IF_NAME.io_writeback_13_bits_wflags; \
        force RTL_PATH.io_writeback_13_bits_vxsat = U_IF_NAME.io_writeback_13_bits_vxsat; \
        force RTL_PATH.io_writeback_13_bits_exceptionVec_2 = U_IF_NAME.io_writeback_13_bits_exceptionVec_2; \
        force RTL_PATH.io_writeback_13_bits_debugInfo_eliminatedMove = U_IF_NAME.io_writeback_13_bits_debugInfo_eliminatedMove; \
        force RTL_PATH.io_writeback_13_bits_debugInfo_renameTime = U_IF_NAME.io_writeback_13_bits_debugInfo_renameTime; \
        force RTL_PATH.io_writeback_13_bits_debugInfo_dispatchTime = U_IF_NAME.io_writeback_13_bits_debugInfo_dispatchTime; \
        force RTL_PATH.io_writeback_13_bits_debugInfo_enqRsTime = U_IF_NAME.io_writeback_13_bits_debugInfo_enqRsTime; \
        force RTL_PATH.io_writeback_13_bits_debugInfo_selectTime = U_IF_NAME.io_writeback_13_bits_debugInfo_selectTime; \
        force RTL_PATH.io_writeback_13_bits_debugInfo_issueTime = U_IF_NAME.io_writeback_13_bits_debugInfo_issueTime; \
        force RTL_PATH.io_writeback_13_bits_debugInfo_writebackTime = U_IF_NAME.io_writeback_13_bits_debugInfo_writebackTime; \
        force RTL_PATH.io_writeback_13_bits_debugInfo_runahead_checkpoint_id = U_IF_NAME.io_writeback_13_bits_debugInfo_runahead_checkpoint_id; \
        force RTL_PATH.io_writeback_13_bits_debugInfo_tlbFirstReqTime = U_IF_NAME.io_writeback_13_bits_debugInfo_tlbFirstReqTime; \
        force RTL_PATH.io_writeback_13_bits_debugInfo_tlbRespTime = U_IF_NAME.io_writeback_13_bits_debugInfo_tlbRespTime; \
        force RTL_PATH.io_writeback_13_bits_debug_seqNum = U_IF_NAME.io_writeback_13_bits_debug_seqNum; \
        force RTL_PATH.io_writeback_7_valid = U_IF_NAME.io_writeback_7_valid; \
        force RTL_PATH.io_writeback_7_bits_data_0 = U_IF_NAME.io_writeback_7_bits_data_0; \
        force RTL_PATH.io_writeback_7_bits_data_1 = U_IF_NAME.io_writeback_7_bits_data_1; \
        force RTL_PATH.io_writeback_7_bits_pdest = U_IF_NAME.io_writeback_7_bits_pdest; \
        force RTL_PATH.io_writeback_7_bits_robIdx_flag = U_IF_NAME.io_writeback_7_bits_robIdx_flag; \
        force RTL_PATH.io_writeback_7_bits_robIdx_value = U_IF_NAME.io_writeback_7_bits_robIdx_value; \
        force RTL_PATH.io_writeback_7_bits_intWen = U_IF_NAME.io_writeback_7_bits_intWen; \
        force RTL_PATH.io_writeback_7_bits_redirect_valid = U_IF_NAME.io_writeback_7_bits_redirect_valid; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_isRVC = U_IF_NAME.io_writeback_7_bits_redirect_bits_isRVC; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_robIdx_flag = U_IF_NAME.io_writeback_7_bits_redirect_bits_robIdx_flag; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_robIdx_value = U_IF_NAME.io_writeback_7_bits_redirect_bits_robIdx_value; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_ftqIdx_flag = U_IF_NAME.io_writeback_7_bits_redirect_bits_ftqIdx_flag; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_ftqIdx_value = U_IF_NAME.io_writeback_7_bits_redirect_bits_ftqIdx_value; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_ftqOffset = U_IF_NAME.io_writeback_7_bits_redirect_bits_ftqOffset; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_level = U_IF_NAME.io_writeback_7_bits_redirect_bits_level; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_interrupt = U_IF_NAME.io_writeback_7_bits_redirect_bits_interrupt; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_pc = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_pc; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_ssp = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_ssp; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_sctr = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_sctr; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0 = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1 = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2 = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3 = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0 = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1 = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2 = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3 = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0 = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1 = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2 = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3 = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0 = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1 = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2 = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3 = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0 = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1 = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2 = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3 = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0 = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1 = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2 = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3 = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_ghr = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_ghr; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0 = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1 = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_target = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_target; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_taken = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_taken; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_shift = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_shift; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF = U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_fullTarget = U_IF_NAME.io_writeback_7_bits_redirect_bits_fullTarget; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_stFtqIdx_flag = U_IF_NAME.io_writeback_7_bits_redirect_bits_stFtqIdx_flag; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_stFtqIdx_value = U_IF_NAME.io_writeback_7_bits_redirect_bits_stFtqIdx_value; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_stFtqOffset = U_IF_NAME.io_writeback_7_bits_redirect_bits_stFtqOffset; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id = U_IF_NAME.io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_debugIsCtrl = U_IF_NAME.io_writeback_7_bits_redirect_bits_debugIsCtrl; \
        force RTL_PATH.io_writeback_7_bits_redirect_bits_debugIsMemVio = U_IF_NAME.io_writeback_7_bits_redirect_bits_debugIsMemVio; \
        force RTL_PATH.io_writeback_7_bits_exceptionVec_2 = U_IF_NAME.io_writeback_7_bits_exceptionVec_2; \
        force RTL_PATH.io_writeback_7_bits_exceptionVec_3 = U_IF_NAME.io_writeback_7_bits_exceptionVec_3; \
        force RTL_PATH.io_writeback_7_bits_exceptionVec_8 = U_IF_NAME.io_writeback_7_bits_exceptionVec_8; \
        force RTL_PATH.io_writeback_7_bits_exceptionVec_9 = U_IF_NAME.io_writeback_7_bits_exceptionVec_9; \
        force RTL_PATH.io_writeback_7_bits_exceptionVec_10 = U_IF_NAME.io_writeback_7_bits_exceptionVec_10; \
        force RTL_PATH.io_writeback_7_bits_exceptionVec_11 = U_IF_NAME.io_writeback_7_bits_exceptionVec_11; \
        force RTL_PATH.io_writeback_7_bits_exceptionVec_22 = U_IF_NAME.io_writeback_7_bits_exceptionVec_22; \
        force RTL_PATH.io_writeback_7_bits_flushPipe = U_IF_NAME.io_writeback_7_bits_flushPipe; \
        force RTL_PATH.io_writeback_7_bits_predecodeInfo_valid = U_IF_NAME.io_writeback_7_bits_predecodeInfo_valid; \
        force RTL_PATH.io_writeback_7_bits_predecodeInfo_isRVC = U_IF_NAME.io_writeback_7_bits_predecodeInfo_isRVC; \
        force RTL_PATH.io_writeback_7_bits_predecodeInfo_brType = U_IF_NAME.io_writeback_7_bits_predecodeInfo_brType; \
        force RTL_PATH.io_writeback_7_bits_predecodeInfo_isCall = U_IF_NAME.io_writeback_7_bits_predecodeInfo_isCall; \
        force RTL_PATH.io_writeback_7_bits_predecodeInfo_isRet = U_IF_NAME.io_writeback_7_bits_predecodeInfo_isRet; \
        force RTL_PATH.io_writeback_7_bits_debug_isPerfCnt = U_IF_NAME.io_writeback_7_bits_debug_isPerfCnt; \
        force RTL_PATH.io_writeback_7_bits_debugInfo_eliminatedMove = U_IF_NAME.io_writeback_7_bits_debugInfo_eliminatedMove; \
        force RTL_PATH.io_writeback_7_bits_debugInfo_renameTime = U_IF_NAME.io_writeback_7_bits_debugInfo_renameTime; \
        force RTL_PATH.io_writeback_7_bits_debugInfo_dispatchTime = U_IF_NAME.io_writeback_7_bits_debugInfo_dispatchTime; \
        force RTL_PATH.io_writeback_7_bits_debugInfo_enqRsTime = U_IF_NAME.io_writeback_7_bits_debugInfo_enqRsTime; \
        force RTL_PATH.io_writeback_7_bits_debugInfo_selectTime = U_IF_NAME.io_writeback_7_bits_debugInfo_selectTime; \
        force RTL_PATH.io_writeback_7_bits_debugInfo_issueTime = U_IF_NAME.io_writeback_7_bits_debugInfo_issueTime; \
        force RTL_PATH.io_writeback_7_bits_debugInfo_writebackTime = U_IF_NAME.io_writeback_7_bits_debugInfo_writebackTime; \
        force RTL_PATH.io_writeback_7_bits_debugInfo_runahead_checkpoint_id = U_IF_NAME.io_writeback_7_bits_debugInfo_runahead_checkpoint_id; \
        force RTL_PATH.io_writeback_7_bits_debugInfo_tlbFirstReqTime = U_IF_NAME.io_writeback_7_bits_debugInfo_tlbFirstReqTime; \
        force RTL_PATH.io_writeback_7_bits_debugInfo_tlbRespTime = U_IF_NAME.io_writeback_7_bits_debugInfo_tlbRespTime; \
        force RTL_PATH.io_writeback_7_bits_debug_seqNum = U_IF_NAME.io_writeback_7_bits_debug_seqNum; \
        force RTL_PATH.io_writeback_5_valid = U_IF_NAME.io_writeback_5_valid; \
        force RTL_PATH.io_writeback_5_bits_redirect_valid = U_IF_NAME.io_writeback_5_bits_redirect_valid; \
        force RTL_PATH.io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred = U_IF_NAME.io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred; \
        force RTL_PATH.io_writeback_3_valid = U_IF_NAME.io_writeback_3_valid; \
        force RTL_PATH.io_writeback_3_bits_redirect_valid = U_IF_NAME.io_writeback_3_bits_redirect_valid; \
        force RTL_PATH.io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred = U_IF_NAME.io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred; \
        force RTL_PATH.io_writeback_1_valid = U_IF_NAME.io_writeback_1_valid; \
        force RTL_PATH.io_writeback_1_bits_redirect_valid = U_IF_NAME.io_writeback_1_bits_redirect_valid; \
        force RTL_PATH.io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred = U_IF_NAME.io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred; \
        force RTL_PATH.io_exuWriteback_26_valid = U_IF_NAME.io_exuWriteback_26_valid; \
        force RTL_PATH.io_exuWriteback_26_bits_robIdx_value = U_IF_NAME.io_exuWriteback_26_bits_robIdx_value; \
        force RTL_PATH.io_exuWriteback_25_valid = U_IF_NAME.io_exuWriteback_25_valid; \
        force RTL_PATH.io_exuWriteback_25_bits_robIdx_value = U_IF_NAME.io_exuWriteback_25_bits_robIdx_value; \
        force RTL_PATH.io_exuWriteback_24_valid = U_IF_NAME.io_exuWriteback_24_valid; \
        force RTL_PATH.io_exuWriteback_24_bits_data_0 = U_IF_NAME.io_exuWriteback_24_bits_data_0; \
        force RTL_PATH.io_exuWriteback_24_bits_pdest = U_IF_NAME.io_exuWriteback_24_bits_pdest; \
        force RTL_PATH.io_exuWriteback_24_bits_robIdx_value = U_IF_NAME.io_exuWriteback_24_bits_robIdx_value; \
        force RTL_PATH.io_exuWriteback_24_bits_vecWen = U_IF_NAME.io_exuWriteback_24_bits_vecWen; \
        force RTL_PATH.io_exuWriteback_24_bits_v0Wen = U_IF_NAME.io_exuWriteback_24_bits_v0Wen; \
        force RTL_PATH.io_exuWriteback_24_bits_vls_vdIdx = U_IF_NAME.io_exuWriteback_24_bits_vls_vdIdx; \
        force RTL_PATH.io_exuWriteback_24_bits_debug_isMMIO = U_IF_NAME.io_exuWriteback_24_bits_debug_isMMIO; \
        force RTL_PATH.io_exuWriteback_24_bits_debug_isNCIO = U_IF_NAME.io_exuWriteback_24_bits_debug_isNCIO; \
        force RTL_PATH.io_exuWriteback_24_bits_debug_isPerfCnt = U_IF_NAME.io_exuWriteback_24_bits_debug_isPerfCnt; \
        force RTL_PATH.io_exuWriteback_24_bits_debug_paddr = U_IF_NAME.io_exuWriteback_24_bits_debug_paddr; \
        force RTL_PATH.io_exuWriteback_23_valid = U_IF_NAME.io_exuWriteback_23_valid; \
        force RTL_PATH.io_exuWriteback_23_bits_data_0 = U_IF_NAME.io_exuWriteback_23_bits_data_0; \
        force RTL_PATH.io_exuWriteback_23_bits_pdest = U_IF_NAME.io_exuWriteback_23_bits_pdest; \
        force RTL_PATH.io_exuWriteback_23_bits_robIdx_value = U_IF_NAME.io_exuWriteback_23_bits_robIdx_value; \
        force RTL_PATH.io_exuWriteback_23_bits_vecWen = U_IF_NAME.io_exuWriteback_23_bits_vecWen; \
        force RTL_PATH.io_exuWriteback_23_bits_v0Wen = U_IF_NAME.io_exuWriteback_23_bits_v0Wen; \
        force RTL_PATH.io_exuWriteback_23_bits_vls_vdIdx = U_IF_NAME.io_exuWriteback_23_bits_vls_vdIdx; \
        force RTL_PATH.io_exuWriteback_23_bits_debug_isMMIO = U_IF_NAME.io_exuWriteback_23_bits_debug_isMMIO; \
        force RTL_PATH.io_exuWriteback_23_bits_debug_isNCIO = U_IF_NAME.io_exuWriteback_23_bits_debug_isNCIO; \
        force RTL_PATH.io_exuWriteback_23_bits_debug_isPerfCnt = U_IF_NAME.io_exuWriteback_23_bits_debug_isPerfCnt; \
        force RTL_PATH.io_exuWriteback_23_bits_debug_paddr = U_IF_NAME.io_exuWriteback_23_bits_debug_paddr; \
        force RTL_PATH.io_exuWriteback_22_valid = U_IF_NAME.io_exuWriteback_22_valid; \
        force RTL_PATH.io_exuWriteback_22_bits_data_0 = U_IF_NAME.io_exuWriteback_22_bits_data_0; \
        force RTL_PATH.io_exuWriteback_22_bits_robIdx_value = U_IF_NAME.io_exuWriteback_22_bits_robIdx_value; \
        force RTL_PATH.io_exuWriteback_22_bits_lqIdx_value = U_IF_NAME.io_exuWriteback_22_bits_lqIdx_value; \
        force RTL_PATH.io_exuWriteback_22_bits_debug_isMMIO = U_IF_NAME.io_exuWriteback_22_bits_debug_isMMIO; \
        force RTL_PATH.io_exuWriteback_22_bits_debug_isNCIO = U_IF_NAME.io_exuWriteback_22_bits_debug_isNCIO; \
        force RTL_PATH.io_exuWriteback_22_bits_debug_isPerfCnt = U_IF_NAME.io_exuWriteback_22_bits_debug_isPerfCnt; \
        force RTL_PATH.io_exuWriteback_22_bits_debug_paddr = U_IF_NAME.io_exuWriteback_22_bits_debug_paddr; \
        force RTL_PATH.io_exuWriteback_21_valid = U_IF_NAME.io_exuWriteback_21_valid; \
        force RTL_PATH.io_exuWriteback_21_bits_data_0 = U_IF_NAME.io_exuWriteback_21_bits_data_0; \
        force RTL_PATH.io_exuWriteback_21_bits_robIdx_value = U_IF_NAME.io_exuWriteback_21_bits_robIdx_value; \
        force RTL_PATH.io_exuWriteback_21_bits_lqIdx_value = U_IF_NAME.io_exuWriteback_21_bits_lqIdx_value; \
        force RTL_PATH.io_exuWriteback_21_bits_debug_isMMIO = U_IF_NAME.io_exuWriteback_21_bits_debug_isMMIO; \
        force RTL_PATH.io_exuWriteback_21_bits_debug_isNCIO = U_IF_NAME.io_exuWriteback_21_bits_debug_isNCIO; \
        force RTL_PATH.io_exuWriteback_21_bits_debug_isPerfCnt = U_IF_NAME.io_exuWriteback_21_bits_debug_isPerfCnt; \
        force RTL_PATH.io_exuWriteback_21_bits_debug_paddr = U_IF_NAME.io_exuWriteback_21_bits_debug_paddr; \
        force RTL_PATH.io_exuWriteback_20_valid = U_IF_NAME.io_exuWriteback_20_valid; \
        force RTL_PATH.io_exuWriteback_20_bits_data_0 = U_IF_NAME.io_exuWriteback_20_bits_data_0; \
        force RTL_PATH.io_exuWriteback_20_bits_robIdx_value = U_IF_NAME.io_exuWriteback_20_bits_robIdx_value; \
        force RTL_PATH.io_exuWriteback_20_bits_lqIdx_value = U_IF_NAME.io_exuWriteback_20_bits_lqIdx_value; \
        force RTL_PATH.io_exuWriteback_20_bits_debug_isMMIO = U_IF_NAME.io_exuWriteback_20_bits_debug_isMMIO; \
        force RTL_PATH.io_exuWriteback_20_bits_debug_isNCIO = U_IF_NAME.io_exuWriteback_20_bits_debug_isNCIO; \
        force RTL_PATH.io_exuWriteback_20_bits_debug_isPerfCnt = U_IF_NAME.io_exuWriteback_20_bits_debug_isPerfCnt; \
        force RTL_PATH.io_exuWriteback_20_bits_debug_paddr = U_IF_NAME.io_exuWriteback_20_bits_debug_paddr; \
        force RTL_PATH.io_exuWriteback_19_valid = U_IF_NAME.io_exuWriteback_19_valid; \
        force RTL_PATH.io_exuWriteback_19_bits_data_0 = U_IF_NAME.io_exuWriteback_19_bits_data_0; \
        force RTL_PATH.io_exuWriteback_19_bits_robIdx_value = U_IF_NAME.io_exuWriteback_19_bits_robIdx_value; \
        force RTL_PATH.io_exuWriteback_19_bits_sqIdx_value = U_IF_NAME.io_exuWriteback_19_bits_sqIdx_value; \
        force RTL_PATH.io_exuWriteback_19_bits_debug_isMMIO = U_IF_NAME.io_exuWriteback_19_bits_debug_isMMIO; \
        force RTL_PATH.io_exuWriteback_19_bits_debug_isNCIO = U_IF_NAME.io_exuWriteback_19_bits_debug_isNCIO; \
        force RTL_PATH.io_exuWriteback_19_bits_debug_isPerfCnt = U_IF_NAME.io_exuWriteback_19_bits_debug_isPerfCnt; \
        force RTL_PATH.io_exuWriteback_19_bits_debug_paddr = U_IF_NAME.io_exuWriteback_19_bits_debug_paddr; \
        force RTL_PATH.io_exuWriteback_18_valid = U_IF_NAME.io_exuWriteback_18_valid; \
        force RTL_PATH.io_exuWriteback_18_bits_data_0 = U_IF_NAME.io_exuWriteback_18_bits_data_0; \
        force RTL_PATH.io_exuWriteback_18_bits_robIdx_value = U_IF_NAME.io_exuWriteback_18_bits_robIdx_value; \
        force RTL_PATH.io_exuWriteback_18_bits_sqIdx_value = U_IF_NAME.io_exuWriteback_18_bits_sqIdx_value; \
        force RTL_PATH.io_exuWriteback_18_bits_debug_isMMIO = U_IF_NAME.io_exuWriteback_18_bits_debug_isMMIO; \
        force RTL_PATH.io_exuWriteback_18_bits_debug_isNCIO = U_IF_NAME.io_exuWriteback_18_bits_debug_isNCIO; \
        force RTL_PATH.io_exuWriteback_18_bits_debug_isPerfCnt = U_IF_NAME.io_exuWriteback_18_bits_debug_isPerfCnt; \
        force RTL_PATH.io_exuWriteback_18_bits_debug_paddr = U_IF_NAME.io_exuWriteback_18_bits_debug_paddr; \
        force RTL_PATH.io_exuWriteback_17_valid = U_IF_NAME.io_exuWriteback_17_valid; \
        force RTL_PATH.io_exuWriteback_17_bits_data_0 = U_IF_NAME.io_exuWriteback_17_bits_data_0; \
        force RTL_PATH.io_exuWriteback_17_bits_robIdx_value = U_IF_NAME.io_exuWriteback_17_bits_robIdx_value; \
        force RTL_PATH.io_exuWriteback_17_bits_fflags = U_IF_NAME.io_exuWriteback_17_bits_fflags; \
        force RTL_PATH.io_exuWriteback_17_bits_wflags = U_IF_NAME.io_exuWriteback_17_bits_wflags; \
        force RTL_PATH.io_exuWriteback_16_valid = U_IF_NAME.io_exuWriteback_16_valid; \
        force RTL_PATH.io_exuWriteback_16_bits_data_0 = U_IF_NAME.io_exuWriteback_16_bits_data_0; \
        force RTL_PATH.io_exuWriteback_16_bits_robIdx_value = U_IF_NAME.io_exuWriteback_16_bits_robIdx_value; \
        force RTL_PATH.io_exuWriteback_16_bits_fflags = U_IF_NAME.io_exuWriteback_16_bits_fflags; \
        force RTL_PATH.io_exuWriteback_16_bits_wflags = U_IF_NAME.io_exuWriteback_16_bits_wflags; \
        force RTL_PATH.io_exuWriteback_15_valid = U_IF_NAME.io_exuWriteback_15_valid; \
        force RTL_PATH.io_exuWriteback_15_bits_data_0 = U_IF_NAME.io_exuWriteback_15_bits_data_0; \
        force RTL_PATH.io_exuWriteback_15_bits_robIdx_value = U_IF_NAME.io_exuWriteback_15_bits_robIdx_value; \
        force RTL_PATH.io_exuWriteback_15_bits_fflags = U_IF_NAME.io_exuWriteback_15_bits_fflags; \
        force RTL_PATH.io_exuWriteback_15_bits_wflags = U_IF_NAME.io_exuWriteback_15_bits_wflags; \
        force RTL_PATH.io_exuWriteback_15_bits_vxsat = U_IF_NAME.io_exuWriteback_15_bits_vxsat; \
        force RTL_PATH.io_exuWriteback_14_valid = U_IF_NAME.io_exuWriteback_14_valid; \
        force RTL_PATH.io_exuWriteback_14_bits_data_0 = U_IF_NAME.io_exuWriteback_14_bits_data_0; \
        force RTL_PATH.io_exuWriteback_14_bits_robIdx_value = U_IF_NAME.io_exuWriteback_14_bits_robIdx_value; \
        force RTL_PATH.io_exuWriteback_14_bits_fflags = U_IF_NAME.io_exuWriteback_14_bits_fflags; \
        force RTL_PATH.io_exuWriteback_14_bits_wflags = U_IF_NAME.io_exuWriteback_14_bits_wflags; \
        force RTL_PATH.io_exuWriteback_13_valid = U_IF_NAME.io_exuWriteback_13_valid; \
        force RTL_PATH.io_exuWriteback_13_bits_data_0 = U_IF_NAME.io_exuWriteback_13_bits_data_0; \
        force RTL_PATH.io_exuWriteback_13_bits_robIdx_value = U_IF_NAME.io_exuWriteback_13_bits_robIdx_value; \
        force RTL_PATH.io_exuWriteback_13_bits_fflags = U_IF_NAME.io_exuWriteback_13_bits_fflags; \
        force RTL_PATH.io_exuWriteback_13_bits_wflags = U_IF_NAME.io_exuWriteback_13_bits_wflags; \
        force RTL_PATH.io_exuWriteback_13_bits_vxsat = U_IF_NAME.io_exuWriteback_13_bits_vxsat; \
        force RTL_PATH.io_exuWriteback_12_valid = U_IF_NAME.io_exuWriteback_12_valid; \
        force RTL_PATH.io_exuWriteback_12_bits_data_0 = U_IF_NAME.io_exuWriteback_12_bits_data_0; \
        force RTL_PATH.io_exuWriteback_12_bits_robIdx_value = U_IF_NAME.io_exuWriteback_12_bits_robIdx_value; \
        force RTL_PATH.io_exuWriteback_12_bits_fflags = U_IF_NAME.io_exuWriteback_12_bits_fflags; \
        force RTL_PATH.io_exuWriteback_12_bits_wflags = U_IF_NAME.io_exuWriteback_12_bits_wflags; \
        force RTL_PATH.io_exuWriteback_11_valid = U_IF_NAME.io_exuWriteback_11_valid; \
        force RTL_PATH.io_exuWriteback_11_bits_data_0 = U_IF_NAME.io_exuWriteback_11_bits_data_0; \
        force RTL_PATH.io_exuWriteback_11_bits_robIdx_value = U_IF_NAME.io_exuWriteback_11_bits_robIdx_value; \
        force RTL_PATH.io_exuWriteback_11_bits_fflags = U_IF_NAME.io_exuWriteback_11_bits_fflags; \
        force RTL_PATH.io_exuWriteback_11_bits_wflags = U_IF_NAME.io_exuWriteback_11_bits_wflags; \
        force RTL_PATH.io_exuWriteback_10_valid = U_IF_NAME.io_exuWriteback_10_valid; \
        force RTL_PATH.io_exuWriteback_10_bits_data_0 = U_IF_NAME.io_exuWriteback_10_bits_data_0; \
        force RTL_PATH.io_exuWriteback_10_bits_robIdx_value = U_IF_NAME.io_exuWriteback_10_bits_robIdx_value; \
        force RTL_PATH.io_exuWriteback_10_bits_fflags = U_IF_NAME.io_exuWriteback_10_bits_fflags; \
        force RTL_PATH.io_exuWriteback_10_bits_wflags = U_IF_NAME.io_exuWriteback_10_bits_wflags; \
        force RTL_PATH.io_exuWriteback_9_valid = U_IF_NAME.io_exuWriteback_9_valid; \
        force RTL_PATH.io_exuWriteback_9_bits_data_0 = U_IF_NAME.io_exuWriteback_9_bits_data_0; \
        force RTL_PATH.io_exuWriteback_9_bits_robIdx_value = U_IF_NAME.io_exuWriteback_9_bits_robIdx_value; \
        force RTL_PATH.io_exuWriteback_9_bits_fflags = U_IF_NAME.io_exuWriteback_9_bits_fflags; \
        force RTL_PATH.io_exuWriteback_9_bits_wflags = U_IF_NAME.io_exuWriteback_9_bits_wflags; \
        force RTL_PATH.io_exuWriteback_8_valid = U_IF_NAME.io_exuWriteback_8_valid; \
        force RTL_PATH.io_exuWriteback_8_bits_data_0 = U_IF_NAME.io_exuWriteback_8_bits_data_0; \
        force RTL_PATH.io_exuWriteback_8_bits_robIdx_value = U_IF_NAME.io_exuWriteback_8_bits_robIdx_value; \
        force RTL_PATH.io_exuWriteback_8_bits_fflags = U_IF_NAME.io_exuWriteback_8_bits_fflags; \
        force RTL_PATH.io_exuWriteback_8_bits_wflags = U_IF_NAME.io_exuWriteback_8_bits_wflags; \
        force RTL_PATH.io_exuWriteback_7_valid = U_IF_NAME.io_exuWriteback_7_valid; \
        force RTL_PATH.io_exuWriteback_7_bits_data_0 = U_IF_NAME.io_exuWriteback_7_bits_data_0; \
        force RTL_PATH.io_exuWriteback_7_bits_robIdx_value = U_IF_NAME.io_exuWriteback_7_bits_robIdx_value; \
        force RTL_PATH.io_exuWriteback_7_bits_debug_isPerfCnt = U_IF_NAME.io_exuWriteback_7_bits_debug_isPerfCnt; \
        force RTL_PATH.io_exuWriteback_6_valid = U_IF_NAME.io_exuWriteback_6_valid; \
        force RTL_PATH.io_exuWriteback_6_bits_data_0 = U_IF_NAME.io_exuWriteback_6_bits_data_0; \
        force RTL_PATH.io_exuWriteback_6_bits_robIdx_value = U_IF_NAME.io_exuWriteback_6_bits_robIdx_value; \
        force RTL_PATH.io_exuWriteback_5_valid = U_IF_NAME.io_exuWriteback_5_valid; \
        force RTL_PATH.io_exuWriteback_5_bits_data_0 = U_IF_NAME.io_exuWriteback_5_bits_data_0; \
        force RTL_PATH.io_exuWriteback_5_bits_robIdx_value = U_IF_NAME.io_exuWriteback_5_bits_robIdx_value; \
        force RTL_PATH.io_exuWriteback_5_bits_redirect_valid = U_IF_NAME.io_exuWriteback_5_bits_redirect_valid; \
        force RTL_PATH.io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken = U_IF_NAME.io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken; \
        force RTL_PATH.io_exuWriteback_5_bits_fflags = U_IF_NAME.io_exuWriteback_5_bits_fflags; \
        force RTL_PATH.io_exuWriteback_5_bits_wflags = U_IF_NAME.io_exuWriteback_5_bits_wflags; \
        force RTL_PATH.io_exuWriteback_4_valid = U_IF_NAME.io_exuWriteback_4_valid; \
        force RTL_PATH.io_exuWriteback_4_bits_data_0 = U_IF_NAME.io_exuWriteback_4_bits_data_0; \
        force RTL_PATH.io_exuWriteback_4_bits_robIdx_value = U_IF_NAME.io_exuWriteback_4_bits_robIdx_value; \
        force RTL_PATH.io_exuWriteback_3_valid = U_IF_NAME.io_exuWriteback_3_valid; \
        force RTL_PATH.io_exuWriteback_3_bits_data_0 = U_IF_NAME.io_exuWriteback_3_bits_data_0; \
        force RTL_PATH.io_exuWriteback_3_bits_robIdx_value = U_IF_NAME.io_exuWriteback_3_bits_robIdx_value; \
        force RTL_PATH.io_exuWriteback_3_bits_redirect_valid = U_IF_NAME.io_exuWriteback_3_bits_redirect_valid; \
        force RTL_PATH.io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken = U_IF_NAME.io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken; \
        force RTL_PATH.io_exuWriteback_2_valid = U_IF_NAME.io_exuWriteback_2_valid; \
        force RTL_PATH.io_exuWriteback_2_bits_data_0 = U_IF_NAME.io_exuWriteback_2_bits_data_0; \
        force RTL_PATH.io_exuWriteback_2_bits_robIdx_value = U_IF_NAME.io_exuWriteback_2_bits_robIdx_value; \
        force RTL_PATH.io_exuWriteback_1_valid = U_IF_NAME.io_exuWriteback_1_valid; \
        force RTL_PATH.io_exuWriteback_1_bits_data_0 = U_IF_NAME.io_exuWriteback_1_bits_data_0; \
        force RTL_PATH.io_exuWriteback_1_bits_robIdx_value = U_IF_NAME.io_exuWriteback_1_bits_robIdx_value; \
        force RTL_PATH.io_exuWriteback_1_bits_redirect_valid = U_IF_NAME.io_exuWriteback_1_bits_redirect_valid; \
        force RTL_PATH.io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken = U_IF_NAME.io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken; \
        force RTL_PATH.io_exuWriteback_0_valid = U_IF_NAME.io_exuWriteback_0_valid; \
        force RTL_PATH.io_exuWriteback_0_bits_data_0 = U_IF_NAME.io_exuWriteback_0_bits_data_0; \
        force RTL_PATH.io_exuWriteback_0_bits_robIdx_value = U_IF_NAME.io_exuWriteback_0_bits_robIdx_value; \
        force RTL_PATH.io_writebackNums_0_bits = U_IF_NAME.io_writebackNums_0_bits; \
        force RTL_PATH.io_writebackNums_1_bits = U_IF_NAME.io_writebackNums_1_bits; \
        force RTL_PATH.io_writebackNums_2_bits = U_IF_NAME.io_writebackNums_2_bits; \
        force RTL_PATH.io_writebackNums_3_bits = U_IF_NAME.io_writebackNums_3_bits; \
        force RTL_PATH.io_writebackNums_4_bits = U_IF_NAME.io_writebackNums_4_bits; \
        force RTL_PATH.io_writebackNums_5_bits = U_IF_NAME.io_writebackNums_5_bits; \
        force RTL_PATH.io_writebackNums_6_bits = U_IF_NAME.io_writebackNums_6_bits; \
        force RTL_PATH.io_writebackNums_7_bits = U_IF_NAME.io_writebackNums_7_bits; \
        force RTL_PATH.io_writebackNums_8_bits = U_IF_NAME.io_writebackNums_8_bits; \
        force RTL_PATH.io_writebackNums_9_bits = U_IF_NAME.io_writebackNums_9_bits; \
        force RTL_PATH.io_writebackNums_10_bits = U_IF_NAME.io_writebackNums_10_bits; \
        force RTL_PATH.io_writebackNums_11_bits = U_IF_NAME.io_writebackNums_11_bits; \
        force RTL_PATH.io_writebackNums_12_bits = U_IF_NAME.io_writebackNums_12_bits; \
        force RTL_PATH.io_writebackNums_13_bits = U_IF_NAME.io_writebackNums_13_bits; \
        force RTL_PATH.io_writebackNums_14_bits = U_IF_NAME.io_writebackNums_14_bits; \
        force RTL_PATH.io_writebackNums_15_bits = U_IF_NAME.io_writebackNums_15_bits; \
        force RTL_PATH.io_writebackNums_16_bits = U_IF_NAME.io_writebackNums_16_bits; \
        force RTL_PATH.io_writebackNums_17_bits = U_IF_NAME.io_writebackNums_17_bits; \
        force RTL_PATH.io_writebackNums_18_bits = U_IF_NAME.io_writebackNums_18_bits; \
        force RTL_PATH.io_writebackNums_19_bits = U_IF_NAME.io_writebackNums_19_bits; \
        force RTL_PATH.io_writebackNums_20_bits = U_IF_NAME.io_writebackNums_20_bits; \
        force RTL_PATH.io_writebackNums_21_bits = U_IF_NAME.io_writebackNums_21_bits; \
        force RTL_PATH.io_writebackNums_22_bits = U_IF_NAME.io_writebackNums_22_bits; \
        force RTL_PATH.io_writebackNums_23_bits = U_IF_NAME.io_writebackNums_23_bits; \
        force RTL_PATH.io_writebackNums_24_bits = U_IF_NAME.io_writebackNums_24_bits; \
        force RTL_PATH.io_writebackNeedFlush_0 = U_IF_NAME.io_writebackNeedFlush_0; \
        force RTL_PATH.io_writebackNeedFlush_1 = U_IF_NAME.io_writebackNeedFlush_1; \
        force RTL_PATH.io_writebackNeedFlush_2 = U_IF_NAME.io_writebackNeedFlush_2; \
        force RTL_PATH.io_writebackNeedFlush_6 = U_IF_NAME.io_writebackNeedFlush_6; \
        force RTL_PATH.io_writebackNeedFlush_7 = U_IF_NAME.io_writebackNeedFlush_7; \
        force RTL_PATH.io_writebackNeedFlush_8 = U_IF_NAME.io_writebackNeedFlush_8; \
        force RTL_PATH.io_writebackNeedFlush_9 = U_IF_NAME.io_writebackNeedFlush_9; \
        force RTL_PATH.io_writebackNeedFlush_10 = U_IF_NAME.io_writebackNeedFlush_10; \
        force RTL_PATH.io_writebackNeedFlush_11 = U_IF_NAME.io_writebackNeedFlush_11; \
        force RTL_PATH.io_writebackNeedFlush_12 = U_IF_NAME.io_writebackNeedFlush_12; \
    end \
    `else \
    initial begin \
        force U_IF_NAME.io_writeback_24_valid = RTL_PATH.io_writeback_24_valid; \
        force U_IF_NAME.io_writeback_24_bits_data_0 = RTL_PATH.io_writeback_24_bits_data_0; \
        force U_IF_NAME.io_writeback_24_bits_pdest = RTL_PATH.io_writeback_24_bits_pdest; \
        force U_IF_NAME.io_writeback_24_bits_robIdx_flag = RTL_PATH.io_writeback_24_bits_robIdx_flag; \
        force U_IF_NAME.io_writeback_24_bits_robIdx_value = RTL_PATH.io_writeback_24_bits_robIdx_value; \
        force U_IF_NAME.io_writeback_24_bits_vecWen = RTL_PATH.io_writeback_24_bits_vecWen; \
        force U_IF_NAME.io_writeback_24_bits_v0Wen = RTL_PATH.io_writeback_24_bits_v0Wen; \
        force U_IF_NAME.io_writeback_24_bits_vlWen = RTL_PATH.io_writeback_24_bits_vlWen; \
        force U_IF_NAME.io_writeback_24_bits_exceptionVec_0 = RTL_PATH.io_writeback_24_bits_exceptionVec_0; \
        force U_IF_NAME.io_writeback_24_bits_exceptionVec_1 = RTL_PATH.io_writeback_24_bits_exceptionVec_1; \
        force U_IF_NAME.io_writeback_24_bits_exceptionVec_2 = RTL_PATH.io_writeback_24_bits_exceptionVec_2; \
        force U_IF_NAME.io_writeback_24_bits_exceptionVec_3 = RTL_PATH.io_writeback_24_bits_exceptionVec_3; \
        force U_IF_NAME.io_writeback_24_bits_exceptionVec_4 = RTL_PATH.io_writeback_24_bits_exceptionVec_4; \
        force U_IF_NAME.io_writeback_24_bits_exceptionVec_5 = RTL_PATH.io_writeback_24_bits_exceptionVec_5; \
        force U_IF_NAME.io_writeback_24_bits_exceptionVec_6 = RTL_PATH.io_writeback_24_bits_exceptionVec_6; \
        force U_IF_NAME.io_writeback_24_bits_exceptionVec_7 = RTL_PATH.io_writeback_24_bits_exceptionVec_7; \
        force U_IF_NAME.io_writeback_24_bits_exceptionVec_8 = RTL_PATH.io_writeback_24_bits_exceptionVec_8; \
        force U_IF_NAME.io_writeback_24_bits_exceptionVec_9 = RTL_PATH.io_writeback_24_bits_exceptionVec_9; \
        force U_IF_NAME.io_writeback_24_bits_exceptionVec_10 = RTL_PATH.io_writeback_24_bits_exceptionVec_10; \
        force U_IF_NAME.io_writeback_24_bits_exceptionVec_11 = RTL_PATH.io_writeback_24_bits_exceptionVec_11; \
        force U_IF_NAME.io_writeback_24_bits_exceptionVec_12 = RTL_PATH.io_writeback_24_bits_exceptionVec_12; \
        force U_IF_NAME.io_writeback_24_bits_exceptionVec_13 = RTL_PATH.io_writeback_24_bits_exceptionVec_13; \
        force U_IF_NAME.io_writeback_24_bits_exceptionVec_14 = RTL_PATH.io_writeback_24_bits_exceptionVec_14; \
        force U_IF_NAME.io_writeback_24_bits_exceptionVec_15 = RTL_PATH.io_writeback_24_bits_exceptionVec_15; \
        force U_IF_NAME.io_writeback_24_bits_exceptionVec_16 = RTL_PATH.io_writeback_24_bits_exceptionVec_16; \
        force U_IF_NAME.io_writeback_24_bits_exceptionVec_17 = RTL_PATH.io_writeback_24_bits_exceptionVec_17; \
        force U_IF_NAME.io_writeback_24_bits_exceptionVec_18 = RTL_PATH.io_writeback_24_bits_exceptionVec_18; \
        force U_IF_NAME.io_writeback_24_bits_exceptionVec_19 = RTL_PATH.io_writeback_24_bits_exceptionVec_19; \
        force U_IF_NAME.io_writeback_24_bits_exceptionVec_20 = RTL_PATH.io_writeback_24_bits_exceptionVec_20; \
        force U_IF_NAME.io_writeback_24_bits_exceptionVec_21 = RTL_PATH.io_writeback_24_bits_exceptionVec_21; \
        force U_IF_NAME.io_writeback_24_bits_exceptionVec_22 = RTL_PATH.io_writeback_24_bits_exceptionVec_22; \
        force U_IF_NAME.io_writeback_24_bits_exceptionVec_23 = RTL_PATH.io_writeback_24_bits_exceptionVec_23; \
        force U_IF_NAME.io_writeback_24_bits_flushPipe = RTL_PATH.io_writeback_24_bits_flushPipe; \
        force U_IF_NAME.io_writeback_24_bits_replay = RTL_PATH.io_writeback_24_bits_replay; \
        force U_IF_NAME.io_writeback_24_bits_trigger = RTL_PATH.io_writeback_24_bits_trigger; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_vill = RTL_PATH.io_writeback_24_bits_vls_vpu_vill; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_vma = RTL_PATH.io_writeback_24_bits_vls_vpu_vma; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_vta = RTL_PATH.io_writeback_24_bits_vls_vpu_vta; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_vsew = RTL_PATH.io_writeback_24_bits_vls_vpu_vsew; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_vlmul = RTL_PATH.io_writeback_24_bits_vls_vpu_vlmul; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_specVill = RTL_PATH.io_writeback_24_bits_vls_vpu_specVill; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_specVma = RTL_PATH.io_writeback_24_bits_vls_vpu_specVma; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_specVta = RTL_PATH.io_writeback_24_bits_vls_vpu_specVta; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_specVsew = RTL_PATH.io_writeback_24_bits_vls_vpu_specVsew; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_specVlmul = RTL_PATH.io_writeback_24_bits_vls_vpu_specVlmul; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_vm = RTL_PATH.io_writeback_24_bits_vls_vpu_vm; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_vstart = RTL_PATH.io_writeback_24_bits_vls_vpu_vstart; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_frm = RTL_PATH.io_writeback_24_bits_vls_vpu_frm; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst = RTL_PATH.io_writeback_24_bits_vls_vpu_fpu_isFpToVecInst; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_fpu_isFP32Instr = RTL_PATH.io_writeback_24_bits_vls_vpu_fpu_isFP32Instr; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_fpu_isFP64Instr = RTL_PATH.io_writeback_24_bits_vls_vpu_fpu_isFP64Instr; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_fpu_isReduction = RTL_PATH.io_writeback_24_bits_vls_vpu_fpu_isReduction; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2 = RTL_PATH.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_2; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4 = RTL_PATH.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_4; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8 = RTL_PATH.io_writeback_24_bits_vls_vpu_fpu_isFoldTo1_8; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_vxrm = RTL_PATH.io_writeback_24_bits_vls_vpu_vxrm; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_vuopIdx = RTL_PATH.io_writeback_24_bits_vls_vpu_vuopIdx; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_lastUop = RTL_PATH.io_writeback_24_bits_vls_vpu_lastUop; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_vmask = RTL_PATH.io_writeback_24_bits_vls_vpu_vmask; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_vl = RTL_PATH.io_writeback_24_bits_vls_vpu_vl; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_nf = RTL_PATH.io_writeback_24_bits_vls_vpu_nf; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_veew = RTL_PATH.io_writeback_24_bits_vls_vpu_veew; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_isReverse = RTL_PATH.io_writeback_24_bits_vls_vpu_isReverse; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_isExt = RTL_PATH.io_writeback_24_bits_vls_vpu_isExt; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_isNarrow = RTL_PATH.io_writeback_24_bits_vls_vpu_isNarrow; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_isDstMask = RTL_PATH.io_writeback_24_bits_vls_vpu_isDstMask; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_isOpMask = RTL_PATH.io_writeback_24_bits_vls_vpu_isOpMask; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_isMove = RTL_PATH.io_writeback_24_bits_vls_vpu_isMove; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_isDependOldVd = RTL_PATH.io_writeback_24_bits_vls_vpu_isDependOldVd; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_isWritePartVd = RTL_PATH.io_writeback_24_bits_vls_vpu_isWritePartVd; \
        force U_IF_NAME.io_writeback_24_bits_vls_vpu_isVleff = RTL_PATH.io_writeback_24_bits_vls_vpu_isVleff; \
        force U_IF_NAME.io_writeback_24_bits_vls_oldVdPsrc = RTL_PATH.io_writeback_24_bits_vls_oldVdPsrc; \
        force U_IF_NAME.io_writeback_24_bits_vls_vdIdx = RTL_PATH.io_writeback_24_bits_vls_vdIdx; \
        force U_IF_NAME.io_writeback_24_bits_vls_vdIdxInField = RTL_PATH.io_writeback_24_bits_vls_vdIdxInField; \
        force U_IF_NAME.io_writeback_24_bits_vls_isIndexed = RTL_PATH.io_writeback_24_bits_vls_isIndexed; \
        force U_IF_NAME.io_writeback_24_bits_vls_isMasked = RTL_PATH.io_writeback_24_bits_vls_isMasked; \
        force U_IF_NAME.io_writeback_24_bits_vls_isStrided = RTL_PATH.io_writeback_24_bits_vls_isStrided; \
        force U_IF_NAME.io_writeback_24_bits_vls_isWhole = RTL_PATH.io_writeback_24_bits_vls_isWhole; \
        force U_IF_NAME.io_writeback_24_bits_vls_isVecLoad = RTL_PATH.io_writeback_24_bits_vls_isVecLoad; \
        force U_IF_NAME.io_writeback_24_bits_vls_isVlm = RTL_PATH.io_writeback_24_bits_vls_isVlm; \
        force U_IF_NAME.io_writeback_24_bits_debug_isMMIO = RTL_PATH.io_writeback_24_bits_debug_isMMIO; \
        force U_IF_NAME.io_writeback_24_bits_debug_isNCIO = RTL_PATH.io_writeback_24_bits_debug_isNCIO; \
        force U_IF_NAME.io_writeback_24_bits_debug_isPerfCnt = RTL_PATH.io_writeback_24_bits_debug_isPerfCnt; \
        force U_IF_NAME.io_writeback_24_bits_debug_paddr = RTL_PATH.io_writeback_24_bits_debug_paddr; \
        force U_IF_NAME.io_writeback_24_bits_debug_vaddr = RTL_PATH.io_writeback_24_bits_debug_vaddr; \
        force U_IF_NAME.io_writeback_24_bits_debugInfo_eliminatedMove = RTL_PATH.io_writeback_24_bits_debugInfo_eliminatedMove; \
        force U_IF_NAME.io_writeback_24_bits_debugInfo_renameTime = RTL_PATH.io_writeback_24_bits_debugInfo_renameTime; \
        force U_IF_NAME.io_writeback_24_bits_debugInfo_dispatchTime = RTL_PATH.io_writeback_24_bits_debugInfo_dispatchTime; \
        force U_IF_NAME.io_writeback_24_bits_debugInfo_enqRsTime = RTL_PATH.io_writeback_24_bits_debugInfo_enqRsTime; \
        force U_IF_NAME.io_writeback_24_bits_debugInfo_selectTime = RTL_PATH.io_writeback_24_bits_debugInfo_selectTime; \
        force U_IF_NAME.io_writeback_24_bits_debugInfo_issueTime = RTL_PATH.io_writeback_24_bits_debugInfo_issueTime; \
        force U_IF_NAME.io_writeback_24_bits_debugInfo_writebackTime = RTL_PATH.io_writeback_24_bits_debugInfo_writebackTime; \
        force U_IF_NAME.io_writeback_24_bits_debugInfo_runahead_checkpoint_id = RTL_PATH.io_writeback_24_bits_debugInfo_runahead_checkpoint_id; \
        force U_IF_NAME.io_writeback_24_bits_debugInfo_tlbFirstReqTime = RTL_PATH.io_writeback_24_bits_debugInfo_tlbFirstReqTime; \
        force U_IF_NAME.io_writeback_24_bits_debugInfo_tlbRespTime = RTL_PATH.io_writeback_24_bits_debugInfo_tlbRespTime; \
        force U_IF_NAME.io_writeback_24_bits_debug_seqNum = RTL_PATH.io_writeback_24_bits_debug_seqNum; \
        force U_IF_NAME.io_writeback_23_valid = RTL_PATH.io_writeback_23_valid; \
        force U_IF_NAME.io_writeback_23_bits_data_0 = RTL_PATH.io_writeback_23_bits_data_0; \
        force U_IF_NAME.io_writeback_23_bits_pdest = RTL_PATH.io_writeback_23_bits_pdest; \
        force U_IF_NAME.io_writeback_23_bits_robIdx_flag = RTL_PATH.io_writeback_23_bits_robIdx_flag; \
        force U_IF_NAME.io_writeback_23_bits_robIdx_value = RTL_PATH.io_writeback_23_bits_robIdx_value; \
        force U_IF_NAME.io_writeback_23_bits_vecWen = RTL_PATH.io_writeback_23_bits_vecWen; \
        force U_IF_NAME.io_writeback_23_bits_v0Wen = RTL_PATH.io_writeback_23_bits_v0Wen; \
        force U_IF_NAME.io_writeback_23_bits_vlWen = RTL_PATH.io_writeback_23_bits_vlWen; \
        force U_IF_NAME.io_writeback_23_bits_exceptionVec_0 = RTL_PATH.io_writeback_23_bits_exceptionVec_0; \
        force U_IF_NAME.io_writeback_23_bits_exceptionVec_1 = RTL_PATH.io_writeback_23_bits_exceptionVec_1; \
        force U_IF_NAME.io_writeback_23_bits_exceptionVec_2 = RTL_PATH.io_writeback_23_bits_exceptionVec_2; \
        force U_IF_NAME.io_writeback_23_bits_exceptionVec_3 = RTL_PATH.io_writeback_23_bits_exceptionVec_3; \
        force U_IF_NAME.io_writeback_23_bits_exceptionVec_4 = RTL_PATH.io_writeback_23_bits_exceptionVec_4; \
        force U_IF_NAME.io_writeback_23_bits_exceptionVec_5 = RTL_PATH.io_writeback_23_bits_exceptionVec_5; \
        force U_IF_NAME.io_writeback_23_bits_exceptionVec_6 = RTL_PATH.io_writeback_23_bits_exceptionVec_6; \
        force U_IF_NAME.io_writeback_23_bits_exceptionVec_7 = RTL_PATH.io_writeback_23_bits_exceptionVec_7; \
        force U_IF_NAME.io_writeback_23_bits_exceptionVec_8 = RTL_PATH.io_writeback_23_bits_exceptionVec_8; \
        force U_IF_NAME.io_writeback_23_bits_exceptionVec_9 = RTL_PATH.io_writeback_23_bits_exceptionVec_9; \
        force U_IF_NAME.io_writeback_23_bits_exceptionVec_10 = RTL_PATH.io_writeback_23_bits_exceptionVec_10; \
        force U_IF_NAME.io_writeback_23_bits_exceptionVec_11 = RTL_PATH.io_writeback_23_bits_exceptionVec_11; \
        force U_IF_NAME.io_writeback_23_bits_exceptionVec_12 = RTL_PATH.io_writeback_23_bits_exceptionVec_12; \
        force U_IF_NAME.io_writeback_23_bits_exceptionVec_13 = RTL_PATH.io_writeback_23_bits_exceptionVec_13; \
        force U_IF_NAME.io_writeback_23_bits_exceptionVec_14 = RTL_PATH.io_writeback_23_bits_exceptionVec_14; \
        force U_IF_NAME.io_writeback_23_bits_exceptionVec_15 = RTL_PATH.io_writeback_23_bits_exceptionVec_15; \
        force U_IF_NAME.io_writeback_23_bits_exceptionVec_16 = RTL_PATH.io_writeback_23_bits_exceptionVec_16; \
        force U_IF_NAME.io_writeback_23_bits_exceptionVec_17 = RTL_PATH.io_writeback_23_bits_exceptionVec_17; \
        force U_IF_NAME.io_writeback_23_bits_exceptionVec_18 = RTL_PATH.io_writeback_23_bits_exceptionVec_18; \
        force U_IF_NAME.io_writeback_23_bits_exceptionVec_19 = RTL_PATH.io_writeback_23_bits_exceptionVec_19; \
        force U_IF_NAME.io_writeback_23_bits_exceptionVec_20 = RTL_PATH.io_writeback_23_bits_exceptionVec_20; \
        force U_IF_NAME.io_writeback_23_bits_exceptionVec_21 = RTL_PATH.io_writeback_23_bits_exceptionVec_21; \
        force U_IF_NAME.io_writeback_23_bits_exceptionVec_22 = RTL_PATH.io_writeback_23_bits_exceptionVec_22; \
        force U_IF_NAME.io_writeback_23_bits_exceptionVec_23 = RTL_PATH.io_writeback_23_bits_exceptionVec_23; \
        force U_IF_NAME.io_writeback_23_bits_flushPipe = RTL_PATH.io_writeback_23_bits_flushPipe; \
        force U_IF_NAME.io_writeback_23_bits_replay = RTL_PATH.io_writeback_23_bits_replay; \
        force U_IF_NAME.io_writeback_23_bits_trigger = RTL_PATH.io_writeback_23_bits_trigger; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_vill = RTL_PATH.io_writeback_23_bits_vls_vpu_vill; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_vma = RTL_PATH.io_writeback_23_bits_vls_vpu_vma; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_vta = RTL_PATH.io_writeback_23_bits_vls_vpu_vta; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_vsew = RTL_PATH.io_writeback_23_bits_vls_vpu_vsew; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_vlmul = RTL_PATH.io_writeback_23_bits_vls_vpu_vlmul; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_specVill = RTL_PATH.io_writeback_23_bits_vls_vpu_specVill; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_specVma = RTL_PATH.io_writeback_23_bits_vls_vpu_specVma; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_specVta = RTL_PATH.io_writeback_23_bits_vls_vpu_specVta; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_specVsew = RTL_PATH.io_writeback_23_bits_vls_vpu_specVsew; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_specVlmul = RTL_PATH.io_writeback_23_bits_vls_vpu_specVlmul; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_vm = RTL_PATH.io_writeback_23_bits_vls_vpu_vm; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_vstart = RTL_PATH.io_writeback_23_bits_vls_vpu_vstart; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_frm = RTL_PATH.io_writeback_23_bits_vls_vpu_frm; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst = RTL_PATH.io_writeback_23_bits_vls_vpu_fpu_isFpToVecInst; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_fpu_isFP32Instr = RTL_PATH.io_writeback_23_bits_vls_vpu_fpu_isFP32Instr; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_fpu_isFP64Instr = RTL_PATH.io_writeback_23_bits_vls_vpu_fpu_isFP64Instr; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_fpu_isReduction = RTL_PATH.io_writeback_23_bits_vls_vpu_fpu_isReduction; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2 = RTL_PATH.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_2; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4 = RTL_PATH.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_4; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8 = RTL_PATH.io_writeback_23_bits_vls_vpu_fpu_isFoldTo1_8; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_vxrm = RTL_PATH.io_writeback_23_bits_vls_vpu_vxrm; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_vuopIdx = RTL_PATH.io_writeback_23_bits_vls_vpu_vuopIdx; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_lastUop = RTL_PATH.io_writeback_23_bits_vls_vpu_lastUop; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_vmask = RTL_PATH.io_writeback_23_bits_vls_vpu_vmask; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_vl = RTL_PATH.io_writeback_23_bits_vls_vpu_vl; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_nf = RTL_PATH.io_writeback_23_bits_vls_vpu_nf; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_veew = RTL_PATH.io_writeback_23_bits_vls_vpu_veew; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_isReverse = RTL_PATH.io_writeback_23_bits_vls_vpu_isReverse; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_isExt = RTL_PATH.io_writeback_23_bits_vls_vpu_isExt; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_isNarrow = RTL_PATH.io_writeback_23_bits_vls_vpu_isNarrow; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_isDstMask = RTL_PATH.io_writeback_23_bits_vls_vpu_isDstMask; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_isOpMask = RTL_PATH.io_writeback_23_bits_vls_vpu_isOpMask; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_isMove = RTL_PATH.io_writeback_23_bits_vls_vpu_isMove; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_isDependOldVd = RTL_PATH.io_writeback_23_bits_vls_vpu_isDependOldVd; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_isWritePartVd = RTL_PATH.io_writeback_23_bits_vls_vpu_isWritePartVd; \
        force U_IF_NAME.io_writeback_23_bits_vls_vpu_isVleff = RTL_PATH.io_writeback_23_bits_vls_vpu_isVleff; \
        force U_IF_NAME.io_writeback_23_bits_vls_oldVdPsrc = RTL_PATH.io_writeback_23_bits_vls_oldVdPsrc; \
        force U_IF_NAME.io_writeback_23_bits_vls_vdIdx = RTL_PATH.io_writeback_23_bits_vls_vdIdx; \
        force U_IF_NAME.io_writeback_23_bits_vls_vdIdxInField = RTL_PATH.io_writeback_23_bits_vls_vdIdxInField; \
        force U_IF_NAME.io_writeback_23_bits_vls_isIndexed = RTL_PATH.io_writeback_23_bits_vls_isIndexed; \
        force U_IF_NAME.io_writeback_23_bits_vls_isMasked = RTL_PATH.io_writeback_23_bits_vls_isMasked; \
        force U_IF_NAME.io_writeback_23_bits_vls_isStrided = RTL_PATH.io_writeback_23_bits_vls_isStrided; \
        force U_IF_NAME.io_writeback_23_bits_vls_isWhole = RTL_PATH.io_writeback_23_bits_vls_isWhole; \
        force U_IF_NAME.io_writeback_23_bits_vls_isVecLoad = RTL_PATH.io_writeback_23_bits_vls_isVecLoad; \
        force U_IF_NAME.io_writeback_23_bits_vls_isVlm = RTL_PATH.io_writeback_23_bits_vls_isVlm; \
        force U_IF_NAME.io_writeback_23_bits_debug_isMMIO = RTL_PATH.io_writeback_23_bits_debug_isMMIO; \
        force U_IF_NAME.io_writeback_23_bits_debug_isNCIO = RTL_PATH.io_writeback_23_bits_debug_isNCIO; \
        force U_IF_NAME.io_writeback_23_bits_debug_isPerfCnt = RTL_PATH.io_writeback_23_bits_debug_isPerfCnt; \
        force U_IF_NAME.io_writeback_23_bits_debug_paddr = RTL_PATH.io_writeback_23_bits_debug_paddr; \
        force U_IF_NAME.io_writeback_23_bits_debug_vaddr = RTL_PATH.io_writeback_23_bits_debug_vaddr; \
        force U_IF_NAME.io_writeback_23_bits_debugInfo_eliminatedMove = RTL_PATH.io_writeback_23_bits_debugInfo_eliminatedMove; \
        force U_IF_NAME.io_writeback_23_bits_debugInfo_renameTime = RTL_PATH.io_writeback_23_bits_debugInfo_renameTime; \
        force U_IF_NAME.io_writeback_23_bits_debugInfo_dispatchTime = RTL_PATH.io_writeback_23_bits_debugInfo_dispatchTime; \
        force U_IF_NAME.io_writeback_23_bits_debugInfo_enqRsTime = RTL_PATH.io_writeback_23_bits_debugInfo_enqRsTime; \
        force U_IF_NAME.io_writeback_23_bits_debugInfo_selectTime = RTL_PATH.io_writeback_23_bits_debugInfo_selectTime; \
        force U_IF_NAME.io_writeback_23_bits_debugInfo_issueTime = RTL_PATH.io_writeback_23_bits_debugInfo_issueTime; \
        force U_IF_NAME.io_writeback_23_bits_debugInfo_writebackTime = RTL_PATH.io_writeback_23_bits_debugInfo_writebackTime; \
        force U_IF_NAME.io_writeback_23_bits_debugInfo_runahead_checkpoint_id = RTL_PATH.io_writeback_23_bits_debugInfo_runahead_checkpoint_id; \
        force U_IF_NAME.io_writeback_23_bits_debugInfo_tlbFirstReqTime = RTL_PATH.io_writeback_23_bits_debugInfo_tlbFirstReqTime; \
        force U_IF_NAME.io_writeback_23_bits_debugInfo_tlbRespTime = RTL_PATH.io_writeback_23_bits_debugInfo_tlbRespTime; \
        force U_IF_NAME.io_writeback_23_bits_debug_seqNum = RTL_PATH.io_writeback_23_bits_debug_seqNum; \
        force U_IF_NAME.io_writeback_22_valid = RTL_PATH.io_writeback_22_valid; \
        force U_IF_NAME.io_writeback_22_bits_data_0 = RTL_PATH.io_writeback_22_bits_data_0; \
        force U_IF_NAME.io_writeback_22_bits_pdest = RTL_PATH.io_writeback_22_bits_pdest; \
        force U_IF_NAME.io_writeback_22_bits_robIdx_flag = RTL_PATH.io_writeback_22_bits_robIdx_flag; \
        force U_IF_NAME.io_writeback_22_bits_robIdx_value = RTL_PATH.io_writeback_22_bits_robIdx_value; \
        force U_IF_NAME.io_writeback_22_bits_intWen = RTL_PATH.io_writeback_22_bits_intWen; \
        force U_IF_NAME.io_writeback_22_bits_fpWen = RTL_PATH.io_writeback_22_bits_fpWen; \
        force U_IF_NAME.io_writeback_22_bits_exceptionVec_0 = RTL_PATH.io_writeback_22_bits_exceptionVec_0; \
        force U_IF_NAME.io_writeback_22_bits_exceptionVec_1 = RTL_PATH.io_writeback_22_bits_exceptionVec_1; \
        force U_IF_NAME.io_writeback_22_bits_exceptionVec_2 = RTL_PATH.io_writeback_22_bits_exceptionVec_2; \
        force U_IF_NAME.io_writeback_22_bits_exceptionVec_3 = RTL_PATH.io_writeback_22_bits_exceptionVec_3; \
        force U_IF_NAME.io_writeback_22_bits_exceptionVec_4 = RTL_PATH.io_writeback_22_bits_exceptionVec_4; \
        force U_IF_NAME.io_writeback_22_bits_exceptionVec_5 = RTL_PATH.io_writeback_22_bits_exceptionVec_5; \
        force U_IF_NAME.io_writeback_22_bits_exceptionVec_6 = RTL_PATH.io_writeback_22_bits_exceptionVec_6; \
        force U_IF_NAME.io_writeback_22_bits_exceptionVec_7 = RTL_PATH.io_writeback_22_bits_exceptionVec_7; \
        force U_IF_NAME.io_writeback_22_bits_exceptionVec_8 = RTL_PATH.io_writeback_22_bits_exceptionVec_8; \
        force U_IF_NAME.io_writeback_22_bits_exceptionVec_9 = RTL_PATH.io_writeback_22_bits_exceptionVec_9; \
        force U_IF_NAME.io_writeback_22_bits_exceptionVec_10 = RTL_PATH.io_writeback_22_bits_exceptionVec_10; \
        force U_IF_NAME.io_writeback_22_bits_exceptionVec_11 = RTL_PATH.io_writeback_22_bits_exceptionVec_11; \
        force U_IF_NAME.io_writeback_22_bits_exceptionVec_12 = RTL_PATH.io_writeback_22_bits_exceptionVec_12; \
        force U_IF_NAME.io_writeback_22_bits_exceptionVec_13 = RTL_PATH.io_writeback_22_bits_exceptionVec_13; \
        force U_IF_NAME.io_writeback_22_bits_exceptionVec_14 = RTL_PATH.io_writeback_22_bits_exceptionVec_14; \
        force U_IF_NAME.io_writeback_22_bits_exceptionVec_15 = RTL_PATH.io_writeback_22_bits_exceptionVec_15; \
        force U_IF_NAME.io_writeback_22_bits_exceptionVec_16 = RTL_PATH.io_writeback_22_bits_exceptionVec_16; \
        force U_IF_NAME.io_writeback_22_bits_exceptionVec_17 = RTL_PATH.io_writeback_22_bits_exceptionVec_17; \
        force U_IF_NAME.io_writeback_22_bits_exceptionVec_18 = RTL_PATH.io_writeback_22_bits_exceptionVec_18; \
        force U_IF_NAME.io_writeback_22_bits_exceptionVec_19 = RTL_PATH.io_writeback_22_bits_exceptionVec_19; \
        force U_IF_NAME.io_writeback_22_bits_exceptionVec_20 = RTL_PATH.io_writeback_22_bits_exceptionVec_20; \
        force U_IF_NAME.io_writeback_22_bits_exceptionVec_21 = RTL_PATH.io_writeback_22_bits_exceptionVec_21; \
        force U_IF_NAME.io_writeback_22_bits_exceptionVec_22 = RTL_PATH.io_writeback_22_bits_exceptionVec_22; \
        force U_IF_NAME.io_writeback_22_bits_exceptionVec_23 = RTL_PATH.io_writeback_22_bits_exceptionVec_23; \
        force U_IF_NAME.io_writeback_22_bits_flushPipe = RTL_PATH.io_writeback_22_bits_flushPipe; \
        force U_IF_NAME.io_writeback_22_bits_replay = RTL_PATH.io_writeback_22_bits_replay; \
        force U_IF_NAME.io_writeback_22_bits_lqIdx_flag = RTL_PATH.io_writeback_22_bits_lqIdx_flag; \
        force U_IF_NAME.io_writeback_22_bits_lqIdx_value = RTL_PATH.io_writeback_22_bits_lqIdx_value; \
        force U_IF_NAME.io_writeback_22_bits_trigger = RTL_PATH.io_writeback_22_bits_trigger; \
        force U_IF_NAME.io_writeback_22_bits_predecodeInfo_valid = RTL_PATH.io_writeback_22_bits_predecodeInfo_valid; \
        force U_IF_NAME.io_writeback_22_bits_predecodeInfo_isRVC = RTL_PATH.io_writeback_22_bits_predecodeInfo_isRVC; \
        force U_IF_NAME.io_writeback_22_bits_predecodeInfo_brType = RTL_PATH.io_writeback_22_bits_predecodeInfo_brType; \
        force U_IF_NAME.io_writeback_22_bits_predecodeInfo_isCall = RTL_PATH.io_writeback_22_bits_predecodeInfo_isCall; \
        force U_IF_NAME.io_writeback_22_bits_predecodeInfo_isRet = RTL_PATH.io_writeback_22_bits_predecodeInfo_isRet; \
        force U_IF_NAME.io_writeback_22_bits_debug_isMMIO = RTL_PATH.io_writeback_22_bits_debug_isMMIO; \
        force U_IF_NAME.io_writeback_22_bits_debug_isNCIO = RTL_PATH.io_writeback_22_bits_debug_isNCIO; \
        force U_IF_NAME.io_writeback_22_bits_debug_isPerfCnt = RTL_PATH.io_writeback_22_bits_debug_isPerfCnt; \
        force U_IF_NAME.io_writeback_22_bits_debug_paddr = RTL_PATH.io_writeback_22_bits_debug_paddr; \
        force U_IF_NAME.io_writeback_22_bits_debug_vaddr = RTL_PATH.io_writeback_22_bits_debug_vaddr; \
        force U_IF_NAME.io_writeback_22_bits_debugInfo_eliminatedMove = RTL_PATH.io_writeback_22_bits_debugInfo_eliminatedMove; \
        force U_IF_NAME.io_writeback_22_bits_debugInfo_renameTime = RTL_PATH.io_writeback_22_bits_debugInfo_renameTime; \
        force U_IF_NAME.io_writeback_22_bits_debugInfo_dispatchTime = RTL_PATH.io_writeback_22_bits_debugInfo_dispatchTime; \
        force U_IF_NAME.io_writeback_22_bits_debugInfo_enqRsTime = RTL_PATH.io_writeback_22_bits_debugInfo_enqRsTime; \
        force U_IF_NAME.io_writeback_22_bits_debugInfo_selectTime = RTL_PATH.io_writeback_22_bits_debugInfo_selectTime; \
        force U_IF_NAME.io_writeback_22_bits_debugInfo_issueTime = RTL_PATH.io_writeback_22_bits_debugInfo_issueTime; \
        force U_IF_NAME.io_writeback_22_bits_debugInfo_writebackTime = RTL_PATH.io_writeback_22_bits_debugInfo_writebackTime; \
        force U_IF_NAME.io_writeback_22_bits_debugInfo_runahead_checkpoint_id = RTL_PATH.io_writeback_22_bits_debugInfo_runahead_checkpoint_id; \
        force U_IF_NAME.io_writeback_22_bits_debugInfo_tlbFirstReqTime = RTL_PATH.io_writeback_22_bits_debugInfo_tlbFirstReqTime; \
        force U_IF_NAME.io_writeback_22_bits_debugInfo_tlbRespTime = RTL_PATH.io_writeback_22_bits_debugInfo_tlbRespTime; \
        force U_IF_NAME.io_writeback_22_bits_debug_seqNum = RTL_PATH.io_writeback_22_bits_debug_seqNum; \
        force U_IF_NAME.io_writeback_21_valid = RTL_PATH.io_writeback_21_valid; \
        force U_IF_NAME.io_writeback_21_bits_data_0 = RTL_PATH.io_writeback_21_bits_data_0; \
        force U_IF_NAME.io_writeback_21_bits_pdest = RTL_PATH.io_writeback_21_bits_pdest; \
        force U_IF_NAME.io_writeback_21_bits_robIdx_flag = RTL_PATH.io_writeback_21_bits_robIdx_flag; \
        force U_IF_NAME.io_writeback_21_bits_robIdx_value = RTL_PATH.io_writeback_21_bits_robIdx_value; \
        force U_IF_NAME.io_writeback_21_bits_intWen = RTL_PATH.io_writeback_21_bits_intWen; \
        force U_IF_NAME.io_writeback_21_bits_fpWen = RTL_PATH.io_writeback_21_bits_fpWen; \
        force U_IF_NAME.io_writeback_21_bits_exceptionVec_0 = RTL_PATH.io_writeback_21_bits_exceptionVec_0; \
        force U_IF_NAME.io_writeback_21_bits_exceptionVec_1 = RTL_PATH.io_writeback_21_bits_exceptionVec_1; \
        force U_IF_NAME.io_writeback_21_bits_exceptionVec_2 = RTL_PATH.io_writeback_21_bits_exceptionVec_2; \
        force U_IF_NAME.io_writeback_21_bits_exceptionVec_3 = RTL_PATH.io_writeback_21_bits_exceptionVec_3; \
        force U_IF_NAME.io_writeback_21_bits_exceptionVec_4 = RTL_PATH.io_writeback_21_bits_exceptionVec_4; \
        force U_IF_NAME.io_writeback_21_bits_exceptionVec_5 = RTL_PATH.io_writeback_21_bits_exceptionVec_5; \
        force U_IF_NAME.io_writeback_21_bits_exceptionVec_6 = RTL_PATH.io_writeback_21_bits_exceptionVec_6; \
        force U_IF_NAME.io_writeback_21_bits_exceptionVec_7 = RTL_PATH.io_writeback_21_bits_exceptionVec_7; \
        force U_IF_NAME.io_writeback_21_bits_exceptionVec_8 = RTL_PATH.io_writeback_21_bits_exceptionVec_8; \
        force U_IF_NAME.io_writeback_21_bits_exceptionVec_9 = RTL_PATH.io_writeback_21_bits_exceptionVec_9; \
        force U_IF_NAME.io_writeback_21_bits_exceptionVec_10 = RTL_PATH.io_writeback_21_bits_exceptionVec_10; \
        force U_IF_NAME.io_writeback_21_bits_exceptionVec_11 = RTL_PATH.io_writeback_21_bits_exceptionVec_11; \
        force U_IF_NAME.io_writeback_21_bits_exceptionVec_12 = RTL_PATH.io_writeback_21_bits_exceptionVec_12; \
        force U_IF_NAME.io_writeback_21_bits_exceptionVec_13 = RTL_PATH.io_writeback_21_bits_exceptionVec_13; \
        force U_IF_NAME.io_writeback_21_bits_exceptionVec_14 = RTL_PATH.io_writeback_21_bits_exceptionVec_14; \
        force U_IF_NAME.io_writeback_21_bits_exceptionVec_15 = RTL_PATH.io_writeback_21_bits_exceptionVec_15; \
        force U_IF_NAME.io_writeback_21_bits_exceptionVec_16 = RTL_PATH.io_writeback_21_bits_exceptionVec_16; \
        force U_IF_NAME.io_writeback_21_bits_exceptionVec_17 = RTL_PATH.io_writeback_21_bits_exceptionVec_17; \
        force U_IF_NAME.io_writeback_21_bits_exceptionVec_18 = RTL_PATH.io_writeback_21_bits_exceptionVec_18; \
        force U_IF_NAME.io_writeback_21_bits_exceptionVec_19 = RTL_PATH.io_writeback_21_bits_exceptionVec_19; \
        force U_IF_NAME.io_writeback_21_bits_exceptionVec_20 = RTL_PATH.io_writeback_21_bits_exceptionVec_20; \
        force U_IF_NAME.io_writeback_21_bits_exceptionVec_21 = RTL_PATH.io_writeback_21_bits_exceptionVec_21; \
        force U_IF_NAME.io_writeback_21_bits_exceptionVec_22 = RTL_PATH.io_writeback_21_bits_exceptionVec_22; \
        force U_IF_NAME.io_writeback_21_bits_exceptionVec_23 = RTL_PATH.io_writeback_21_bits_exceptionVec_23; \
        force U_IF_NAME.io_writeback_21_bits_flushPipe = RTL_PATH.io_writeback_21_bits_flushPipe; \
        force U_IF_NAME.io_writeback_21_bits_replay = RTL_PATH.io_writeback_21_bits_replay; \
        force U_IF_NAME.io_writeback_21_bits_lqIdx_flag = RTL_PATH.io_writeback_21_bits_lqIdx_flag; \
        force U_IF_NAME.io_writeback_21_bits_lqIdx_value = RTL_PATH.io_writeback_21_bits_lqIdx_value; \
        force U_IF_NAME.io_writeback_21_bits_trigger = RTL_PATH.io_writeback_21_bits_trigger; \
        force U_IF_NAME.io_writeback_21_bits_predecodeInfo_valid = RTL_PATH.io_writeback_21_bits_predecodeInfo_valid; \
        force U_IF_NAME.io_writeback_21_bits_predecodeInfo_isRVC = RTL_PATH.io_writeback_21_bits_predecodeInfo_isRVC; \
        force U_IF_NAME.io_writeback_21_bits_predecodeInfo_brType = RTL_PATH.io_writeback_21_bits_predecodeInfo_brType; \
        force U_IF_NAME.io_writeback_21_bits_predecodeInfo_isCall = RTL_PATH.io_writeback_21_bits_predecodeInfo_isCall; \
        force U_IF_NAME.io_writeback_21_bits_predecodeInfo_isRet = RTL_PATH.io_writeback_21_bits_predecodeInfo_isRet; \
        force U_IF_NAME.io_writeback_21_bits_debug_isMMIO = RTL_PATH.io_writeback_21_bits_debug_isMMIO; \
        force U_IF_NAME.io_writeback_21_bits_debug_isNCIO = RTL_PATH.io_writeback_21_bits_debug_isNCIO; \
        force U_IF_NAME.io_writeback_21_bits_debug_isPerfCnt = RTL_PATH.io_writeback_21_bits_debug_isPerfCnt; \
        force U_IF_NAME.io_writeback_21_bits_debug_paddr = RTL_PATH.io_writeback_21_bits_debug_paddr; \
        force U_IF_NAME.io_writeback_21_bits_debug_vaddr = RTL_PATH.io_writeback_21_bits_debug_vaddr; \
        force U_IF_NAME.io_writeback_21_bits_debugInfo_eliminatedMove = RTL_PATH.io_writeback_21_bits_debugInfo_eliminatedMove; \
        force U_IF_NAME.io_writeback_21_bits_debugInfo_renameTime = RTL_PATH.io_writeback_21_bits_debugInfo_renameTime; \
        force U_IF_NAME.io_writeback_21_bits_debugInfo_dispatchTime = RTL_PATH.io_writeback_21_bits_debugInfo_dispatchTime; \
        force U_IF_NAME.io_writeback_21_bits_debugInfo_enqRsTime = RTL_PATH.io_writeback_21_bits_debugInfo_enqRsTime; \
        force U_IF_NAME.io_writeback_21_bits_debugInfo_selectTime = RTL_PATH.io_writeback_21_bits_debugInfo_selectTime; \
        force U_IF_NAME.io_writeback_21_bits_debugInfo_issueTime = RTL_PATH.io_writeback_21_bits_debugInfo_issueTime; \
        force U_IF_NAME.io_writeback_21_bits_debugInfo_writebackTime = RTL_PATH.io_writeback_21_bits_debugInfo_writebackTime; \
        force U_IF_NAME.io_writeback_21_bits_debugInfo_runahead_checkpoint_id = RTL_PATH.io_writeback_21_bits_debugInfo_runahead_checkpoint_id; \
        force U_IF_NAME.io_writeback_21_bits_debugInfo_tlbFirstReqTime = RTL_PATH.io_writeback_21_bits_debugInfo_tlbFirstReqTime; \
        force U_IF_NAME.io_writeback_21_bits_debugInfo_tlbRespTime = RTL_PATH.io_writeback_21_bits_debugInfo_tlbRespTime; \
        force U_IF_NAME.io_writeback_21_bits_debug_seqNum = RTL_PATH.io_writeback_21_bits_debug_seqNum; \
        force U_IF_NAME.io_writeback_20_valid = RTL_PATH.io_writeback_20_valid; \
        force U_IF_NAME.io_writeback_20_bits_data_0 = RTL_PATH.io_writeback_20_bits_data_0; \
        force U_IF_NAME.io_writeback_20_bits_pdest = RTL_PATH.io_writeback_20_bits_pdest; \
        force U_IF_NAME.io_writeback_20_bits_robIdx_flag = RTL_PATH.io_writeback_20_bits_robIdx_flag; \
        force U_IF_NAME.io_writeback_20_bits_robIdx_value = RTL_PATH.io_writeback_20_bits_robIdx_value; \
        force U_IF_NAME.io_writeback_20_bits_intWen = RTL_PATH.io_writeback_20_bits_intWen; \
        force U_IF_NAME.io_writeback_20_bits_fpWen = RTL_PATH.io_writeback_20_bits_fpWen; \
        force U_IF_NAME.io_writeback_20_bits_exceptionVec_0 = RTL_PATH.io_writeback_20_bits_exceptionVec_0; \
        force U_IF_NAME.io_writeback_20_bits_exceptionVec_1 = RTL_PATH.io_writeback_20_bits_exceptionVec_1; \
        force U_IF_NAME.io_writeback_20_bits_exceptionVec_2 = RTL_PATH.io_writeback_20_bits_exceptionVec_2; \
        force U_IF_NAME.io_writeback_20_bits_exceptionVec_3 = RTL_PATH.io_writeback_20_bits_exceptionVec_3; \
        force U_IF_NAME.io_writeback_20_bits_exceptionVec_4 = RTL_PATH.io_writeback_20_bits_exceptionVec_4; \
        force U_IF_NAME.io_writeback_20_bits_exceptionVec_5 = RTL_PATH.io_writeback_20_bits_exceptionVec_5; \
        force U_IF_NAME.io_writeback_20_bits_exceptionVec_6 = RTL_PATH.io_writeback_20_bits_exceptionVec_6; \
        force U_IF_NAME.io_writeback_20_bits_exceptionVec_7 = RTL_PATH.io_writeback_20_bits_exceptionVec_7; \
        force U_IF_NAME.io_writeback_20_bits_exceptionVec_8 = RTL_PATH.io_writeback_20_bits_exceptionVec_8; \
        force U_IF_NAME.io_writeback_20_bits_exceptionVec_9 = RTL_PATH.io_writeback_20_bits_exceptionVec_9; \
        force U_IF_NAME.io_writeback_20_bits_exceptionVec_10 = RTL_PATH.io_writeback_20_bits_exceptionVec_10; \
        force U_IF_NAME.io_writeback_20_bits_exceptionVec_11 = RTL_PATH.io_writeback_20_bits_exceptionVec_11; \
        force U_IF_NAME.io_writeback_20_bits_exceptionVec_12 = RTL_PATH.io_writeback_20_bits_exceptionVec_12; \
        force U_IF_NAME.io_writeback_20_bits_exceptionVec_13 = RTL_PATH.io_writeback_20_bits_exceptionVec_13; \
        force U_IF_NAME.io_writeback_20_bits_exceptionVec_14 = RTL_PATH.io_writeback_20_bits_exceptionVec_14; \
        force U_IF_NAME.io_writeback_20_bits_exceptionVec_15 = RTL_PATH.io_writeback_20_bits_exceptionVec_15; \
        force U_IF_NAME.io_writeback_20_bits_exceptionVec_16 = RTL_PATH.io_writeback_20_bits_exceptionVec_16; \
        force U_IF_NAME.io_writeback_20_bits_exceptionVec_17 = RTL_PATH.io_writeback_20_bits_exceptionVec_17; \
        force U_IF_NAME.io_writeback_20_bits_exceptionVec_18 = RTL_PATH.io_writeback_20_bits_exceptionVec_18; \
        force U_IF_NAME.io_writeback_20_bits_exceptionVec_19 = RTL_PATH.io_writeback_20_bits_exceptionVec_19; \
        force U_IF_NAME.io_writeback_20_bits_exceptionVec_20 = RTL_PATH.io_writeback_20_bits_exceptionVec_20; \
        force U_IF_NAME.io_writeback_20_bits_exceptionVec_21 = RTL_PATH.io_writeback_20_bits_exceptionVec_21; \
        force U_IF_NAME.io_writeback_20_bits_exceptionVec_22 = RTL_PATH.io_writeback_20_bits_exceptionVec_22; \
        force U_IF_NAME.io_writeback_20_bits_exceptionVec_23 = RTL_PATH.io_writeback_20_bits_exceptionVec_23; \
        force U_IF_NAME.io_writeback_20_bits_flushPipe = RTL_PATH.io_writeback_20_bits_flushPipe; \
        force U_IF_NAME.io_writeback_20_bits_replay = RTL_PATH.io_writeback_20_bits_replay; \
        force U_IF_NAME.io_writeback_20_bits_lqIdx_flag = RTL_PATH.io_writeback_20_bits_lqIdx_flag; \
        force U_IF_NAME.io_writeback_20_bits_lqIdx_value = RTL_PATH.io_writeback_20_bits_lqIdx_value; \
        force U_IF_NAME.io_writeback_20_bits_trigger = RTL_PATH.io_writeback_20_bits_trigger; \
        force U_IF_NAME.io_writeback_20_bits_predecodeInfo_valid = RTL_PATH.io_writeback_20_bits_predecodeInfo_valid; \
        force U_IF_NAME.io_writeback_20_bits_predecodeInfo_isRVC = RTL_PATH.io_writeback_20_bits_predecodeInfo_isRVC; \
        force U_IF_NAME.io_writeback_20_bits_predecodeInfo_brType = RTL_PATH.io_writeback_20_bits_predecodeInfo_brType; \
        force U_IF_NAME.io_writeback_20_bits_predecodeInfo_isCall = RTL_PATH.io_writeback_20_bits_predecodeInfo_isCall; \
        force U_IF_NAME.io_writeback_20_bits_predecodeInfo_isRet = RTL_PATH.io_writeback_20_bits_predecodeInfo_isRet; \
        force U_IF_NAME.io_writeback_20_bits_debug_isMMIO = RTL_PATH.io_writeback_20_bits_debug_isMMIO; \
        force U_IF_NAME.io_writeback_20_bits_debug_isNCIO = RTL_PATH.io_writeback_20_bits_debug_isNCIO; \
        force U_IF_NAME.io_writeback_20_bits_debug_isPerfCnt = RTL_PATH.io_writeback_20_bits_debug_isPerfCnt; \
        force U_IF_NAME.io_writeback_20_bits_debug_paddr = RTL_PATH.io_writeback_20_bits_debug_paddr; \
        force U_IF_NAME.io_writeback_20_bits_debug_vaddr = RTL_PATH.io_writeback_20_bits_debug_vaddr; \
        force U_IF_NAME.io_writeback_20_bits_debugInfo_eliminatedMove = RTL_PATH.io_writeback_20_bits_debugInfo_eliminatedMove; \
        force U_IF_NAME.io_writeback_20_bits_debugInfo_renameTime = RTL_PATH.io_writeback_20_bits_debugInfo_renameTime; \
        force U_IF_NAME.io_writeback_20_bits_debugInfo_dispatchTime = RTL_PATH.io_writeback_20_bits_debugInfo_dispatchTime; \
        force U_IF_NAME.io_writeback_20_bits_debugInfo_enqRsTime = RTL_PATH.io_writeback_20_bits_debugInfo_enqRsTime; \
        force U_IF_NAME.io_writeback_20_bits_debugInfo_selectTime = RTL_PATH.io_writeback_20_bits_debugInfo_selectTime; \
        force U_IF_NAME.io_writeback_20_bits_debugInfo_issueTime = RTL_PATH.io_writeback_20_bits_debugInfo_issueTime; \
        force U_IF_NAME.io_writeback_20_bits_debugInfo_writebackTime = RTL_PATH.io_writeback_20_bits_debugInfo_writebackTime; \
        force U_IF_NAME.io_writeback_20_bits_debugInfo_runahead_checkpoint_id = RTL_PATH.io_writeback_20_bits_debugInfo_runahead_checkpoint_id; \
        force U_IF_NAME.io_writeback_20_bits_debugInfo_tlbFirstReqTime = RTL_PATH.io_writeback_20_bits_debugInfo_tlbFirstReqTime; \
        force U_IF_NAME.io_writeback_20_bits_debugInfo_tlbRespTime = RTL_PATH.io_writeback_20_bits_debugInfo_tlbRespTime; \
        force U_IF_NAME.io_writeback_20_bits_debug_seqNum = RTL_PATH.io_writeback_20_bits_debug_seqNum; \
        force U_IF_NAME.io_writeback_19_valid = RTL_PATH.io_writeback_19_valid; \
        force U_IF_NAME.io_writeback_19_bits_data_0 = RTL_PATH.io_writeback_19_bits_data_0; \
        force U_IF_NAME.io_writeback_19_bits_pdest = RTL_PATH.io_writeback_19_bits_pdest; \
        force U_IF_NAME.io_writeback_19_bits_robIdx_flag = RTL_PATH.io_writeback_19_bits_robIdx_flag; \
        force U_IF_NAME.io_writeback_19_bits_robIdx_value = RTL_PATH.io_writeback_19_bits_robIdx_value; \
        force U_IF_NAME.io_writeback_19_bits_intWen = RTL_PATH.io_writeback_19_bits_intWen; \
        force U_IF_NAME.io_writeback_19_bits_exceptionVec_0 = RTL_PATH.io_writeback_19_bits_exceptionVec_0; \
        force U_IF_NAME.io_writeback_19_bits_exceptionVec_1 = RTL_PATH.io_writeback_19_bits_exceptionVec_1; \
        force U_IF_NAME.io_writeback_19_bits_exceptionVec_2 = RTL_PATH.io_writeback_19_bits_exceptionVec_2; \
        force U_IF_NAME.io_writeback_19_bits_exceptionVec_3 = RTL_PATH.io_writeback_19_bits_exceptionVec_3; \
        force U_IF_NAME.io_writeback_19_bits_exceptionVec_4 = RTL_PATH.io_writeback_19_bits_exceptionVec_4; \
        force U_IF_NAME.io_writeback_19_bits_exceptionVec_5 = RTL_PATH.io_writeback_19_bits_exceptionVec_5; \
        force U_IF_NAME.io_writeback_19_bits_exceptionVec_6 = RTL_PATH.io_writeback_19_bits_exceptionVec_6; \
        force U_IF_NAME.io_writeback_19_bits_exceptionVec_7 = RTL_PATH.io_writeback_19_bits_exceptionVec_7; \
        force U_IF_NAME.io_writeback_19_bits_exceptionVec_8 = RTL_PATH.io_writeback_19_bits_exceptionVec_8; \
        force U_IF_NAME.io_writeback_19_bits_exceptionVec_9 = RTL_PATH.io_writeback_19_bits_exceptionVec_9; \
        force U_IF_NAME.io_writeback_19_bits_exceptionVec_10 = RTL_PATH.io_writeback_19_bits_exceptionVec_10; \
        force U_IF_NAME.io_writeback_19_bits_exceptionVec_11 = RTL_PATH.io_writeback_19_bits_exceptionVec_11; \
        force U_IF_NAME.io_writeback_19_bits_exceptionVec_12 = RTL_PATH.io_writeback_19_bits_exceptionVec_12; \
        force U_IF_NAME.io_writeback_19_bits_exceptionVec_13 = RTL_PATH.io_writeback_19_bits_exceptionVec_13; \
        force U_IF_NAME.io_writeback_19_bits_exceptionVec_14 = RTL_PATH.io_writeback_19_bits_exceptionVec_14; \
        force U_IF_NAME.io_writeback_19_bits_exceptionVec_15 = RTL_PATH.io_writeback_19_bits_exceptionVec_15; \
        force U_IF_NAME.io_writeback_19_bits_exceptionVec_16 = RTL_PATH.io_writeback_19_bits_exceptionVec_16; \
        force U_IF_NAME.io_writeback_19_bits_exceptionVec_17 = RTL_PATH.io_writeback_19_bits_exceptionVec_17; \
        force U_IF_NAME.io_writeback_19_bits_exceptionVec_18 = RTL_PATH.io_writeback_19_bits_exceptionVec_18; \
        force U_IF_NAME.io_writeback_19_bits_exceptionVec_19 = RTL_PATH.io_writeback_19_bits_exceptionVec_19; \
        force U_IF_NAME.io_writeback_19_bits_exceptionVec_20 = RTL_PATH.io_writeback_19_bits_exceptionVec_20; \
        force U_IF_NAME.io_writeback_19_bits_exceptionVec_21 = RTL_PATH.io_writeback_19_bits_exceptionVec_21; \
        force U_IF_NAME.io_writeback_19_bits_exceptionVec_22 = RTL_PATH.io_writeback_19_bits_exceptionVec_22; \
        force U_IF_NAME.io_writeback_19_bits_exceptionVec_23 = RTL_PATH.io_writeback_19_bits_exceptionVec_23; \
        force U_IF_NAME.io_writeback_19_bits_flushPipe = RTL_PATH.io_writeback_19_bits_flushPipe; \
        force U_IF_NAME.io_writeback_19_bits_sqIdx_flag = RTL_PATH.io_writeback_19_bits_sqIdx_flag; \
        force U_IF_NAME.io_writeback_19_bits_sqIdx_value = RTL_PATH.io_writeback_19_bits_sqIdx_value; \
        force U_IF_NAME.io_writeback_19_bits_trigger = RTL_PATH.io_writeback_19_bits_trigger; \
        force U_IF_NAME.io_writeback_19_bits_debug_isMMIO = RTL_PATH.io_writeback_19_bits_debug_isMMIO; \
        force U_IF_NAME.io_writeback_19_bits_debug_isNCIO = RTL_PATH.io_writeback_19_bits_debug_isNCIO; \
        force U_IF_NAME.io_writeback_19_bits_debug_isPerfCnt = RTL_PATH.io_writeback_19_bits_debug_isPerfCnt; \
        force U_IF_NAME.io_writeback_19_bits_debug_paddr = RTL_PATH.io_writeback_19_bits_debug_paddr; \
        force U_IF_NAME.io_writeback_19_bits_debug_vaddr = RTL_PATH.io_writeback_19_bits_debug_vaddr; \
        force U_IF_NAME.io_writeback_19_bits_debugInfo_eliminatedMove = RTL_PATH.io_writeback_19_bits_debugInfo_eliminatedMove; \
        force U_IF_NAME.io_writeback_19_bits_debugInfo_renameTime = RTL_PATH.io_writeback_19_bits_debugInfo_renameTime; \
        force U_IF_NAME.io_writeback_19_bits_debugInfo_dispatchTime = RTL_PATH.io_writeback_19_bits_debugInfo_dispatchTime; \
        force U_IF_NAME.io_writeback_19_bits_debugInfo_enqRsTime = RTL_PATH.io_writeback_19_bits_debugInfo_enqRsTime; \
        force U_IF_NAME.io_writeback_19_bits_debugInfo_selectTime = RTL_PATH.io_writeback_19_bits_debugInfo_selectTime; \
        force U_IF_NAME.io_writeback_19_bits_debugInfo_issueTime = RTL_PATH.io_writeback_19_bits_debugInfo_issueTime; \
        force U_IF_NAME.io_writeback_19_bits_debugInfo_writebackTime = RTL_PATH.io_writeback_19_bits_debugInfo_writebackTime; \
        force U_IF_NAME.io_writeback_19_bits_debugInfo_runahead_checkpoint_id = RTL_PATH.io_writeback_19_bits_debugInfo_runahead_checkpoint_id; \
        force U_IF_NAME.io_writeback_19_bits_debugInfo_tlbFirstReqTime = RTL_PATH.io_writeback_19_bits_debugInfo_tlbFirstReqTime; \
        force U_IF_NAME.io_writeback_19_bits_debugInfo_tlbRespTime = RTL_PATH.io_writeback_19_bits_debugInfo_tlbRespTime; \
        force U_IF_NAME.io_writeback_19_bits_debug_seqNum = RTL_PATH.io_writeback_19_bits_debug_seqNum; \
        force U_IF_NAME.io_writeback_18_valid = RTL_PATH.io_writeback_18_valid; \
        force U_IF_NAME.io_writeback_18_bits_data_0 = RTL_PATH.io_writeback_18_bits_data_0; \
        force U_IF_NAME.io_writeback_18_bits_pdest = RTL_PATH.io_writeback_18_bits_pdest; \
        force U_IF_NAME.io_writeback_18_bits_robIdx_flag = RTL_PATH.io_writeback_18_bits_robIdx_flag; \
        force U_IF_NAME.io_writeback_18_bits_robIdx_value = RTL_PATH.io_writeback_18_bits_robIdx_value; \
        force U_IF_NAME.io_writeback_18_bits_intWen = RTL_PATH.io_writeback_18_bits_intWen; \
        force U_IF_NAME.io_writeback_18_bits_exceptionVec_0 = RTL_PATH.io_writeback_18_bits_exceptionVec_0; \
        force U_IF_NAME.io_writeback_18_bits_exceptionVec_1 = RTL_PATH.io_writeback_18_bits_exceptionVec_1; \
        force U_IF_NAME.io_writeback_18_bits_exceptionVec_2 = RTL_PATH.io_writeback_18_bits_exceptionVec_2; \
        force U_IF_NAME.io_writeback_18_bits_exceptionVec_3 = RTL_PATH.io_writeback_18_bits_exceptionVec_3; \
        force U_IF_NAME.io_writeback_18_bits_exceptionVec_4 = RTL_PATH.io_writeback_18_bits_exceptionVec_4; \
        force U_IF_NAME.io_writeback_18_bits_exceptionVec_5 = RTL_PATH.io_writeback_18_bits_exceptionVec_5; \
        force U_IF_NAME.io_writeback_18_bits_exceptionVec_6 = RTL_PATH.io_writeback_18_bits_exceptionVec_6; \
        force U_IF_NAME.io_writeback_18_bits_exceptionVec_7 = RTL_PATH.io_writeback_18_bits_exceptionVec_7; \
        force U_IF_NAME.io_writeback_18_bits_exceptionVec_8 = RTL_PATH.io_writeback_18_bits_exceptionVec_8; \
        force U_IF_NAME.io_writeback_18_bits_exceptionVec_9 = RTL_PATH.io_writeback_18_bits_exceptionVec_9; \
        force U_IF_NAME.io_writeback_18_bits_exceptionVec_10 = RTL_PATH.io_writeback_18_bits_exceptionVec_10; \
        force U_IF_NAME.io_writeback_18_bits_exceptionVec_11 = RTL_PATH.io_writeback_18_bits_exceptionVec_11; \
        force U_IF_NAME.io_writeback_18_bits_exceptionVec_12 = RTL_PATH.io_writeback_18_bits_exceptionVec_12; \
        force U_IF_NAME.io_writeback_18_bits_exceptionVec_13 = RTL_PATH.io_writeback_18_bits_exceptionVec_13; \
        force U_IF_NAME.io_writeback_18_bits_exceptionVec_14 = RTL_PATH.io_writeback_18_bits_exceptionVec_14; \
        force U_IF_NAME.io_writeback_18_bits_exceptionVec_15 = RTL_PATH.io_writeback_18_bits_exceptionVec_15; \
        force U_IF_NAME.io_writeback_18_bits_exceptionVec_16 = RTL_PATH.io_writeback_18_bits_exceptionVec_16; \
        force U_IF_NAME.io_writeback_18_bits_exceptionVec_17 = RTL_PATH.io_writeback_18_bits_exceptionVec_17; \
        force U_IF_NAME.io_writeback_18_bits_exceptionVec_18 = RTL_PATH.io_writeback_18_bits_exceptionVec_18; \
        force U_IF_NAME.io_writeback_18_bits_exceptionVec_19 = RTL_PATH.io_writeback_18_bits_exceptionVec_19; \
        force U_IF_NAME.io_writeback_18_bits_exceptionVec_20 = RTL_PATH.io_writeback_18_bits_exceptionVec_20; \
        force U_IF_NAME.io_writeback_18_bits_exceptionVec_21 = RTL_PATH.io_writeback_18_bits_exceptionVec_21; \
        force U_IF_NAME.io_writeback_18_bits_exceptionVec_22 = RTL_PATH.io_writeback_18_bits_exceptionVec_22; \
        force U_IF_NAME.io_writeback_18_bits_exceptionVec_23 = RTL_PATH.io_writeback_18_bits_exceptionVec_23; \
        force U_IF_NAME.io_writeback_18_bits_flushPipe = RTL_PATH.io_writeback_18_bits_flushPipe; \
        force U_IF_NAME.io_writeback_18_bits_sqIdx_flag = RTL_PATH.io_writeback_18_bits_sqIdx_flag; \
        force U_IF_NAME.io_writeback_18_bits_sqIdx_value = RTL_PATH.io_writeback_18_bits_sqIdx_value; \
        force U_IF_NAME.io_writeback_18_bits_trigger = RTL_PATH.io_writeback_18_bits_trigger; \
        force U_IF_NAME.io_writeback_18_bits_debug_isMMIO = RTL_PATH.io_writeback_18_bits_debug_isMMIO; \
        force U_IF_NAME.io_writeback_18_bits_debug_isNCIO = RTL_PATH.io_writeback_18_bits_debug_isNCIO; \
        force U_IF_NAME.io_writeback_18_bits_debug_isPerfCnt = RTL_PATH.io_writeback_18_bits_debug_isPerfCnt; \
        force U_IF_NAME.io_writeback_18_bits_debug_paddr = RTL_PATH.io_writeback_18_bits_debug_paddr; \
        force U_IF_NAME.io_writeback_18_bits_debug_vaddr = RTL_PATH.io_writeback_18_bits_debug_vaddr; \
        force U_IF_NAME.io_writeback_18_bits_debugInfo_eliminatedMove = RTL_PATH.io_writeback_18_bits_debugInfo_eliminatedMove; \
        force U_IF_NAME.io_writeback_18_bits_debugInfo_renameTime = RTL_PATH.io_writeback_18_bits_debugInfo_renameTime; \
        force U_IF_NAME.io_writeback_18_bits_debugInfo_dispatchTime = RTL_PATH.io_writeback_18_bits_debugInfo_dispatchTime; \
        force U_IF_NAME.io_writeback_18_bits_debugInfo_enqRsTime = RTL_PATH.io_writeback_18_bits_debugInfo_enqRsTime; \
        force U_IF_NAME.io_writeback_18_bits_debugInfo_selectTime = RTL_PATH.io_writeback_18_bits_debugInfo_selectTime; \
        force U_IF_NAME.io_writeback_18_bits_debugInfo_issueTime = RTL_PATH.io_writeback_18_bits_debugInfo_issueTime; \
        force U_IF_NAME.io_writeback_18_bits_debugInfo_writebackTime = RTL_PATH.io_writeback_18_bits_debugInfo_writebackTime; \
        force U_IF_NAME.io_writeback_18_bits_debugInfo_runahead_checkpoint_id = RTL_PATH.io_writeback_18_bits_debugInfo_runahead_checkpoint_id; \
        force U_IF_NAME.io_writeback_18_bits_debugInfo_tlbFirstReqTime = RTL_PATH.io_writeback_18_bits_debugInfo_tlbFirstReqTime; \
        force U_IF_NAME.io_writeback_18_bits_debugInfo_tlbRespTime = RTL_PATH.io_writeback_18_bits_debugInfo_tlbRespTime; \
        force U_IF_NAME.io_writeback_18_bits_debug_seqNum = RTL_PATH.io_writeback_18_bits_debug_seqNum; \
        force U_IF_NAME.io_writeback_17_valid = RTL_PATH.io_writeback_17_valid; \
        force U_IF_NAME.io_writeback_17_bits_data_0 = RTL_PATH.io_writeback_17_bits_data_0; \
        force U_IF_NAME.io_writeback_17_bits_data_1 = RTL_PATH.io_writeback_17_bits_data_1; \
        force U_IF_NAME.io_writeback_17_bits_data_2 = RTL_PATH.io_writeback_17_bits_data_2; \
        force U_IF_NAME.io_writeback_17_bits_pdest = RTL_PATH.io_writeback_17_bits_pdest; \
        force U_IF_NAME.io_writeback_17_bits_robIdx_flag = RTL_PATH.io_writeback_17_bits_robIdx_flag; \
        force U_IF_NAME.io_writeback_17_bits_robIdx_value = RTL_PATH.io_writeback_17_bits_robIdx_value; \
        force U_IF_NAME.io_writeback_17_bits_vecWen = RTL_PATH.io_writeback_17_bits_vecWen; \
        force U_IF_NAME.io_writeback_17_bits_v0Wen = RTL_PATH.io_writeback_17_bits_v0Wen; \
        force U_IF_NAME.io_writeback_17_bits_fflags = RTL_PATH.io_writeback_17_bits_fflags; \
        force U_IF_NAME.io_writeback_17_bits_wflags = RTL_PATH.io_writeback_17_bits_wflags; \
        force U_IF_NAME.io_writeback_17_bits_debugInfo_eliminatedMove = RTL_PATH.io_writeback_17_bits_debugInfo_eliminatedMove; \
        force U_IF_NAME.io_writeback_17_bits_debugInfo_renameTime = RTL_PATH.io_writeback_17_bits_debugInfo_renameTime; \
        force U_IF_NAME.io_writeback_17_bits_debugInfo_dispatchTime = RTL_PATH.io_writeback_17_bits_debugInfo_dispatchTime; \
        force U_IF_NAME.io_writeback_17_bits_debugInfo_enqRsTime = RTL_PATH.io_writeback_17_bits_debugInfo_enqRsTime; \
        force U_IF_NAME.io_writeback_17_bits_debugInfo_selectTime = RTL_PATH.io_writeback_17_bits_debugInfo_selectTime; \
        force U_IF_NAME.io_writeback_17_bits_debugInfo_issueTime = RTL_PATH.io_writeback_17_bits_debugInfo_issueTime; \
        force U_IF_NAME.io_writeback_17_bits_debugInfo_writebackTime = RTL_PATH.io_writeback_17_bits_debugInfo_writebackTime; \
        force U_IF_NAME.io_writeback_17_bits_debugInfo_runahead_checkpoint_id = RTL_PATH.io_writeback_17_bits_debugInfo_runahead_checkpoint_id; \
        force U_IF_NAME.io_writeback_17_bits_debugInfo_tlbFirstReqTime = RTL_PATH.io_writeback_17_bits_debugInfo_tlbFirstReqTime; \
        force U_IF_NAME.io_writeback_17_bits_debugInfo_tlbRespTime = RTL_PATH.io_writeback_17_bits_debugInfo_tlbRespTime; \
        force U_IF_NAME.io_writeback_17_bits_debug_seqNum = RTL_PATH.io_writeback_17_bits_debug_seqNum; \
        force U_IF_NAME.io_writeback_16_valid = RTL_PATH.io_writeback_16_valid; \
        force U_IF_NAME.io_writeback_16_bits_data_0 = RTL_PATH.io_writeback_16_bits_data_0; \
        force U_IF_NAME.io_writeback_16_bits_data_1 = RTL_PATH.io_writeback_16_bits_data_1; \
        force U_IF_NAME.io_writeback_16_bits_data_2 = RTL_PATH.io_writeback_16_bits_data_2; \
        force U_IF_NAME.io_writeback_16_bits_data_3 = RTL_PATH.io_writeback_16_bits_data_3; \
        force U_IF_NAME.io_writeback_16_bits_pdest = RTL_PATH.io_writeback_16_bits_pdest; \
        force U_IF_NAME.io_writeback_16_bits_robIdx_flag = RTL_PATH.io_writeback_16_bits_robIdx_flag; \
        force U_IF_NAME.io_writeback_16_bits_robIdx_value = RTL_PATH.io_writeback_16_bits_robIdx_value; \
        force U_IF_NAME.io_writeback_16_bits_fpWen = RTL_PATH.io_writeback_16_bits_fpWen; \
        force U_IF_NAME.io_writeback_16_bits_vecWen = RTL_PATH.io_writeback_16_bits_vecWen; \
        force U_IF_NAME.io_writeback_16_bits_v0Wen = RTL_PATH.io_writeback_16_bits_v0Wen; \
        force U_IF_NAME.io_writeback_16_bits_fflags = RTL_PATH.io_writeback_16_bits_fflags; \
        force U_IF_NAME.io_writeback_16_bits_wflags = RTL_PATH.io_writeback_16_bits_wflags; \
        force U_IF_NAME.io_writeback_16_bits_debugInfo_eliminatedMove = RTL_PATH.io_writeback_16_bits_debugInfo_eliminatedMove; \
        force U_IF_NAME.io_writeback_16_bits_debugInfo_renameTime = RTL_PATH.io_writeback_16_bits_debugInfo_renameTime; \
        force U_IF_NAME.io_writeback_16_bits_debugInfo_dispatchTime = RTL_PATH.io_writeback_16_bits_debugInfo_dispatchTime; \
        force U_IF_NAME.io_writeback_16_bits_debugInfo_enqRsTime = RTL_PATH.io_writeback_16_bits_debugInfo_enqRsTime; \
        force U_IF_NAME.io_writeback_16_bits_debugInfo_selectTime = RTL_PATH.io_writeback_16_bits_debugInfo_selectTime; \
        force U_IF_NAME.io_writeback_16_bits_debugInfo_issueTime = RTL_PATH.io_writeback_16_bits_debugInfo_issueTime; \
        force U_IF_NAME.io_writeback_16_bits_debugInfo_writebackTime = RTL_PATH.io_writeback_16_bits_debugInfo_writebackTime; \
        force U_IF_NAME.io_writeback_16_bits_debugInfo_runahead_checkpoint_id = RTL_PATH.io_writeback_16_bits_debugInfo_runahead_checkpoint_id; \
        force U_IF_NAME.io_writeback_16_bits_debugInfo_tlbFirstReqTime = RTL_PATH.io_writeback_16_bits_debugInfo_tlbFirstReqTime; \
        force U_IF_NAME.io_writeback_16_bits_debugInfo_tlbRespTime = RTL_PATH.io_writeback_16_bits_debugInfo_tlbRespTime; \
        force U_IF_NAME.io_writeback_16_bits_debug_seqNum = RTL_PATH.io_writeback_16_bits_debug_seqNum; \
        force U_IF_NAME.io_writeback_15_valid = RTL_PATH.io_writeback_15_valid; \
        force U_IF_NAME.io_writeback_15_bits_data_0 = RTL_PATH.io_writeback_15_bits_data_0; \
        force U_IF_NAME.io_writeback_15_bits_data_1 = RTL_PATH.io_writeback_15_bits_data_1; \
        force U_IF_NAME.io_writeback_15_bits_data_2 = RTL_PATH.io_writeback_15_bits_data_2; \
        force U_IF_NAME.io_writeback_15_bits_pdest = RTL_PATH.io_writeback_15_bits_pdest; \
        force U_IF_NAME.io_writeback_15_bits_robIdx_flag = RTL_PATH.io_writeback_15_bits_robIdx_flag; \
        force U_IF_NAME.io_writeback_15_bits_robIdx_value = RTL_PATH.io_writeback_15_bits_robIdx_value; \
        force U_IF_NAME.io_writeback_15_bits_vecWen = RTL_PATH.io_writeback_15_bits_vecWen; \
        force U_IF_NAME.io_writeback_15_bits_v0Wen = RTL_PATH.io_writeback_15_bits_v0Wen; \
        force U_IF_NAME.io_writeback_15_bits_fflags = RTL_PATH.io_writeback_15_bits_fflags; \
        force U_IF_NAME.io_writeback_15_bits_wflags = RTL_PATH.io_writeback_15_bits_wflags; \
        force U_IF_NAME.io_writeback_15_bits_vxsat = RTL_PATH.io_writeback_15_bits_vxsat; \
        force U_IF_NAME.io_writeback_15_bits_debugInfo_eliminatedMove = RTL_PATH.io_writeback_15_bits_debugInfo_eliminatedMove; \
        force U_IF_NAME.io_writeback_15_bits_debugInfo_renameTime = RTL_PATH.io_writeback_15_bits_debugInfo_renameTime; \
        force U_IF_NAME.io_writeback_15_bits_debugInfo_dispatchTime = RTL_PATH.io_writeback_15_bits_debugInfo_dispatchTime; \
        force U_IF_NAME.io_writeback_15_bits_debugInfo_enqRsTime = RTL_PATH.io_writeback_15_bits_debugInfo_enqRsTime; \
        force U_IF_NAME.io_writeback_15_bits_debugInfo_selectTime = RTL_PATH.io_writeback_15_bits_debugInfo_selectTime; \
        force U_IF_NAME.io_writeback_15_bits_debugInfo_issueTime = RTL_PATH.io_writeback_15_bits_debugInfo_issueTime; \
        force U_IF_NAME.io_writeback_15_bits_debugInfo_writebackTime = RTL_PATH.io_writeback_15_bits_debugInfo_writebackTime; \
        force U_IF_NAME.io_writeback_15_bits_debugInfo_runahead_checkpoint_id = RTL_PATH.io_writeback_15_bits_debugInfo_runahead_checkpoint_id; \
        force U_IF_NAME.io_writeback_15_bits_debugInfo_tlbFirstReqTime = RTL_PATH.io_writeback_15_bits_debugInfo_tlbFirstReqTime; \
        force U_IF_NAME.io_writeback_15_bits_debugInfo_tlbRespTime = RTL_PATH.io_writeback_15_bits_debugInfo_tlbRespTime; \
        force U_IF_NAME.io_writeback_15_bits_debug_seqNum = RTL_PATH.io_writeback_15_bits_debug_seqNum; \
        force U_IF_NAME.io_writeback_14_valid = RTL_PATH.io_writeback_14_valid; \
        force U_IF_NAME.io_writeback_14_bits_data_0 = RTL_PATH.io_writeback_14_bits_data_0; \
        force U_IF_NAME.io_writeback_14_bits_data_1 = RTL_PATH.io_writeback_14_bits_data_1; \
        force U_IF_NAME.io_writeback_14_bits_data_2 = RTL_PATH.io_writeback_14_bits_data_2; \
        force U_IF_NAME.io_writeback_14_bits_data_3 = RTL_PATH.io_writeback_14_bits_data_3; \
        force U_IF_NAME.io_writeback_14_bits_data_4 = RTL_PATH.io_writeback_14_bits_data_4; \
        force U_IF_NAME.io_writeback_14_bits_data_5 = RTL_PATH.io_writeback_14_bits_data_5; \
        force U_IF_NAME.io_writeback_14_bits_pdest = RTL_PATH.io_writeback_14_bits_pdest; \
        force U_IF_NAME.io_writeback_14_bits_robIdx_flag = RTL_PATH.io_writeback_14_bits_robIdx_flag; \
        force U_IF_NAME.io_writeback_14_bits_robIdx_value = RTL_PATH.io_writeback_14_bits_robIdx_value; \
        force U_IF_NAME.io_writeback_14_bits_intWen = RTL_PATH.io_writeback_14_bits_intWen; \
        force U_IF_NAME.io_writeback_14_bits_fpWen = RTL_PATH.io_writeback_14_bits_fpWen; \
        force U_IF_NAME.io_writeback_14_bits_vecWen = RTL_PATH.io_writeback_14_bits_vecWen; \
        force U_IF_NAME.io_writeback_14_bits_v0Wen = RTL_PATH.io_writeback_14_bits_v0Wen; \
        force U_IF_NAME.io_writeback_14_bits_vlWen = RTL_PATH.io_writeback_14_bits_vlWen; \
        force U_IF_NAME.io_writeback_14_bits_fflags = RTL_PATH.io_writeback_14_bits_fflags; \
        force U_IF_NAME.io_writeback_14_bits_wflags = RTL_PATH.io_writeback_14_bits_wflags; \
        force U_IF_NAME.io_writeback_14_bits_exceptionVec_2 = RTL_PATH.io_writeback_14_bits_exceptionVec_2; \
        force U_IF_NAME.io_writeback_14_bits_debugInfo_eliminatedMove = RTL_PATH.io_writeback_14_bits_debugInfo_eliminatedMove; \
        force U_IF_NAME.io_writeback_14_bits_debugInfo_renameTime = RTL_PATH.io_writeback_14_bits_debugInfo_renameTime; \
        force U_IF_NAME.io_writeback_14_bits_debugInfo_dispatchTime = RTL_PATH.io_writeback_14_bits_debugInfo_dispatchTime; \
        force U_IF_NAME.io_writeback_14_bits_debugInfo_enqRsTime = RTL_PATH.io_writeback_14_bits_debugInfo_enqRsTime; \
        force U_IF_NAME.io_writeback_14_bits_debugInfo_selectTime = RTL_PATH.io_writeback_14_bits_debugInfo_selectTime; \
        force U_IF_NAME.io_writeback_14_bits_debugInfo_issueTime = RTL_PATH.io_writeback_14_bits_debugInfo_issueTime; \
        force U_IF_NAME.io_writeback_14_bits_debugInfo_writebackTime = RTL_PATH.io_writeback_14_bits_debugInfo_writebackTime; \
        force U_IF_NAME.io_writeback_14_bits_debugInfo_runahead_checkpoint_id = RTL_PATH.io_writeback_14_bits_debugInfo_runahead_checkpoint_id; \
        force U_IF_NAME.io_writeback_14_bits_debugInfo_tlbFirstReqTime = RTL_PATH.io_writeback_14_bits_debugInfo_tlbFirstReqTime; \
        force U_IF_NAME.io_writeback_14_bits_debugInfo_tlbRespTime = RTL_PATH.io_writeback_14_bits_debugInfo_tlbRespTime; \
        force U_IF_NAME.io_writeback_14_bits_debug_seqNum = RTL_PATH.io_writeback_14_bits_debug_seqNum; \
        force U_IF_NAME.io_writeback_13_valid = RTL_PATH.io_writeback_13_valid; \
        force U_IF_NAME.io_writeback_13_bits_data_0 = RTL_PATH.io_writeback_13_bits_data_0; \
        force U_IF_NAME.io_writeback_13_bits_data_1 = RTL_PATH.io_writeback_13_bits_data_1; \
        force U_IF_NAME.io_writeback_13_bits_data_2 = RTL_PATH.io_writeback_13_bits_data_2; \
        force U_IF_NAME.io_writeback_13_bits_pdest = RTL_PATH.io_writeback_13_bits_pdest; \
        force U_IF_NAME.io_writeback_13_bits_robIdx_flag = RTL_PATH.io_writeback_13_bits_robIdx_flag; \
        force U_IF_NAME.io_writeback_13_bits_robIdx_value = RTL_PATH.io_writeback_13_bits_robIdx_value; \
        force U_IF_NAME.io_writeback_13_bits_vecWen = RTL_PATH.io_writeback_13_bits_vecWen; \
        force U_IF_NAME.io_writeback_13_bits_v0Wen = RTL_PATH.io_writeback_13_bits_v0Wen; \
        force U_IF_NAME.io_writeback_13_bits_fflags = RTL_PATH.io_writeback_13_bits_fflags; \
        force U_IF_NAME.io_writeback_13_bits_wflags = RTL_PATH.io_writeback_13_bits_wflags; \
        force U_IF_NAME.io_writeback_13_bits_vxsat = RTL_PATH.io_writeback_13_bits_vxsat; \
        force U_IF_NAME.io_writeback_13_bits_exceptionVec_2 = RTL_PATH.io_writeback_13_bits_exceptionVec_2; \
        force U_IF_NAME.io_writeback_13_bits_debugInfo_eliminatedMove = RTL_PATH.io_writeback_13_bits_debugInfo_eliminatedMove; \
        force U_IF_NAME.io_writeback_13_bits_debugInfo_renameTime = RTL_PATH.io_writeback_13_bits_debugInfo_renameTime; \
        force U_IF_NAME.io_writeback_13_bits_debugInfo_dispatchTime = RTL_PATH.io_writeback_13_bits_debugInfo_dispatchTime; \
        force U_IF_NAME.io_writeback_13_bits_debugInfo_enqRsTime = RTL_PATH.io_writeback_13_bits_debugInfo_enqRsTime; \
        force U_IF_NAME.io_writeback_13_bits_debugInfo_selectTime = RTL_PATH.io_writeback_13_bits_debugInfo_selectTime; \
        force U_IF_NAME.io_writeback_13_bits_debugInfo_issueTime = RTL_PATH.io_writeback_13_bits_debugInfo_issueTime; \
        force U_IF_NAME.io_writeback_13_bits_debugInfo_writebackTime = RTL_PATH.io_writeback_13_bits_debugInfo_writebackTime; \
        force U_IF_NAME.io_writeback_13_bits_debugInfo_runahead_checkpoint_id = RTL_PATH.io_writeback_13_bits_debugInfo_runahead_checkpoint_id; \
        force U_IF_NAME.io_writeback_13_bits_debugInfo_tlbFirstReqTime = RTL_PATH.io_writeback_13_bits_debugInfo_tlbFirstReqTime; \
        force U_IF_NAME.io_writeback_13_bits_debugInfo_tlbRespTime = RTL_PATH.io_writeback_13_bits_debugInfo_tlbRespTime; \
        force U_IF_NAME.io_writeback_13_bits_debug_seqNum = RTL_PATH.io_writeback_13_bits_debug_seqNum; \
        force U_IF_NAME.io_writeback_7_valid = RTL_PATH.io_writeback_7_valid; \
        force U_IF_NAME.io_writeback_7_bits_data_0 = RTL_PATH.io_writeback_7_bits_data_0; \
        force U_IF_NAME.io_writeback_7_bits_data_1 = RTL_PATH.io_writeback_7_bits_data_1; \
        force U_IF_NAME.io_writeback_7_bits_pdest = RTL_PATH.io_writeback_7_bits_pdest; \
        force U_IF_NAME.io_writeback_7_bits_robIdx_flag = RTL_PATH.io_writeback_7_bits_robIdx_flag; \
        force U_IF_NAME.io_writeback_7_bits_robIdx_value = RTL_PATH.io_writeback_7_bits_robIdx_value; \
        force U_IF_NAME.io_writeback_7_bits_intWen = RTL_PATH.io_writeback_7_bits_intWen; \
        force U_IF_NAME.io_writeback_7_bits_redirect_valid = RTL_PATH.io_writeback_7_bits_redirect_valid; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_isRVC = RTL_PATH.io_writeback_7_bits_redirect_bits_isRVC; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_robIdx_flag = RTL_PATH.io_writeback_7_bits_redirect_bits_robIdx_flag; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_robIdx_value = RTL_PATH.io_writeback_7_bits_redirect_bits_robIdx_value; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_ftqIdx_flag = RTL_PATH.io_writeback_7_bits_redirect_bits_ftqIdx_flag; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_ftqIdx_value = RTL_PATH.io_writeback_7_bits_redirect_bits_ftqIdx_value; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_ftqOffset = RTL_PATH.io_writeback_7_bits_redirect_bits_ftqOffset; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_level = RTL_PATH.io_writeback_7_bits_redirect_bits_level; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_interrupt = RTL_PATH.io_writeback_7_bits_redirect_bits_interrupt; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_pc = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_pc; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_valid; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRVC; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_brType; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isCall; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_pd_isRet; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_ssp = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_ssp; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_sctr = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_sctr; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_flag; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSW_value; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_flag; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_TOSR_value; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_flag; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_NOS_value; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_topAddr; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0 = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1 = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2 = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3 = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0 = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1 = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2 = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3 = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_4_bits_3; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0 = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1 = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2 = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3 = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0 = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1 = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2 = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3 = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0 = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1 = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2 = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3 = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0 = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1 = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2 = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3 = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_lastBrNumOH; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_ghr = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_ghr; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_flag; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_histPtr_value; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0 = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_0; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1 = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_specCnt_1; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_br_hit; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_jr_hit; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_sc_hit; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_predTaken; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_target = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_target; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_taken = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_taken; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_isMisPred; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_shift = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_shift; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_addIntoHist; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIGPF; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIPF; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF = RTL_PATH.io_writeback_7_bits_redirect_bits_cfiUpdate_backendIAF; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_fullTarget = RTL_PATH.io_writeback_7_bits_redirect_bits_fullTarget; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_stFtqIdx_flag = RTL_PATH.io_writeback_7_bits_redirect_bits_stFtqIdx_flag; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_stFtqIdx_value = RTL_PATH.io_writeback_7_bits_redirect_bits_stFtqIdx_value; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_stFtqOffset = RTL_PATH.io_writeback_7_bits_redirect_bits_stFtqOffset; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id = RTL_PATH.io_writeback_7_bits_redirect_bits_debug_runahead_checkpoint_id; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_debugIsCtrl = RTL_PATH.io_writeback_7_bits_redirect_bits_debugIsCtrl; \
        force U_IF_NAME.io_writeback_7_bits_redirect_bits_debugIsMemVio = RTL_PATH.io_writeback_7_bits_redirect_bits_debugIsMemVio; \
        force U_IF_NAME.io_writeback_7_bits_exceptionVec_2 = RTL_PATH.io_writeback_7_bits_exceptionVec_2; \
        force U_IF_NAME.io_writeback_7_bits_exceptionVec_3 = RTL_PATH.io_writeback_7_bits_exceptionVec_3; \
        force U_IF_NAME.io_writeback_7_bits_exceptionVec_8 = RTL_PATH.io_writeback_7_bits_exceptionVec_8; \
        force U_IF_NAME.io_writeback_7_bits_exceptionVec_9 = RTL_PATH.io_writeback_7_bits_exceptionVec_9; \
        force U_IF_NAME.io_writeback_7_bits_exceptionVec_10 = RTL_PATH.io_writeback_7_bits_exceptionVec_10; \
        force U_IF_NAME.io_writeback_7_bits_exceptionVec_11 = RTL_PATH.io_writeback_7_bits_exceptionVec_11; \
        force U_IF_NAME.io_writeback_7_bits_exceptionVec_22 = RTL_PATH.io_writeback_7_bits_exceptionVec_22; \
        force U_IF_NAME.io_writeback_7_bits_flushPipe = RTL_PATH.io_writeback_7_bits_flushPipe; \
        force U_IF_NAME.io_writeback_7_bits_predecodeInfo_valid = RTL_PATH.io_writeback_7_bits_predecodeInfo_valid; \
        force U_IF_NAME.io_writeback_7_bits_predecodeInfo_isRVC = RTL_PATH.io_writeback_7_bits_predecodeInfo_isRVC; \
        force U_IF_NAME.io_writeback_7_bits_predecodeInfo_brType = RTL_PATH.io_writeback_7_bits_predecodeInfo_brType; \
        force U_IF_NAME.io_writeback_7_bits_predecodeInfo_isCall = RTL_PATH.io_writeback_7_bits_predecodeInfo_isCall; \
        force U_IF_NAME.io_writeback_7_bits_predecodeInfo_isRet = RTL_PATH.io_writeback_7_bits_predecodeInfo_isRet; \
        force U_IF_NAME.io_writeback_7_bits_debug_isPerfCnt = RTL_PATH.io_writeback_7_bits_debug_isPerfCnt; \
        force U_IF_NAME.io_writeback_7_bits_debugInfo_eliminatedMove = RTL_PATH.io_writeback_7_bits_debugInfo_eliminatedMove; \
        force U_IF_NAME.io_writeback_7_bits_debugInfo_renameTime = RTL_PATH.io_writeback_7_bits_debugInfo_renameTime; \
        force U_IF_NAME.io_writeback_7_bits_debugInfo_dispatchTime = RTL_PATH.io_writeback_7_bits_debugInfo_dispatchTime; \
        force U_IF_NAME.io_writeback_7_bits_debugInfo_enqRsTime = RTL_PATH.io_writeback_7_bits_debugInfo_enqRsTime; \
        force U_IF_NAME.io_writeback_7_bits_debugInfo_selectTime = RTL_PATH.io_writeback_7_bits_debugInfo_selectTime; \
        force U_IF_NAME.io_writeback_7_bits_debugInfo_issueTime = RTL_PATH.io_writeback_7_bits_debugInfo_issueTime; \
        force U_IF_NAME.io_writeback_7_bits_debugInfo_writebackTime = RTL_PATH.io_writeback_7_bits_debugInfo_writebackTime; \
        force U_IF_NAME.io_writeback_7_bits_debugInfo_runahead_checkpoint_id = RTL_PATH.io_writeback_7_bits_debugInfo_runahead_checkpoint_id; \
        force U_IF_NAME.io_writeback_7_bits_debugInfo_tlbFirstReqTime = RTL_PATH.io_writeback_7_bits_debugInfo_tlbFirstReqTime; \
        force U_IF_NAME.io_writeback_7_bits_debugInfo_tlbRespTime = RTL_PATH.io_writeback_7_bits_debugInfo_tlbRespTime; \
        force U_IF_NAME.io_writeback_7_bits_debug_seqNum = RTL_PATH.io_writeback_7_bits_debug_seqNum; \
        force U_IF_NAME.io_writeback_5_valid = RTL_PATH.io_writeback_5_valid; \
        force U_IF_NAME.io_writeback_5_bits_redirect_valid = RTL_PATH.io_writeback_5_bits_redirect_valid; \
        force U_IF_NAME.io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred = RTL_PATH.io_writeback_5_bits_redirect_bits_cfiUpdate_isMisPred; \
        force U_IF_NAME.io_writeback_3_valid = RTL_PATH.io_writeback_3_valid; \
        force U_IF_NAME.io_writeback_3_bits_redirect_valid = RTL_PATH.io_writeback_3_bits_redirect_valid; \
        force U_IF_NAME.io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred = RTL_PATH.io_writeback_3_bits_redirect_bits_cfiUpdate_isMisPred; \
        force U_IF_NAME.io_writeback_1_valid = RTL_PATH.io_writeback_1_valid; \
        force U_IF_NAME.io_writeback_1_bits_redirect_valid = RTL_PATH.io_writeback_1_bits_redirect_valid; \
        force U_IF_NAME.io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred = RTL_PATH.io_writeback_1_bits_redirect_bits_cfiUpdate_isMisPred; \
        force U_IF_NAME.io_exuWriteback_26_valid = RTL_PATH.io_exuWriteback_26_valid; \
        force U_IF_NAME.io_exuWriteback_26_bits_robIdx_value = RTL_PATH.io_exuWriteback_26_bits_robIdx_value; \
        force U_IF_NAME.io_exuWriteback_25_valid = RTL_PATH.io_exuWriteback_25_valid; \
        force U_IF_NAME.io_exuWriteback_25_bits_robIdx_value = RTL_PATH.io_exuWriteback_25_bits_robIdx_value; \
        force U_IF_NAME.io_exuWriteback_24_valid = RTL_PATH.io_exuWriteback_24_valid; \
        force U_IF_NAME.io_exuWriteback_24_bits_data_0 = RTL_PATH.io_exuWriteback_24_bits_data_0; \
        force U_IF_NAME.io_exuWriteback_24_bits_pdest = RTL_PATH.io_exuWriteback_24_bits_pdest; \
        force U_IF_NAME.io_exuWriteback_24_bits_robIdx_value = RTL_PATH.io_exuWriteback_24_bits_robIdx_value; \
        force U_IF_NAME.io_exuWriteback_24_bits_vecWen = RTL_PATH.io_exuWriteback_24_bits_vecWen; \
        force U_IF_NAME.io_exuWriteback_24_bits_v0Wen = RTL_PATH.io_exuWriteback_24_bits_v0Wen; \
        force U_IF_NAME.io_exuWriteback_24_bits_vls_vdIdx = RTL_PATH.io_exuWriteback_24_bits_vls_vdIdx; \
        force U_IF_NAME.io_exuWriteback_24_bits_debug_isMMIO = RTL_PATH.io_exuWriteback_24_bits_debug_isMMIO; \
        force U_IF_NAME.io_exuWriteback_24_bits_debug_isNCIO = RTL_PATH.io_exuWriteback_24_bits_debug_isNCIO; \
        force U_IF_NAME.io_exuWriteback_24_bits_debug_isPerfCnt = RTL_PATH.io_exuWriteback_24_bits_debug_isPerfCnt; \
        force U_IF_NAME.io_exuWriteback_24_bits_debug_paddr = RTL_PATH.io_exuWriteback_24_bits_debug_paddr; \
        force U_IF_NAME.io_exuWriteback_23_valid = RTL_PATH.io_exuWriteback_23_valid; \
        force U_IF_NAME.io_exuWriteback_23_bits_data_0 = RTL_PATH.io_exuWriteback_23_bits_data_0; \
        force U_IF_NAME.io_exuWriteback_23_bits_pdest = RTL_PATH.io_exuWriteback_23_bits_pdest; \
        force U_IF_NAME.io_exuWriteback_23_bits_robIdx_value = RTL_PATH.io_exuWriteback_23_bits_robIdx_value; \
        force U_IF_NAME.io_exuWriteback_23_bits_vecWen = RTL_PATH.io_exuWriteback_23_bits_vecWen; \
        force U_IF_NAME.io_exuWriteback_23_bits_v0Wen = RTL_PATH.io_exuWriteback_23_bits_v0Wen; \
        force U_IF_NAME.io_exuWriteback_23_bits_vls_vdIdx = RTL_PATH.io_exuWriteback_23_bits_vls_vdIdx; \
        force U_IF_NAME.io_exuWriteback_23_bits_debug_isMMIO = RTL_PATH.io_exuWriteback_23_bits_debug_isMMIO; \
        force U_IF_NAME.io_exuWriteback_23_bits_debug_isNCIO = RTL_PATH.io_exuWriteback_23_bits_debug_isNCIO; \
        force U_IF_NAME.io_exuWriteback_23_bits_debug_isPerfCnt = RTL_PATH.io_exuWriteback_23_bits_debug_isPerfCnt; \
        force U_IF_NAME.io_exuWriteback_23_bits_debug_paddr = RTL_PATH.io_exuWriteback_23_bits_debug_paddr; \
        force U_IF_NAME.io_exuWriteback_22_valid = RTL_PATH.io_exuWriteback_22_valid; \
        force U_IF_NAME.io_exuWriteback_22_bits_data_0 = RTL_PATH.io_exuWriteback_22_bits_data_0; \
        force U_IF_NAME.io_exuWriteback_22_bits_robIdx_value = RTL_PATH.io_exuWriteback_22_bits_robIdx_value; \
        force U_IF_NAME.io_exuWriteback_22_bits_lqIdx_value = RTL_PATH.io_exuWriteback_22_bits_lqIdx_value; \
        force U_IF_NAME.io_exuWriteback_22_bits_debug_isMMIO = RTL_PATH.io_exuWriteback_22_bits_debug_isMMIO; \
        force U_IF_NAME.io_exuWriteback_22_bits_debug_isNCIO = RTL_PATH.io_exuWriteback_22_bits_debug_isNCIO; \
        force U_IF_NAME.io_exuWriteback_22_bits_debug_isPerfCnt = RTL_PATH.io_exuWriteback_22_bits_debug_isPerfCnt; \
        force U_IF_NAME.io_exuWriteback_22_bits_debug_paddr = RTL_PATH.io_exuWriteback_22_bits_debug_paddr; \
        force U_IF_NAME.io_exuWriteback_21_valid = RTL_PATH.io_exuWriteback_21_valid; \
        force U_IF_NAME.io_exuWriteback_21_bits_data_0 = RTL_PATH.io_exuWriteback_21_bits_data_0; \
        force U_IF_NAME.io_exuWriteback_21_bits_robIdx_value = RTL_PATH.io_exuWriteback_21_bits_robIdx_value; \
        force U_IF_NAME.io_exuWriteback_21_bits_lqIdx_value = RTL_PATH.io_exuWriteback_21_bits_lqIdx_value; \
        force U_IF_NAME.io_exuWriteback_21_bits_debug_isMMIO = RTL_PATH.io_exuWriteback_21_bits_debug_isMMIO; \
        force U_IF_NAME.io_exuWriteback_21_bits_debug_isNCIO = RTL_PATH.io_exuWriteback_21_bits_debug_isNCIO; \
        force U_IF_NAME.io_exuWriteback_21_bits_debug_isPerfCnt = RTL_PATH.io_exuWriteback_21_bits_debug_isPerfCnt; \
        force U_IF_NAME.io_exuWriteback_21_bits_debug_paddr = RTL_PATH.io_exuWriteback_21_bits_debug_paddr; \
        force U_IF_NAME.io_exuWriteback_20_valid = RTL_PATH.io_exuWriteback_20_valid; \
        force U_IF_NAME.io_exuWriteback_20_bits_data_0 = RTL_PATH.io_exuWriteback_20_bits_data_0; \
        force U_IF_NAME.io_exuWriteback_20_bits_robIdx_value = RTL_PATH.io_exuWriteback_20_bits_robIdx_value; \
        force U_IF_NAME.io_exuWriteback_20_bits_lqIdx_value = RTL_PATH.io_exuWriteback_20_bits_lqIdx_value; \
        force U_IF_NAME.io_exuWriteback_20_bits_debug_isMMIO = RTL_PATH.io_exuWriteback_20_bits_debug_isMMIO; \
        force U_IF_NAME.io_exuWriteback_20_bits_debug_isNCIO = RTL_PATH.io_exuWriteback_20_bits_debug_isNCIO; \
        force U_IF_NAME.io_exuWriteback_20_bits_debug_isPerfCnt = RTL_PATH.io_exuWriteback_20_bits_debug_isPerfCnt; \
        force U_IF_NAME.io_exuWriteback_20_bits_debug_paddr = RTL_PATH.io_exuWriteback_20_bits_debug_paddr; \
        force U_IF_NAME.io_exuWriteback_19_valid = RTL_PATH.io_exuWriteback_19_valid; \
        force U_IF_NAME.io_exuWriteback_19_bits_data_0 = RTL_PATH.io_exuWriteback_19_bits_data_0; \
        force U_IF_NAME.io_exuWriteback_19_bits_robIdx_value = RTL_PATH.io_exuWriteback_19_bits_robIdx_value; \
        force U_IF_NAME.io_exuWriteback_19_bits_sqIdx_value = RTL_PATH.io_exuWriteback_19_bits_sqIdx_value; \
        force U_IF_NAME.io_exuWriteback_19_bits_debug_isMMIO = RTL_PATH.io_exuWriteback_19_bits_debug_isMMIO; \
        force U_IF_NAME.io_exuWriteback_19_bits_debug_isNCIO = RTL_PATH.io_exuWriteback_19_bits_debug_isNCIO; \
        force U_IF_NAME.io_exuWriteback_19_bits_debug_isPerfCnt = RTL_PATH.io_exuWriteback_19_bits_debug_isPerfCnt; \
        force U_IF_NAME.io_exuWriteback_19_bits_debug_paddr = RTL_PATH.io_exuWriteback_19_bits_debug_paddr; \
        force U_IF_NAME.io_exuWriteback_18_valid = RTL_PATH.io_exuWriteback_18_valid; \
        force U_IF_NAME.io_exuWriteback_18_bits_data_0 = RTL_PATH.io_exuWriteback_18_bits_data_0; \
        force U_IF_NAME.io_exuWriteback_18_bits_robIdx_value = RTL_PATH.io_exuWriteback_18_bits_robIdx_value; \
        force U_IF_NAME.io_exuWriteback_18_bits_sqIdx_value = RTL_PATH.io_exuWriteback_18_bits_sqIdx_value; \
        force U_IF_NAME.io_exuWriteback_18_bits_debug_isMMIO = RTL_PATH.io_exuWriteback_18_bits_debug_isMMIO; \
        force U_IF_NAME.io_exuWriteback_18_bits_debug_isNCIO = RTL_PATH.io_exuWriteback_18_bits_debug_isNCIO; \
        force U_IF_NAME.io_exuWriteback_18_bits_debug_isPerfCnt = RTL_PATH.io_exuWriteback_18_bits_debug_isPerfCnt; \
        force U_IF_NAME.io_exuWriteback_18_bits_debug_paddr = RTL_PATH.io_exuWriteback_18_bits_debug_paddr; \
        force U_IF_NAME.io_exuWriteback_17_valid = RTL_PATH.io_exuWriteback_17_valid; \
        force U_IF_NAME.io_exuWriteback_17_bits_data_0 = RTL_PATH.io_exuWriteback_17_bits_data_0; \
        force U_IF_NAME.io_exuWriteback_17_bits_robIdx_value = RTL_PATH.io_exuWriteback_17_bits_robIdx_value; \
        force U_IF_NAME.io_exuWriteback_17_bits_fflags = RTL_PATH.io_exuWriteback_17_bits_fflags; \
        force U_IF_NAME.io_exuWriteback_17_bits_wflags = RTL_PATH.io_exuWriteback_17_bits_wflags; \
        force U_IF_NAME.io_exuWriteback_16_valid = RTL_PATH.io_exuWriteback_16_valid; \
        force U_IF_NAME.io_exuWriteback_16_bits_data_0 = RTL_PATH.io_exuWriteback_16_bits_data_0; \
        force U_IF_NAME.io_exuWriteback_16_bits_robIdx_value = RTL_PATH.io_exuWriteback_16_bits_robIdx_value; \
        force U_IF_NAME.io_exuWriteback_16_bits_fflags = RTL_PATH.io_exuWriteback_16_bits_fflags; \
        force U_IF_NAME.io_exuWriteback_16_bits_wflags = RTL_PATH.io_exuWriteback_16_bits_wflags; \
        force U_IF_NAME.io_exuWriteback_15_valid = RTL_PATH.io_exuWriteback_15_valid; \
        force U_IF_NAME.io_exuWriteback_15_bits_data_0 = RTL_PATH.io_exuWriteback_15_bits_data_0; \
        force U_IF_NAME.io_exuWriteback_15_bits_robIdx_value = RTL_PATH.io_exuWriteback_15_bits_robIdx_value; \
        force U_IF_NAME.io_exuWriteback_15_bits_fflags = RTL_PATH.io_exuWriteback_15_bits_fflags; \
        force U_IF_NAME.io_exuWriteback_15_bits_wflags = RTL_PATH.io_exuWriteback_15_bits_wflags; \
        force U_IF_NAME.io_exuWriteback_15_bits_vxsat = RTL_PATH.io_exuWriteback_15_bits_vxsat; \
        force U_IF_NAME.io_exuWriteback_14_valid = RTL_PATH.io_exuWriteback_14_valid; \
        force U_IF_NAME.io_exuWriteback_14_bits_data_0 = RTL_PATH.io_exuWriteback_14_bits_data_0; \
        force U_IF_NAME.io_exuWriteback_14_bits_robIdx_value = RTL_PATH.io_exuWriteback_14_bits_robIdx_value; \
        force U_IF_NAME.io_exuWriteback_14_bits_fflags = RTL_PATH.io_exuWriteback_14_bits_fflags; \
        force U_IF_NAME.io_exuWriteback_14_bits_wflags = RTL_PATH.io_exuWriteback_14_bits_wflags; \
        force U_IF_NAME.io_exuWriteback_13_valid = RTL_PATH.io_exuWriteback_13_valid; \
        force U_IF_NAME.io_exuWriteback_13_bits_data_0 = RTL_PATH.io_exuWriteback_13_bits_data_0; \
        force U_IF_NAME.io_exuWriteback_13_bits_robIdx_value = RTL_PATH.io_exuWriteback_13_bits_robIdx_value; \
        force U_IF_NAME.io_exuWriteback_13_bits_fflags = RTL_PATH.io_exuWriteback_13_bits_fflags; \
        force U_IF_NAME.io_exuWriteback_13_bits_wflags = RTL_PATH.io_exuWriteback_13_bits_wflags; \
        force U_IF_NAME.io_exuWriteback_13_bits_vxsat = RTL_PATH.io_exuWriteback_13_bits_vxsat; \
        force U_IF_NAME.io_exuWriteback_12_valid = RTL_PATH.io_exuWriteback_12_valid; \
        force U_IF_NAME.io_exuWriteback_12_bits_data_0 = RTL_PATH.io_exuWriteback_12_bits_data_0; \
        force U_IF_NAME.io_exuWriteback_12_bits_robIdx_value = RTL_PATH.io_exuWriteback_12_bits_robIdx_value; \
        force U_IF_NAME.io_exuWriteback_12_bits_fflags = RTL_PATH.io_exuWriteback_12_bits_fflags; \
        force U_IF_NAME.io_exuWriteback_12_bits_wflags = RTL_PATH.io_exuWriteback_12_bits_wflags; \
        force U_IF_NAME.io_exuWriteback_11_valid = RTL_PATH.io_exuWriteback_11_valid; \
        force U_IF_NAME.io_exuWriteback_11_bits_data_0 = RTL_PATH.io_exuWriteback_11_bits_data_0; \
        force U_IF_NAME.io_exuWriteback_11_bits_robIdx_value = RTL_PATH.io_exuWriteback_11_bits_robIdx_value; \
        force U_IF_NAME.io_exuWriteback_11_bits_fflags = RTL_PATH.io_exuWriteback_11_bits_fflags; \
        force U_IF_NAME.io_exuWriteback_11_bits_wflags = RTL_PATH.io_exuWriteback_11_bits_wflags; \
        force U_IF_NAME.io_exuWriteback_10_valid = RTL_PATH.io_exuWriteback_10_valid; \
        force U_IF_NAME.io_exuWriteback_10_bits_data_0 = RTL_PATH.io_exuWriteback_10_bits_data_0; \
        force U_IF_NAME.io_exuWriteback_10_bits_robIdx_value = RTL_PATH.io_exuWriteback_10_bits_robIdx_value; \
        force U_IF_NAME.io_exuWriteback_10_bits_fflags = RTL_PATH.io_exuWriteback_10_bits_fflags; \
        force U_IF_NAME.io_exuWriteback_10_bits_wflags = RTL_PATH.io_exuWriteback_10_bits_wflags; \
        force U_IF_NAME.io_exuWriteback_9_valid = RTL_PATH.io_exuWriteback_9_valid; \
        force U_IF_NAME.io_exuWriteback_9_bits_data_0 = RTL_PATH.io_exuWriteback_9_bits_data_0; \
        force U_IF_NAME.io_exuWriteback_9_bits_robIdx_value = RTL_PATH.io_exuWriteback_9_bits_robIdx_value; \
        force U_IF_NAME.io_exuWriteback_9_bits_fflags = RTL_PATH.io_exuWriteback_9_bits_fflags; \
        force U_IF_NAME.io_exuWriteback_9_bits_wflags = RTL_PATH.io_exuWriteback_9_bits_wflags; \
        force U_IF_NAME.io_exuWriteback_8_valid = RTL_PATH.io_exuWriteback_8_valid; \
        force U_IF_NAME.io_exuWriteback_8_bits_data_0 = RTL_PATH.io_exuWriteback_8_bits_data_0; \
        force U_IF_NAME.io_exuWriteback_8_bits_robIdx_value = RTL_PATH.io_exuWriteback_8_bits_robIdx_value; \
        force U_IF_NAME.io_exuWriteback_8_bits_fflags = RTL_PATH.io_exuWriteback_8_bits_fflags; \
        force U_IF_NAME.io_exuWriteback_8_bits_wflags = RTL_PATH.io_exuWriteback_8_bits_wflags; \
        force U_IF_NAME.io_exuWriteback_7_valid = RTL_PATH.io_exuWriteback_7_valid; \
        force U_IF_NAME.io_exuWriteback_7_bits_data_0 = RTL_PATH.io_exuWriteback_7_bits_data_0; \
        force U_IF_NAME.io_exuWriteback_7_bits_robIdx_value = RTL_PATH.io_exuWriteback_7_bits_robIdx_value; \
        force U_IF_NAME.io_exuWriteback_7_bits_debug_isPerfCnt = RTL_PATH.io_exuWriteback_7_bits_debug_isPerfCnt; \
        force U_IF_NAME.io_exuWriteback_6_valid = RTL_PATH.io_exuWriteback_6_valid; \
        force U_IF_NAME.io_exuWriteback_6_bits_data_0 = RTL_PATH.io_exuWriteback_6_bits_data_0; \
        force U_IF_NAME.io_exuWriteback_6_bits_robIdx_value = RTL_PATH.io_exuWriteback_6_bits_robIdx_value; \
        force U_IF_NAME.io_exuWriteback_5_valid = RTL_PATH.io_exuWriteback_5_valid; \
        force U_IF_NAME.io_exuWriteback_5_bits_data_0 = RTL_PATH.io_exuWriteback_5_bits_data_0; \
        force U_IF_NAME.io_exuWriteback_5_bits_robIdx_value = RTL_PATH.io_exuWriteback_5_bits_robIdx_value; \
        force U_IF_NAME.io_exuWriteback_5_bits_redirect_valid = RTL_PATH.io_exuWriteback_5_bits_redirect_valid; \
        force U_IF_NAME.io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken = RTL_PATH.io_exuWriteback_5_bits_redirect_bits_cfiUpdate_taken; \
        force U_IF_NAME.io_exuWriteback_5_bits_fflags = RTL_PATH.io_exuWriteback_5_bits_fflags; \
        force U_IF_NAME.io_exuWriteback_5_bits_wflags = RTL_PATH.io_exuWriteback_5_bits_wflags; \
        force U_IF_NAME.io_exuWriteback_4_valid = RTL_PATH.io_exuWriteback_4_valid; \
        force U_IF_NAME.io_exuWriteback_4_bits_data_0 = RTL_PATH.io_exuWriteback_4_bits_data_0; \
        force U_IF_NAME.io_exuWriteback_4_bits_robIdx_value = RTL_PATH.io_exuWriteback_4_bits_robIdx_value; \
        force U_IF_NAME.io_exuWriteback_3_valid = RTL_PATH.io_exuWriteback_3_valid; \
        force U_IF_NAME.io_exuWriteback_3_bits_data_0 = RTL_PATH.io_exuWriteback_3_bits_data_0; \
        force U_IF_NAME.io_exuWriteback_3_bits_robIdx_value = RTL_PATH.io_exuWriteback_3_bits_robIdx_value; \
        force U_IF_NAME.io_exuWriteback_3_bits_redirect_valid = RTL_PATH.io_exuWriteback_3_bits_redirect_valid; \
        force U_IF_NAME.io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken = RTL_PATH.io_exuWriteback_3_bits_redirect_bits_cfiUpdate_taken; \
        force U_IF_NAME.io_exuWriteback_2_valid = RTL_PATH.io_exuWriteback_2_valid; \
        force U_IF_NAME.io_exuWriteback_2_bits_data_0 = RTL_PATH.io_exuWriteback_2_bits_data_0; \
        force U_IF_NAME.io_exuWriteback_2_bits_robIdx_value = RTL_PATH.io_exuWriteback_2_bits_robIdx_value; \
        force U_IF_NAME.io_exuWriteback_1_valid = RTL_PATH.io_exuWriteback_1_valid; \
        force U_IF_NAME.io_exuWriteback_1_bits_data_0 = RTL_PATH.io_exuWriteback_1_bits_data_0; \
        force U_IF_NAME.io_exuWriteback_1_bits_robIdx_value = RTL_PATH.io_exuWriteback_1_bits_robIdx_value; \
        force U_IF_NAME.io_exuWriteback_1_bits_redirect_valid = RTL_PATH.io_exuWriteback_1_bits_redirect_valid; \
        force U_IF_NAME.io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken = RTL_PATH.io_exuWriteback_1_bits_redirect_bits_cfiUpdate_taken; \
        force U_IF_NAME.io_exuWriteback_0_valid = RTL_PATH.io_exuWriteback_0_valid; \
        force U_IF_NAME.io_exuWriteback_0_bits_data_0 = RTL_PATH.io_exuWriteback_0_bits_data_0; \
        force U_IF_NAME.io_exuWriteback_0_bits_robIdx_value = RTL_PATH.io_exuWriteback_0_bits_robIdx_value; \
        force U_IF_NAME.io_writebackNums_0_bits = RTL_PATH.io_writebackNums_0_bits; \
        force U_IF_NAME.io_writebackNums_1_bits = RTL_PATH.io_writebackNums_1_bits; \
        force U_IF_NAME.io_writebackNums_2_bits = RTL_PATH.io_writebackNums_2_bits; \
        force U_IF_NAME.io_writebackNums_3_bits = RTL_PATH.io_writebackNums_3_bits; \
        force U_IF_NAME.io_writebackNums_4_bits = RTL_PATH.io_writebackNums_4_bits; \
        force U_IF_NAME.io_writebackNums_5_bits = RTL_PATH.io_writebackNums_5_bits; \
        force U_IF_NAME.io_writebackNums_6_bits = RTL_PATH.io_writebackNums_6_bits; \
        force U_IF_NAME.io_writebackNums_7_bits = RTL_PATH.io_writebackNums_7_bits; \
        force U_IF_NAME.io_writebackNums_8_bits = RTL_PATH.io_writebackNums_8_bits; \
        force U_IF_NAME.io_writebackNums_9_bits = RTL_PATH.io_writebackNums_9_bits; \
        force U_IF_NAME.io_writebackNums_10_bits = RTL_PATH.io_writebackNums_10_bits; \
        force U_IF_NAME.io_writebackNums_11_bits = RTL_PATH.io_writebackNums_11_bits; \
        force U_IF_NAME.io_writebackNums_12_bits = RTL_PATH.io_writebackNums_12_bits; \
        force U_IF_NAME.io_writebackNums_13_bits = RTL_PATH.io_writebackNums_13_bits; \
        force U_IF_NAME.io_writebackNums_14_bits = RTL_PATH.io_writebackNums_14_bits; \
        force U_IF_NAME.io_writebackNums_15_bits = RTL_PATH.io_writebackNums_15_bits; \
        force U_IF_NAME.io_writebackNums_16_bits = RTL_PATH.io_writebackNums_16_bits; \
        force U_IF_NAME.io_writebackNums_17_bits = RTL_PATH.io_writebackNums_17_bits; \
        force U_IF_NAME.io_writebackNums_18_bits = RTL_PATH.io_writebackNums_18_bits; \
        force U_IF_NAME.io_writebackNums_19_bits = RTL_PATH.io_writebackNums_19_bits; \
        force U_IF_NAME.io_writebackNums_20_bits = RTL_PATH.io_writebackNums_20_bits; \
        force U_IF_NAME.io_writebackNums_21_bits = RTL_PATH.io_writebackNums_21_bits; \
        force U_IF_NAME.io_writebackNums_22_bits = RTL_PATH.io_writebackNums_22_bits; \
        force U_IF_NAME.io_writebackNums_23_bits = RTL_PATH.io_writebackNums_23_bits; \
        force U_IF_NAME.io_writebackNums_24_bits = RTL_PATH.io_writebackNums_24_bits; \
        force U_IF_NAME.io_writebackNeedFlush_0 = RTL_PATH.io_writebackNeedFlush_0; \
        force U_IF_NAME.io_writebackNeedFlush_1 = RTL_PATH.io_writebackNeedFlush_1; \
        force U_IF_NAME.io_writebackNeedFlush_2 = RTL_PATH.io_writebackNeedFlush_2; \
        force U_IF_NAME.io_writebackNeedFlush_6 = RTL_PATH.io_writebackNeedFlush_6; \
        force U_IF_NAME.io_writebackNeedFlush_7 = RTL_PATH.io_writebackNeedFlush_7; \
        force U_IF_NAME.io_writebackNeedFlush_8 = RTL_PATH.io_writebackNeedFlush_8; \
        force U_IF_NAME.io_writebackNeedFlush_9 = RTL_PATH.io_writebackNeedFlush_9; \
        force U_IF_NAME.io_writebackNeedFlush_10 = RTL_PATH.io_writebackNeedFlush_10; \
        force U_IF_NAME.io_writebackNeedFlush_11 = RTL_PATH.io_writebackNeedFlush_11; \
        force U_IF_NAME.io_writebackNeedFlush_12 = RTL_PATH.io_writebackNeedFlush_12; \
    end \
    `endif

`endif

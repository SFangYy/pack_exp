//=========================================================
//File name    : rename_in_agent_dec.sv
//Author       : nanyunhao
//Module name  : rename_in_agent_dec
//Discribution : rename_in_agent_dec : parameter
//Date         : 2026-01-22
//=========================================================
`ifndef RENAME_IN_AGENT_DEC__SV
`define RENAME_IN_AGENT_DEC__SV

package rename_in_agent_dec;

endpackage:rename_in_agent_dec

import rename_in_agent_dec::*;

`endif


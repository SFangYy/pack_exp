//=========================================================
//File name    : Mem_in_agent_dec.sv
//Author       : nanyunhao
//Module name  : Mem_in_agent_dec
//Discribution : Mem_in_agent_dec : parameter
//Date         : 2026-01-22
//=========================================================
`ifndef MEM_IN_AGENT_DEC__SV
`define MEM_IN_AGENT_DEC__SV

package Mem_in_agent_dec;

endpackage:Mem_in_agent_dec

import Mem_in_agent_dec::*;

`endif

